library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestArray02_types is
-- No local datatypes implemented!


end package TestArray02_types;