package testfunction2_types;

	import scam_model_types::*;
endpackage