library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestBasic26_types is
-- No local datatypes implemented!


end package TestBasic26_types;