library ieee;
use IEEE.numeric_std.all;

package TestBasic9_types is
end package TestBasic9_types;