package testmasterslave8_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave8_SECTIONS;

endpackage
