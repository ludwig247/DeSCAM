library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave3_types is
type TestMasterSlave3_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave3_types;
