package testarray5_types;

	 import top_level_types::*;
endpackage