package testbasic8_types;

	 import top_level_types::*;
endpackage