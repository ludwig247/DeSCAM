library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave10_types is
type TestMasterSlave10_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave10_types;
