library ieee;
use IEEE.numeric_std.all;

package TestBasic1_types is
type Sections is (SECTION_A, SECTION_B);
end package TestBasic1_types;