package testbasic7_types;

endpackage