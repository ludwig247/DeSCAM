package testbasic3_types;

	typedef enum logic {
		run
	} TestBasic3_SECTIONS;

endpackage
