package testbasic21_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic21_SECTIONS;

endpackage
