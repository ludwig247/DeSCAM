constant number unsigned := 273;
constant number2 unsigned := 273;
constant number3 int := 20;
constant number4 bool := true;
