package testbasic6_types;

	 import top_level_types::*;
endpackage