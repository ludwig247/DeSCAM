library ieee;
use IEEE.numeric_std.all;
use work.SCAM_Model_types.all;

package TestArray4_types is
end package TestArray4_types;