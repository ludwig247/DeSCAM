package testbasic9_types;

	 import top_level_types::*;
endpackage