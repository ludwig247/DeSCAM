module ISA(// @[:@3.2]
    input         clock,
    // @[:@4.4]
    input         reset,
    // @[:@5.4]
    input         io_fromMemoryPort_sync,
    // @[:@6.4]
    input         io_toMemoryPort_sync,
    // @[:@6.4]
    output        io_fromMemoryPort_notify,
    // @[:@6.4]
    output        io_toMemoryPort_notify,
    // @[:@6.4]
    output        io_toRegsPort_notify,
    // @[:@6.4]
    input  [31:0] io_fromMemoryPort_loadedData,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_01,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_02,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_03,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_04,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_05,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_06,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_07,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_08,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_09,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_10,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_11,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_12,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_13,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_14,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_15,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_16,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_17,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_18,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_19,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_20,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_21,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_22,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_23,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_24,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_25,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_26,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_27,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_28,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_29,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_30,
    // @[:@6.4]
    input  [31:0] io_fromRegsPort_reg_file_31,
    // @[:@6.4]
    output [31:0] io_toMemoryPort_addrIn,
    // @[:@6.4]
    output [31:0] io_toMemoryPort_dataIn,
    // @[:@6.4]
    output [31:0] io_toMemoryPort_mask,
    // @[:@6.4]
    output [31:0] io_toMemoryPort_req,
    // @[:@6.4]
    output [31:0] io_toRegsPort_dst,
    // @[:@6.4]
    output [31:0] io_toRegsPort_dstData
    // @[:@6.4]
);
    reg             fromMemoryPort_notify_r; // @[ISA.scala 73:42:@8.4]
    reg [31:0]      _RAND_0;
    reg             toMemoryPort_notify_r; // @[ISA.scala 74:40:@9.4]
    reg [31:0]      _RAND_1;
    reg             toRegsPort_notify_r; // @[ISA.scala 75:38:@10.4]
    reg [31:0]      _RAND_2;
    reg [31:0]      toMemoryPort_r_addrIn; // @[ISA.scala 76:33:@11.4]
    reg [31:0]      _RAND_3;
    reg [31:0]      toMemoryPort_r_dataIn; // @[ISA.scala 76:33:@11.4]
    reg [31:0]      _RAND_4;
    reg [31:0]      toMemoryPort_r_mask; // @[ISA.scala 76:33:@11.4]
    reg [31:0]      _RAND_5;
    reg [31:0]      toMemoryPort_r_req; // @[ISA.scala 76:33:@11.4]
    reg [31:0]      _RAND_6;
    reg [31:0]      toRegsPort_r_dst; // @[ISA.scala 77:31:@12.4]
    reg [31:0]      _RAND_7;
    reg [31:0]      toRegsPort_r_dstData; // @[ISA.scala 77:31:@12.4]
    reg [31:0]      _RAND_8;
    reg [31:0]      memoryAccess_signal_r_addrIn; // @[ISA.scala 78:40:@13.4]
    reg [31:0]      _RAND_9;
    reg [31:0]      memoryAccess_signal_r_dataIn; // @[ISA.scala 78:40:@13.4]
    reg [31:0]      _RAND_10;
    reg [31:0]      memoryAccess_signal_r_mask; // @[ISA.scala 78:40:@13.4]
    reg [31:0]      _RAND_11;
    reg [31:0]      memoryAccess_signal_r_req; // @[ISA.scala 78:40:@13.4]
    reg [31:0]      _RAND_12;
    reg [31:0]      pcReg_signal_r; // @[ISA.scala 79:33:@14.4]
    reg [31:0]      _RAND_13;
    reg [31:0]      regfileWrite_signal_r_dst; // @[ISA.scala 80:40:@15.4]
    reg [31:0]      _RAND_14;
    reg [31:0]      regfileWrite_signal_r_dstData; // @[ISA.scala 80:40:@15.4]
    reg [31:0]      _RAND_15;
    reg [2:0]       state_r; // @[ISA.scala 81:26:@16.4]
    reg [31:0]      _RAND_16;
    wire            _T_43; // @[ISA.scala 105:30:@36.6]
    wire [2:0]      _GEN_0; // @[ISA.scala 106:52:@38.8]
    wire            _GEN_8; // @[ISA.scala 106:52:@38.8]
    wire            _GEN_9; // @[ISA.scala 106:52:@38.8]
    wire            _GEN_10; // @[ISA.scala 106:52:@38.8]
    wire [2:0]      _GEN_11; // @[ISA.scala 105:45:@37.6]
    wire            _GEN_19; // @[ISA.scala 105:45:@37.6]
    wire            _GEN_20; // @[ISA.scala 105:45:@37.6]
    wire            _GEN_21; // @[ISA.scala 105:45:@37.6]
    wire            _T_47; // @[ISA.scala 120:30:@52.6]
    wire [32:0]     _T_49; // @[ISA.scala 123:76:@56.10]
    wire [31:0]     _T_50; // @[ISA.scala 123:76:@57.10]
    wire [2:0]      _GEN_22; // @[ISA.scala 121:54:@54.8]
    wire [31:0]     _GEN_23; // @[ISA.scala 121:54:@54.8]
    wire [31:0]     _GEN_24; // @[ISA.scala 121:54:@54.8]
    wire [31:0]     _GEN_25; // @[ISA.scala 121:54:@54.8]
    wire [31:0]     _GEN_26; // @[ISA.scala 121:54:@54.8]
    wire [31:0]     _GEN_27; // @[ISA.scala 121:54:@54.8]
    wire [31:0]     _GEN_30; // @[ISA.scala 121:54:@54.8]
    wire [31:0]     _GEN_31; // @[ISA.scala 121:54:@54.8]
    wire [31:0]     _GEN_32; // @[ISA.scala 121:54:@54.8]
    wire [31:0]     _GEN_33; // @[ISA.scala 121:54:@54.8]
    wire            _GEN_34; // @[ISA.scala 121:54:@54.8]
    wire            _GEN_35; // @[ISA.scala 121:54:@54.8]
    wire            _GEN_36; // @[ISA.scala 121:54:@54.8]
    wire [2:0]      _GEN_37; // @[ISA.scala 120:45:@53.6]
    wire [31:0]     _GEN_38; // @[ISA.scala 120:45:@53.6]
    wire [31:0]     _GEN_39; // @[ISA.scala 120:45:@53.6]
    wire [31:0]     _GEN_40; // @[ISA.scala 120:45:@53.6]
    wire [31:0]     _GEN_41; // @[ISA.scala 120:45:@53.6]
    wire [31:0]     _GEN_42; // @[ISA.scala 120:45:@53.6]
    wire [31:0]     _GEN_45; // @[ISA.scala 120:45:@53.6]
    wire [31:0]     _GEN_46; // @[ISA.scala 120:45:@53.6]
    wire [31:0]     _GEN_47; // @[ISA.scala 120:45:@53.6]
    wire [31:0]     _GEN_48; // @[ISA.scala 120:45:@53.6]
    wire            _GEN_49; // @[ISA.scala 120:45:@53.6]
    wire            _GEN_50; // @[ISA.scala 120:45:@53.6]
    wire            _GEN_51; // @[ISA.scala 120:45:@53.6]
    wire            _T_62; // @[ISA.scala 139:30:@78.6]
    wire [2:0]      _GEN_52; // @[ISA.scala 140:52:@80.8]
    wire [31:0]     _GEN_53; // @[ISA.scala 140:52:@80.8]
    wire [31:0]     _GEN_54; // @[ISA.scala 140:52:@80.8]
    wire [31:0]     _GEN_55; // @[ISA.scala 140:52:@80.8]
    wire [31:0]     _GEN_56; // @[ISA.scala 140:52:@80.8]
    wire [31:0]     _GEN_57; // @[ISA.scala 140:52:@80.8]
    wire            _GEN_60; // @[ISA.scala 140:52:@80.8]
    wire            _GEN_61; // @[ISA.scala 140:52:@80.8]
    wire            _GEN_62; // @[ISA.scala 140:52:@80.8]
    wire [2:0]      _GEN_63; // @[ISA.scala 139:46:@79.6]
    wire [31:0]     _GEN_64; // @[ISA.scala 139:46:@79.6]
    wire [31:0]     _GEN_65; // @[ISA.scala 139:46:@79.6]
    wire [31:0]     _GEN_66; // @[ISA.scala 139:46:@79.6]
    wire [31:0]     _GEN_67; // @[ISA.scala 139:46:@79.6]
    wire [31:0]     _GEN_68; // @[ISA.scala 139:46:@79.6]
    wire            _GEN_71; // @[ISA.scala 139:46:@79.6]
    wire            _GEN_72; // @[ISA.scala 139:46:@79.6]
    wire            _GEN_73; // @[ISA.scala 139:46:@79.6]
    wire            _T_66; // @[ISA.scala 154:30:@94.6]
    wire [2:0]      _GEN_74; // @[ISA.scala 155:54:@96.8]
    wire [31:0]     _GEN_75; // @[ISA.scala 155:54:@96.8]
    wire [31:0]     _GEN_76; // @[ISA.scala 155:54:@96.8]
    wire [31:0]     _GEN_77; // @[ISA.scala 155:54:@96.8]
    wire [31:0]     _GEN_78; // @[ISA.scala 155:54:@96.8]
    wire [31:0]     _GEN_79; // @[ISA.scala 155:54:@96.8]
    wire [31:0]     _GEN_81; // @[ISA.scala 155:54:@96.8]
    wire [31:0]     _GEN_82; // @[ISA.scala 155:54:@96.8]
    wire [31:0]     _GEN_83; // @[ISA.scala 155:54:@96.8]
    wire [31:0]     _GEN_84; // @[ISA.scala 155:54:@96.8]
    wire [31:0]     _GEN_85; // @[ISA.scala 155:54:@96.8]
    wire [31:0]     _GEN_86; // @[ISA.scala 155:54:@96.8]
    wire [31:0]     _GEN_87; // @[ISA.scala 155:54:@96.8]
    wire            _GEN_88; // @[ISA.scala 155:54:@96.8]
    wire            _GEN_89; // @[ISA.scala 155:54:@96.8]
    wire            _GEN_90; // @[ISA.scala 155:54:@96.8]
    wire [2:0]      _GEN_91; // @[ISA.scala 154:46:@95.6]
    wire [31:0]     _GEN_92; // @[ISA.scala 154:46:@95.6]
    wire [31:0]     _GEN_93; // @[ISA.scala 154:46:@95.6]
    wire [31:0]     _GEN_94; // @[ISA.scala 154:46:@95.6]
    wire [31:0]     _GEN_95; // @[ISA.scala 154:46:@95.6]
    wire [31:0]     _GEN_96; // @[ISA.scala 154:46:@95.6]
    wire [31:0]     _GEN_98; // @[ISA.scala 154:46:@95.6]
    wire [31:0]     _GEN_99; // @[ISA.scala 154:46:@95.6]
    wire [31:0]     _GEN_100; // @[ISA.scala 154:46:@95.6]
    wire [31:0]     _GEN_101; // @[ISA.scala 154:46:@95.6]
    wire [31:0]     _GEN_102; // @[ISA.scala 154:46:@95.6]
    wire [31:0]     _GEN_103; // @[ISA.scala 154:46:@95.6]
    wire [31:0]     _GEN_104; // @[ISA.scala 154:46:@95.6]
    wire            _GEN_105; // @[ISA.scala 154:46:@95.6]
    wire            _GEN_106; // @[ISA.scala 154:46:@95.6]
    wire            _GEN_107; // @[ISA.scala 154:46:@95.6]
    wire            _T_81; // @[ISA.scala 175:30:@122.6]
    wire [2:0]      _GEN_108; // @[ISA.scala 176:52:@124.8]
    wire [31:0]     _GEN_109; // @[ISA.scala 176:52:@124.8]
    wire [31:0]     _GEN_110; // @[ISA.scala 176:52:@124.8]
    wire [31:0]     _GEN_111; // @[ISA.scala 176:52:@124.8]
    wire [31:0]     _GEN_112; // @[ISA.scala 176:52:@124.8]
    wire [31:0]     _GEN_113; // @[ISA.scala 176:52:@124.8]
    wire [31:0]     _GEN_115; // @[ISA.scala 176:52:@124.8]
    wire            _GEN_116; // @[ISA.scala 176:52:@124.8]
    wire            _GEN_117; // @[ISA.scala 176:52:@124.8]
    wire            _GEN_118; // @[ISA.scala 176:52:@124.8]
    wire [2:0]      _GEN_119; // @[ISA.scala 175:44:@123.6]
    wire [31:0]     _GEN_120; // @[ISA.scala 175:44:@123.6]
    wire [31:0]     _GEN_121; // @[ISA.scala 175:44:@123.6]
    wire [31:0]     _GEN_122; // @[ISA.scala 175:44:@123.6]
    wire [31:0]     _GEN_123; // @[ISA.scala 175:44:@123.6]
    wire [31:0]     _GEN_124; // @[ISA.scala 175:44:@123.6]
    wire [31:0]     _GEN_126; // @[ISA.scala 175:44:@123.6]
    wire            _GEN_127; // @[ISA.scala 175:44:@123.6]
    wire            _GEN_128; // @[ISA.scala 175:44:@123.6]
    wire            _GEN_129; // @[ISA.scala 175:44:@123.6]
    wire            _T_85; // @[ISA.scala 190:30:@138.6]
    wire [31:0]     _T_89; // @[ISA_functions.scala 208:38:@141.8]
    wire            _T_91; // @[ISA_functions.scala 208:53:@142.8]
    wire            _T_106; // @[ISA_functions.scala 211:28:@149.10]
    wire            _T_110; // @[ISA_functions.scala 211:108:@151.10]
    wire            _T_111; // @[ISA_functions.scala 211:75:@152.10]
    wire            _T_123; // @[ISA_functions.scala 214:78:@162.12]
    wire            _T_124; // @[ISA_functions.scala 214:75:@163.12]
    wire            _T_128; // @[ISA_functions.scala 214:158:@165.12]
    wire            _T_129; // @[ISA_functions.scala 214:125:@166.12]
    wire            _T_148; // @[ISA_functions.scala 217:128:@180.14]
    wire            _T_149; // @[ISA_functions.scala 217:125:@181.14]
    wire            _T_153; // @[ISA_functions.scala 217:207:@183.14]
    wire            _T_154; // @[ISA_functions.scala 217:174:@184.14]
    wire            _T_180; // @[ISA_functions.scala 220:177:@202.16]
    wire            _T_181; // @[ISA_functions.scala 220:174:@203.16]
    wire            _T_185; // @[ISA_functions.scala 220:258:@205.16]
    wire            _T_186; // @[ISA_functions.scala 220:225:@206.16]
    wire            _T_219; // @[ISA_functions.scala 223:228:@228.18]
    wire            _T_220; // @[ISA_functions.scala 223:225:@229.18]
    wire            _T_224; // @[ISA_functions.scala 223:308:@231.18]
    wire            _T_225; // @[ISA_functions.scala 223:275:@232.18]
    wire            _T_265; // @[ISA_functions.scala 226:278:@258.20]
    wire            _T_266; // @[ISA_functions.scala 226:275:@259.20]
    wire            _T_270; // @[ISA_functions.scala 226:359:@261.20]
    wire            _T_274; // @[ISA_functions.scala 226:408:@263.20]
    wire            _T_275; // @[ISA_functions.scala 226:375:@264.20]
    wire            _T_276; // @[ISA_functions.scala 226:325:@265.20]
    wire            _T_328; // @[ISA_functions.scala 229:328:@298.22]
    wire            _T_329; // @[ISA_functions.scala 229:325:@299.22]
    wire            _T_333; // @[ISA_functions.scala 229:459:@301.22]
    wire            _T_334; // @[ISA_functions.scala 229:426:@302.22]
    wire [31:0]     _GEN_130; // @[ISA_functions.scala 229:477:@303.22]
    wire [31:0]     _GEN_131; // @[ISA_functions.scala 226:426:@266.20]
    wire [31:0]     _GEN_132; // @[ISA_functions.scala 223:325:@233.18]
    wire [31:0]     _GEN_133; // @[ISA_functions.scala 220:275:@207.16]
    wire [31:0]     _GEN_134; // @[ISA_functions.scala 217:225:@185.14]
    wire [31:0]     _GEN_135; // @[ISA_functions.scala 214:174:@167.12]
    wire [31:0]     _GEN_136; // @[ISA_functions.scala 211:125:@153.10]
    wire [31:0]     _GEN_137; // @[ISA_functions.scala 208:70:@143.8]
    wire            _T_335; // @[ISA.scala 191:73:@309.8]
    wire            _T_337; // @[ISA.scala 191:30:@310.8]
    wire            _T_578; // @[ISA.scala 192:81:@481.10]
    wire            _T_580; // @[ISA.scala 192:38:@482.10]
    wire            _T_821; // @[ISA.scala 193:89:@653.12]
    wire            _T_823; // @[ISA.scala 193:46:@654.12]
    wire            _T_1064; // @[ISA.scala 194:97:@825.14]
    wire            _T_1066; // @[ISA.scala 194:54:@826.14]
    wire            _T_1307; // @[ISA.scala 195:105:@997.16]
    wire            _T_1309; // @[ISA.scala 195:62:@998.16]
    wire            _T_1550; // @[ISA.scala 196:113:@1169.18]
    wire            _T_1552; // @[ISA.scala 196:70:@1170.18]
    wire            _T_1793; // @[ISA.scala 197:121:@1341.20]
    wire            _T_1795; // @[ISA.scala 197:78:@1342.20]
    wire            _T_2036; // @[ISA.scala 198:129:@1513.22]
    wire            _T_2038; // @[ISA.scala 198:86:@1514.22]
    wire [2:0]      _GEN_194; // @[ISA.scala 199:118:@1516.24]
    wire [31:0]     _GEN_195; // @[ISA.scala 199:118:@1516.24]
    wire [31:0]     _GEN_196; // @[ISA.scala 199:118:@1516.24]
    wire [31:0]     _GEN_197; // @[ISA.scala 199:118:@1516.24]
    wire [31:0]     _GEN_198; // @[ISA.scala 199:118:@1516.24]
    wire [31:0]     _GEN_199; // @[ISA.scala 199:118:@1516.24]
    wire [31:0]     _GEN_201; // @[ISA.scala 199:118:@1516.24]
    wire [31:0]     _GEN_202; // @[ISA.scala 199:118:@1516.24]
    wire [31:0]     _GEN_203; // @[ISA.scala 199:118:@1516.24]
    wire [31:0]     _GEN_204; // @[ISA.scala 199:118:@1516.24]
    wire [31:0]     _GEN_205; // @[ISA.scala 199:118:@1516.24]
    wire            _GEN_206; // @[ISA.scala 199:118:@1516.24]
    wire            _GEN_207; // @[ISA.scala 199:118:@1516.24]
    wire            _GEN_208; // @[ISA.scala 199:118:@1516.24]
    wire [2:0]      _GEN_209; // @[ISA.scala 198:143:@1515.22]
    wire [31:0]     _GEN_210; // @[ISA.scala 198:143:@1515.22]
    wire [31:0]     _GEN_211; // @[ISA.scala 198:143:@1515.22]
    wire [31:0]     _GEN_212; // @[ISA.scala 198:143:@1515.22]
    wire [31:0]     _GEN_213; // @[ISA.scala 198:143:@1515.22]
    wire [31:0]     _GEN_214; // @[ISA.scala 198:143:@1515.22]
    wire [31:0]     _GEN_216; // @[ISA.scala 198:143:@1515.22]
    wire [31:0]     _GEN_217; // @[ISA.scala 198:143:@1515.22]
    wire [31:0]     _GEN_218; // @[ISA.scala 198:143:@1515.22]
    wire [31:0]     _GEN_219; // @[ISA.scala 198:143:@1515.22]
    wire [31:0]     _GEN_220; // @[ISA.scala 198:143:@1515.22]
    wire            _GEN_221; // @[ISA.scala 198:143:@1515.22]
    wire            _GEN_222; // @[ISA.scala 198:143:@1515.22]
    wire            _GEN_223; // @[ISA.scala 198:143:@1515.22]
    wire [2:0]      _GEN_224; // @[ISA.scala 197:135:@1343.20]
    wire [31:0]     _GEN_225; // @[ISA.scala 197:135:@1343.20]
    wire [31:0]     _GEN_226; // @[ISA.scala 197:135:@1343.20]
    wire [31:0]     _GEN_227; // @[ISA.scala 197:135:@1343.20]
    wire [31:0]     _GEN_228; // @[ISA.scala 197:135:@1343.20]
    wire [31:0]     _GEN_229; // @[ISA.scala 197:135:@1343.20]
    wire [31:0]     _GEN_231; // @[ISA.scala 197:135:@1343.20]
    wire [31:0]     _GEN_232; // @[ISA.scala 197:135:@1343.20]
    wire [31:0]     _GEN_233; // @[ISA.scala 197:135:@1343.20]
    wire [31:0]     _GEN_234; // @[ISA.scala 197:135:@1343.20]
    wire [31:0]     _GEN_235; // @[ISA.scala 197:135:@1343.20]
    wire            _GEN_236; // @[ISA.scala 197:135:@1343.20]
    wire            _GEN_237; // @[ISA.scala 197:135:@1343.20]
    wire            _GEN_238; // @[ISA.scala 197:135:@1343.20]
    wire [2:0]      _GEN_239; // @[ISA.scala 196:127:@1171.18]
    wire [31:0]     _GEN_240; // @[ISA.scala 196:127:@1171.18]
    wire [31:0]     _GEN_241; // @[ISA.scala 196:127:@1171.18]
    wire [31:0]     _GEN_242; // @[ISA.scala 196:127:@1171.18]
    wire [31:0]     _GEN_243; // @[ISA.scala 196:127:@1171.18]
    wire [31:0]     _GEN_244; // @[ISA.scala 196:127:@1171.18]
    wire [31:0]     _GEN_246; // @[ISA.scala 196:127:@1171.18]
    wire [31:0]     _GEN_247; // @[ISA.scala 196:127:@1171.18]
    wire [31:0]     _GEN_248; // @[ISA.scala 196:127:@1171.18]
    wire [31:0]     _GEN_249; // @[ISA.scala 196:127:@1171.18]
    wire [31:0]     _GEN_250; // @[ISA.scala 196:127:@1171.18]
    wire            _GEN_251; // @[ISA.scala 196:127:@1171.18]
    wire            _GEN_252; // @[ISA.scala 196:127:@1171.18]
    wire            _GEN_253; // @[ISA.scala 196:127:@1171.18]
    wire [2:0]      _GEN_254; // @[ISA.scala 195:117:@999.16]
    wire [31:0]     _GEN_255; // @[ISA.scala 195:117:@999.16]
    wire [31:0]     _GEN_256; // @[ISA.scala 195:117:@999.16]
    wire [31:0]     _GEN_257; // @[ISA.scala 195:117:@999.16]
    wire [31:0]     _GEN_258; // @[ISA.scala 195:117:@999.16]
    wire [31:0]     _GEN_259; // @[ISA.scala 195:117:@999.16]
    wire [31:0]     _GEN_261; // @[ISA.scala 195:117:@999.16]
    wire [31:0]     _GEN_262; // @[ISA.scala 195:117:@999.16]
    wire [31:0]     _GEN_263; // @[ISA.scala 195:117:@999.16]
    wire [31:0]     _GEN_264; // @[ISA.scala 195:117:@999.16]
    wire [31:0]     _GEN_265; // @[ISA.scala 195:117:@999.16]
    wire            _GEN_266; // @[ISA.scala 195:117:@999.16]
    wire            _GEN_267; // @[ISA.scala 195:117:@999.16]
    wire            _GEN_268; // @[ISA.scala 195:117:@999.16]
    wire [2:0]      _GEN_269; // @[ISA.scala 194:109:@827.14]
    wire [31:0]     _GEN_270; // @[ISA.scala 194:109:@827.14]
    wire [31:0]     _GEN_271; // @[ISA.scala 194:109:@827.14]
    wire [31:0]     _GEN_272; // @[ISA.scala 194:109:@827.14]
    wire [31:0]     _GEN_273; // @[ISA.scala 194:109:@827.14]
    wire [31:0]     _GEN_274; // @[ISA.scala 194:109:@827.14]
    wire [31:0]     _GEN_276; // @[ISA.scala 194:109:@827.14]
    wire [31:0]     _GEN_277; // @[ISA.scala 194:109:@827.14]
    wire [31:0]     _GEN_278; // @[ISA.scala 194:109:@827.14]
    wire [31:0]     _GEN_279; // @[ISA.scala 194:109:@827.14]
    wire [31:0]     _GEN_280; // @[ISA.scala 194:109:@827.14]
    wire            _GEN_281; // @[ISA.scala 194:109:@827.14]
    wire            _GEN_282; // @[ISA.scala 194:109:@827.14]
    wire            _GEN_283; // @[ISA.scala 194:109:@827.14]
    wire [2:0]      _GEN_284; // @[ISA.scala 193:101:@655.12]
    wire [31:0]     _GEN_285; // @[ISA.scala 193:101:@655.12]
    wire [31:0]     _GEN_286; // @[ISA.scala 193:101:@655.12]
    wire [31:0]     _GEN_287; // @[ISA.scala 193:101:@655.12]
    wire [31:0]     _GEN_288; // @[ISA.scala 193:101:@655.12]
    wire [31:0]     _GEN_289; // @[ISA.scala 193:101:@655.12]
    wire [31:0]     _GEN_291; // @[ISA.scala 193:101:@655.12]
    wire [31:0]     _GEN_292; // @[ISA.scala 193:101:@655.12]
    wire [31:0]     _GEN_293; // @[ISA.scala 193:101:@655.12]
    wire [31:0]     _GEN_294; // @[ISA.scala 193:101:@655.12]
    wire [31:0]     _GEN_295; // @[ISA.scala 193:101:@655.12]
    wire            _GEN_296; // @[ISA.scala 193:101:@655.12]
    wire            _GEN_297; // @[ISA.scala 193:101:@655.12]
    wire            _GEN_298; // @[ISA.scala 193:101:@655.12]
    wire [2:0]      _GEN_299; // @[ISA.scala 192:93:@483.10]
    wire [31:0]     _GEN_300; // @[ISA.scala 192:93:@483.10]
    wire [31:0]     _GEN_301; // @[ISA.scala 192:93:@483.10]
    wire [31:0]     _GEN_302; // @[ISA.scala 192:93:@483.10]
    wire [31:0]     _GEN_303; // @[ISA.scala 192:93:@483.10]
    wire [31:0]     _GEN_304; // @[ISA.scala 192:93:@483.10]
    wire [31:0]     _GEN_306; // @[ISA.scala 192:93:@483.10]
    wire [31:0]     _GEN_307; // @[ISA.scala 192:93:@483.10]
    wire [31:0]     _GEN_308; // @[ISA.scala 192:93:@483.10]
    wire [31:0]     _GEN_309; // @[ISA.scala 192:93:@483.10]
    wire [31:0]     _GEN_310; // @[ISA.scala 192:93:@483.10]
    wire            _GEN_311; // @[ISA.scala 192:93:@483.10]
    wire            _GEN_312; // @[ISA.scala 192:93:@483.10]
    wire            _GEN_313; // @[ISA.scala 192:93:@483.10]
    wire [2:0]      _GEN_314; // @[ISA.scala 191:85:@311.8]
    wire [31:0]     _GEN_315; // @[ISA.scala 191:85:@311.8]
    wire [31:0]     _GEN_316; // @[ISA.scala 191:85:@311.8]
    wire [31:0]     _GEN_317; // @[ISA.scala 191:85:@311.8]
    wire [31:0]     _GEN_318; // @[ISA.scala 191:85:@311.8]
    wire [31:0]     _GEN_319; // @[ISA.scala 191:85:@311.8]
    wire [31:0]     _GEN_321; // @[ISA.scala 191:85:@311.8]
    wire [31:0]     _GEN_322; // @[ISA.scala 191:85:@311.8]
    wire [31:0]     _GEN_323; // @[ISA.scala 191:85:@311.8]
    wire [31:0]     _GEN_324; // @[ISA.scala 191:85:@311.8]
    wire [31:0]     _GEN_325; // @[ISA.scala 191:85:@311.8]
    wire            _GEN_326; // @[ISA.scala 191:85:@311.8]
    wire            _GEN_327; // @[ISA.scala 191:85:@311.8]
    wire            _GEN_328; // @[ISA.scala 191:85:@311.8]
    wire [2:0]      _GEN_329; // @[ISA.scala 190:44:@139.6]
    wire [31:0]     _GEN_330; // @[ISA.scala 190:44:@139.6]
    wire [31:0]     _GEN_331; // @[ISA.scala 190:44:@139.6]
    wire [31:0]     _GEN_332; // @[ISA.scala 190:44:@139.6]
    wire [31:0]     _GEN_333; // @[ISA.scala 190:44:@139.6]
    wire [31:0]     _GEN_334; // @[ISA.scala 190:44:@139.6]
    wire [31:0]     _GEN_336; // @[ISA.scala 190:44:@139.6]
    wire [31:0]     _GEN_337; // @[ISA.scala 190:44:@139.6]
    wire [31:0]     _GEN_338; // @[ISA.scala 190:44:@139.6]
    wire [31:0]     _GEN_339; // @[ISA.scala 190:44:@139.6]
    wire [31:0]     _GEN_340; // @[ISA.scala 190:44:@139.6]
    wire            _GEN_341; // @[ISA.scala 190:44:@139.6]
    wire            _GEN_342; // @[ISA.scala 190:44:@139.6]
    wire            _GEN_343; // @[ISA.scala 190:44:@139.6]
    wire            _T_2303; // @[ISA_functions.scala 452:75:@1731.12]
    wire            _T_2308; // @[ISA_functions.scala 452:125:@1734.12]
    wire            _T_2313; // @[ISA_functions.scala 452:174:@1737.12]
    wire            _T_2318; // @[ISA_functions.scala 452:225:@1740.12]
    wire            _T_2323; // @[ISA_functions.scala 452:275:@1743.12]
    wire            _T_2328; // @[ISA_functions.scala 452:325:@1746.12]
    wire [31:0]     _T_2330; // @[ISA_functions.scala 453:48:@1748.14]
    wire [31:0]     _T_2333; // @[ISA_functions.scala 453:69:@1750.14]
    wire [31:0]     _GEN_352; // @[ISA_functions.scala 452:377:@1747.12]
    wire [31:0]     _T_2342; // @[ISA_functions.scala 286:88:@1760.12]
    wire [31:0]     _T_2345; // @[ISA_functions.scala 286:110:@1762.12]
    wire            _T_2347; // @[ISA_functions.scala 286:123:@1763.12]
    wire            _T_2348; // @[ISA_functions.scala 286:69:@1764.12]
    wire [31:0]     _T_2350; // @[ISA_functions.scala 286:157:@1765.12]
    wire [31:0]     _T_2353; // @[ISA_functions.scala 286:179:@1767.12]
    wire            _T_2355; // @[ISA_functions.scala 286:194:@1768.12]
    wire            _T_2356; // @[ISA_functions.scala 286:138:@1769.12]
    wire            _T_2415; // @[ISA_functions.scala 289:146:@1785.14]
    wire            _T_2416; // @[ISA_functions.scala 289:143:@1786.14]
    wire            _T_2423; // @[ISA_functions.scala 289:271:@1790.14]
    wire            _T_2424; // @[ISA_functions.scala 289:215:@1791.14]
    wire            _T_2455; // @[ISA_functions.scala 292:218:@1813.16]
    wire            _T_2456; // @[ISA_functions.scala 292:215:@1814.16]
    wire            _T_2469; // @[ISA_functions.scala 295:77:@1825.18]
    wire            _T_2470; // @[ISA_functions.scala 295:74:@1826.18]
    wire            _T_2477; // @[ISA_functions.scala 295:198:@1830.18]
    wire            _T_2478; // @[ISA_functions.scala 295:144:@1831.18]
    wire            _T_2501; // @[ISA_functions.scala 298:147:@1848.20]
    wire            _T_2502; // @[ISA_functions.scala 298:144:@1849.20]
    wire            _T_2509; // @[ISA_functions.scala 298:268:@1853.20]
    wire            _T_2510; // @[ISA_functions.scala 298:214:@1854.20]
    wire            _T_2543; // @[ISA_functions.scala 301:217:@1877.22]
    wire            _T_2544; // @[ISA_functions.scala 301:214:@1878.22]
    wire            _T_2551; // @[ISA_functions.scala 301:338:@1882.22]
    wire            _T_2552; // @[ISA_functions.scala 301:284:@1883.22]
    wire            _T_2595; // @[ISA_functions.scala 304:287:@1912.24]
    wire            _T_2596; // @[ISA_functions.scala 304:284:@1913.24]
    wire            _T_2603; // @[ISA_functions.scala 304:408:@1917.24]
    wire            _T_2604; // @[ISA_functions.scala 304:354:@1918.24]
    wire            _T_2657; // @[ISA_functions.scala 307:357:@1953.26]
    wire            _T_2658; // @[ISA_functions.scala 307:354:@1954.26]
    wire            _T_2665; // @[ISA_functions.scala 307:478:@1958.26]
    wire            _T_2666; // @[ISA_functions.scala 307:424:@1959.26]
    wire            _T_2674; // @[ISA_functions.scala 307:493:@1964.26]
    wire            _T_2746; // @[ISA_functions.scala 310:493:@2011.28]
    wire            _T_2754; // @[ISA_functions.scala 310:565:@2016.28]
    wire            _T_2836; // @[ISA_functions.scala 313:565:@2069.30]
    wire            _T_2899; // @[ISA_functions.scala 316:427:@2110.32]
    wire            _T_2900; // @[ISA_functions.scala 316:424:@2111.32]
    wire            _T_2907; // @[ISA_functions.scala 316:548:@2115.32]
    wire            _T_2908; // @[ISA_functions.scala 316:494:@2116.32]
    wire            _T_2981; // @[ISA_functions.scala 319:497:@2163.34]
    wire            _T_2982; // @[ISA_functions.scala 319:494:@2164.34]
    wire            _T_2989; // @[ISA_functions.scala 319:618:@2168.34]
    wire            _T_2990; // @[ISA_functions.scala 319:564:@2169.34]
    wire            _T_3073; // @[ISA_functions.scala 322:567:@2222.36]
    wire            _T_3074; // @[ISA_functions.scala 322:564:@2223.36]
    wire            _T_3093; // @[ISA_functions.scala 325:124:@2238.38]
    wire            _T_3114; // @[ISA_functions.scala 328:124:@2254.40]
    wire            _T_3122; // @[ISA_functions.scala 328:194:@2259.40]
    wire            _T_3153; // @[ISA_functions.scala 331:194:@2281.42]
    wire            _T_3161; // @[ISA_functions.scala 331:264:@2286.42]
    wire            _T_3202; // @[ISA_functions.scala 334:264:@2314.44]
    wire            _T_3210; // @[ISA_functions.scala 334:334:@2319.44]
    wire            _T_3261; // @[ISA_functions.scala 337:334:@2353.46]
    wire            _T_3269; // @[ISA_functions.scala 337:404:@2358.46]
    wire            _T_3330; // @[ISA_functions.scala 340:404:@2398.48]
    wire            _T_3338; // @[ISA_functions.scala 340:474:@2403.48]
    wire            _T_3346; // @[ISA_functions.scala 340:543:@2408.48]
    wire            _T_3425; // @[ISA_functions.scala 343:543:@2459.50]
    wire            _T_3433; // @[ISA_functions.scala 343:615:@2464.50]
    wire            _T_3522; // @[ISA_functions.scala 346:615:@2521.52]
    wire            _T_3593; // @[ISA_functions.scala 349:474:@2567.54]
    wire            _T_3601; // @[ISA_functions.scala 349:544:@2572.54]
    wire            _T_3682; // @[ISA_functions.scala 352:544:@2624.56]
    wire            _T_3690; // @[ISA_functions.scala 352:614:@2629.56]
    wire            _T_3781; // @[ISA_functions.scala 355:614:@2687.58]
    wire            _T_3807; // @[ISA_functions.scala 358:173:@2706.60]
    wire            _T_3835; // @[ISA_functions.scala 361:173:@2726.62]
    wire            _T_3843; // @[ISA_functions.scala 361:243:@2731.62]
    wire            _T_3881; // @[ISA_functions.scala 364:243:@2757.64]
    wire            _T_3889; // @[ISA_functions.scala 364:313:@2762.64]
    wire            _T_3937; // @[ISA_functions.scala 367:313:@2794.66]
    wire            _T_3945; // @[ISA_functions.scala 367:383:@2799.66]
    wire            _T_4003; // @[ISA_functions.scala 370:383:@2837.68]
    wire            _T_4011; // @[ISA_functions.scala 370:453:@2842.68]
    wire            _T_4079; // @[ISA_functions.scala 373:453:@2886.70]
    wire            _T_4144; // @[ISA_functions.scala 379:274:@2931.74]
    wire            _T_4186; // @[ISA_functions.scala 382:274:@2959.76]
    wire            _T_4194; // @[ISA_functions.scala 382:344:@2964.76]
    wire            _T_4246; // @[ISA_functions.scala 385:344:@2998.78]
    wire            _T_4254; // @[ISA_functions.scala 385:414:@3003.78]
    wire            _T_4316; // @[ISA_functions.scala 388:414:@3043.80]
    wire            _T_4363; // @[ISA_functions.scala 391:324:@3074.82]
    wire            _T_4412; // @[ISA_functions.scala 394:324:@3106.84]
    wire            _T_4420; // @[ISA_functions.scala 394:394:@3111.84]
    wire            _T_4479; // @[ISA_functions.scala 397:394:@3149.86]
    wire            _T_4487; // @[ISA_functions.scala 397:464:@3154.86]
    wire            _T_4556; // @[ISA_functions.scala 400:464:@3198.88]
    wire            _T_4564; // @[ISA_functions.scala 400:534:@3203.88]
    wire            _T_4643; // @[ISA_functions.scala 403:534:@3253.90]
    wire            _T_4651; // @[ISA_functions.scala 403:604:@3258.90]
    wire            _T_4740; // @[ISA_functions.scala 406:604:@3314.92]
    wire            _T_4748; // @[ISA_functions.scala 406:674:@3319.92]
    wire            _T_4847; // @[ISA_functions.scala 409:674:@3381.94]
    wire            _T_4893; // @[ISA_functions.scala 412:325:@3411.96]
    wire            _T_4940; // @[ISA_functions.scala 415:328:@3441.98]
    wire            _T_4941; // @[ISA_functions.scala 415:325:@3442.98]
    wire            _T_4946; // @[ISA_functions.scala 415:375:@3445.98]
    wire            _T_5000; // @[ISA_functions.scala 418:378:@3479.100]
    wire            _T_5001; // @[ISA_functions.scala 418:375:@3480.100]
    wire            _T_5006; // @[ISA_functions.scala 418:425:@3483.100]
    wire [31:0]     _GEN_353; // @[ISA_functions.scala 418:476:@3484.100]
    wire [31:0]     _GEN_354; // @[ISA_functions.scala 415:425:@3446.98]
    wire [31:0]     _GEN_355; // @[ISA_functions.scala 412:375:@3412.96]
    wire [31:0]     _GEN_356; // @[ISA_functions.scala 409:745:@3382.94]
    wire [31:0]     _GEN_357; // @[ISA_functions.scala 406:744:@3320.92]
    wire [31:0]     _GEN_358; // @[ISA_functions.scala 403:674:@3259.90]
    wire [31:0]     _GEN_359; // @[ISA_functions.scala 400:604:@3204.88]
    wire [31:0]     _GEN_360; // @[ISA_functions.scala 397:534:@3155.86]
    wire [31:0]     _GEN_361; // @[ISA_functions.scala 394:464:@3112.84]
    wire [31:0]     _GEN_362; // @[ISA_functions.scala 391:394:@3075.82]
    wire [31:0]     _GEN_363; // @[ISA_functions.scala 388:485:@3044.80]
    wire [31:0]     _GEN_364; // @[ISA_functions.scala 385:484:@3004.78]
    wire [31:0]     _GEN_365; // @[ISA_functions.scala 382:414:@2965.76]
    wire [31:0]     _GEN_366; // @[ISA_functions.scala 379:344:@2932.74]
    wire [31:0]     _GEN_367; // @[ISA_functions.scala 376:225:@2905.72]
    wire [31:0]     _GEN_368; // @[ISA_functions.scala 373:524:@2887.70]
    wire [31:0]     _GEN_369; // @[ISA_functions.scala 370:523:@2843.68]
    wire [31:0]     _GEN_370; // @[ISA_functions.scala 367:453:@2800.66]
    wire [31:0]     _GEN_371; // @[ISA_functions.scala 364:383:@2763.64]
    wire [31:0]     _GEN_372; // @[ISA_functions.scala 361:313:@2732.62]
    wire [31:0]     _GEN_373; // @[ISA_functions.scala 358:243:@2707.60]
    wire [31:0]     _GEN_374; // @[ISA_functions.scala 355:685:@2688.58]
    wire [31:0]     _GEN_375; // @[ISA_functions.scala 352:684:@2630.56]
    wire [31:0]     _GEN_376; // @[ISA_functions.scala 349:614:@2573.54]
    wire [31:0]     _GEN_377; // @[ISA_functions.scala 346:689:@2522.52]
    wire [31:0]     _GEN_378; // @[ISA_functions.scala 343:688:@2465.50]
    wire [31:0]     _GEN_379; // @[ISA_functions.scala 340:615:@2409.48]
    wire [31:0]     _GEN_380; // @[ISA_functions.scala 337:474:@2359.46]
    wire [31:0]     _GEN_381; // @[ISA_functions.scala 334:404:@2320.44]
    wire [31:0]     _GEN_382; // @[ISA_functions.scala 331:334:@2287.42]
    wire [31:0]     _GEN_383; // @[ISA_functions.scala 328:264:@2260.40]
    wire [31:0]     _GEN_384; // @[ISA_functions.scala 325:194:@2239.38]
    wire [31:0]     _GEN_385; // @[ISA_functions.scala 322:635:@2224.36]
    wire [31:0]     _GEN_386; // @[ISA_functions.scala 319:634:@2170.34]
    wire [31:0]     _GEN_387; // @[ISA_functions.scala 316:564:@2117.32]
    wire [31:0]     _GEN_388; // @[ISA_functions.scala 313:639:@2070.30]
    wire [31:0]     _GEN_389; // @[ISA_functions.scala 310:638:@2017.28]
    wire [31:0]     _GEN_390; // @[ISA_functions.scala 307:565:@1965.26]
    wire [31:0]     _GEN_391; // @[ISA_functions.scala 304:424:@1919.24]
    wire [31:0]     _GEN_392; // @[ISA_functions.scala 301:354:@1884.22]
    wire [31:0]     _GEN_393; // @[ISA_functions.scala 298:284:@1855.20]
    wire [31:0]     _GEN_394; // @[ISA_functions.scala 295:214:@1832.18]
    wire [31:0]     _GEN_395; // @[ISA_functions.scala 292:289:@1815.16]
    wire [31:0]     _GEN_396; // @[ISA_functions.scala 289:288:@1792.14]
    wire [31:0]     _GEN_397; // @[ISA_functions.scala 286:210:@1770.12]
    wire            _T_5009; // @[ISA_functions.scala 117:40:@3491.12]
    wire            _T_5010; // @[ISA_functions.scala 117:65:@3492.12]
    wire            _T_5011; // @[ISA_functions.scala 117:55:@3493.12]
    wire            _T_5012; // @[ISA_functions.scala 117:92:@3494.12]
    wire            _T_5013; // @[ISA_functions.scala 117:82:@3495.12]
    wire            _T_5014; // @[ISA_functions.scala 117:117:@3496.12]
    wire            _T_5015; // @[ISA_functions.scala 117:107:@3497.12]
    wire            _T_5016; // @[ISA_functions.scala 117:142:@3498.12]
    wire            _T_5017; // @[ISA_functions.scala 117:132:@3499.12]
    wire            _T_5018; // @[ISA_functions.scala 117:167:@3500.12]
    wire            _T_5019; // @[ISA_functions.scala 117:157:@3501.12]
    wire            _T_5020; // @[ISA_functions.scala 117:193:@3502.12]
    wire            _T_5021; // @[ISA_functions.scala 117:183:@3503.12]
    wire            _T_5022; // @[ISA_functions.scala 117:219:@3504.12]
    wire            _T_5023; // @[ISA_functions.scala 117:209:@3505.12]
    wire            _T_5024; // @[ISA_functions.scala 117:244:@3506.12]
    wire            _T_5025; // @[ISA_functions.scala 117:234:@3507.12]
    wire            _T_5026; // @[ISA_functions.scala 117:269:@3508.12]
    wire            _T_5027; // @[ISA_functions.scala 117:259:@3509.12]
    wire            _T_5028; // @[ISA_functions.scala 117:294:@3510.12]
    wire            _T_5029; // @[ISA_functions.scala 117:284:@3511.12]
    wire            _T_5064; // @[ISA_functions.scala 120:28:@3537.14]
    wire            _T_5065; // @[ISA_functions.scala 120:330:@3538.14]
    wire            _T_5066; // @[ISA_functions.scala 120:355:@3539.14]
    wire            _T_5067; // @[ISA_functions.scala 120:345:@3540.14]
    wire            _T_5068; // @[ISA_functions.scala 120:381:@3541.14]
    wire            _T_5069; // @[ISA_functions.scala 120:371:@3542.14]
    wire            _T_5070; // @[ISA_functions.scala 120:318:@3543.14]
    wire            _T_5100; // @[ISA_functions.scala 123:321:@3575.16]
    wire            _T_5101; // @[ISA_functions.scala 123:318:@3576.16]
    wire            _T_5102; // @[ISA_functions.scala 123:409:@3577.16]
    wire            _T_5103; // @[ISA_functions.scala 123:434:@3578.16]
    wire            _T_5104; // @[ISA_functions.scala 123:424:@3579.16]
    wire            _T_5105; // @[ISA_functions.scala 123:398:@3580.16]
    wire            _T_5141; // @[ISA_functions.scala 126:401:@3617.18]
    wire            _T_5142; // @[ISA_functions.scala 126:398:@3618.18]
    wire            _T_5143; // @[ISA_functions.scala 126:465:@3619.18]
    wire            _T_5144; // @[ISA_functions.scala 126:490:@3620.18]
    wire            _T_5145; // @[ISA_functions.scala 126:480:@3621.18]
    wire            _T_5146; // @[ISA_functions.scala 126:517:@3622.18]
    wire            _T_5147; // @[ISA_functions.scala 126:507:@3623.18]
    wire            _T_5148; // @[ISA_functions.scala 126:543:@3624.18]
    wire            _T_5149; // @[ISA_functions.scala 126:533:@3625.18]
    wire            _T_5150; // @[ISA_functions.scala 126:452:@3626.18]
    wire            _T_5196; // @[ISA_functions.scala 129:455:@3672.20]
    wire            _T_5197; // @[ISA_functions.scala 129:452:@3673.20]
    wire            _T_5198; // @[ISA_functions.scala 129:573:@3674.20]
    wire            _T_5199; // @[ISA_functions.scala 129:599:@3675.20]
    wire            _T_5200; // @[ISA_functions.scala 129:589:@3676.20]
    wire            _T_5201; // @[ISA_functions.scala 129:627:@3677.20]
    wire            _T_5202; // @[ISA_functions.scala 129:617:@3678.20]
    wire            _T_5203; // @[ISA_functions.scala 129:654:@3679.20]
    wire            _T_5204; // @[ISA_functions.scala 129:644:@3680.20]
    wire            _T_5205; // @[ISA_functions.scala 129:560:@3681.20]
    wire            _T_5261; // @[ISA_functions.scala 132:563:@3736.22]
    wire            _T_5262; // @[ISA_functions.scala 132:560:@3737.22]
    wire            _T_5263; // @[ISA_functions.scala 132:683:@3738.22]
    wire            _T_5264; // @[ISA_functions.scala 132:708:@3739.22]
    wire            _T_5265; // @[ISA_functions.scala 132:698:@3740.22]
    wire            _T_5266; // @[ISA_functions.scala 132:672:@3741.22]
    wire            _T_5328; // @[ISA_functions.scala 135:675:@3801.24]
    wire            _T_5329; // @[ISA_functions.scala 135:672:@3802.24]
    wire            _T_5330; // @[ISA_functions.scala 135:737:@3803.24]
    wire            _T_5331; // @[ISA_functions.scala 135:762:@3804.24]
    wire            _T_5332; // @[ISA_functions.scala 135:752:@3805.24]
    wire            _T_5333; // @[ISA_functions.scala 135:726:@3806.24]
    wire            _T_5401; // @[ISA_functions.scala 138:729:@3871.26]
    wire            _T_5402; // @[ISA_functions.scala 138:726:@3872.26]
    wire            _T_5403; // @[ISA_functions.scala 138:791:@3873.26]
    wire            _T_5404; // @[ISA_functions.scala 138:816:@3874.26]
    wire            _T_5405; // @[ISA_functions.scala 138:806:@3875.26]
    wire            _T_5406; // @[ISA_functions.scala 138:780:@3876.26]
    wire            _T_5480; // @[ISA_functions.scala 141:783:@3946.28]
    wire            _T_5481; // @[ISA_functions.scala 141:780:@3947.28]
    wire            _T_5482; // @[ISA_functions.scala 141:845:@3948.28]
    wire            _T_5483; // @[ISA_functions.scala 141:869:@3949.28]
    wire            _T_5484; // @[ISA_functions.scala 141:859:@3950.28]
    wire            _T_5485; // @[ISA_functions.scala 141:834:@3951.28]
    wire            _T_5565; // @[ISA_functions.scala 144:837:@4026.30]
    wire            _T_5566; // @[ISA_functions.scala 144:834:@4027.30]
    wire            _T_5567; // @[ISA_functions.scala 144:897:@4028.30]
    wire            _T_5568; // @[ISA_functions.scala 144:922:@4029.30]
    wire            _T_5569; // @[ISA_functions.scala 144:912:@4030.30]
    wire            _T_5570; // @[ISA_functions.scala 144:886:@4031.30]
    wire            _T_5656; // @[ISA_functions.scala 147:889:@4111.32]
    wire            _T_5657; // @[ISA_functions.scala 147:886:@4112.32]
    wire            _T_5658; // @[ISA_functions.scala 147:951:@4113.32]
    wire            _T_5659; // @[ISA_functions.scala 147:977:@4114.32]
    wire            _T_5660; // @[ISA_functions.scala 147:967:@4115.32]
    wire            _T_5661; // @[ISA_functions.scala 147:940:@4116.32]
    wire            _T_5753; // @[ISA_functions.scala 150:943:@4201.34]
    wire            _T_5754; // @[ISA_functions.scala 150:940:@4202.34]
    wire            _T_5755; // @[ISA_functions.scala 150:1004:@4203.34]
    wire            _T_5756; // @[ISA_functions.scala 150:994:@4204.34]
    wire [31:0]     _GEN_398; // @[ISA_functions.scala 150:1020:@4205.34]
    wire [31:0]     _GEN_399; // @[ISA_functions.scala 147:994:@4117.32]
    wire [31:0]     _GEN_400; // @[ISA_functions.scala 144:940:@4032.30]
    wire [31:0]     _GEN_401; // @[ISA_functions.scala 141:886:@3952.28]
    wire [31:0]     _GEN_402; // @[ISA_functions.scala 138:834:@3877.26]
    wire [31:0]     _GEN_403; // @[ISA_functions.scala 135:780:@3807.24]
    wire [31:0]     _GEN_404; // @[ISA_functions.scala 132:726:@3742.22]
    wire [31:0]     _GEN_405; // @[ISA_functions.scala 129:672:@3682.20]
    wire [31:0]     _GEN_406; // @[ISA_functions.scala 126:560:@3627.18]
    wire [31:0]     _GEN_407; // @[ISA_functions.scala 123:452:@3581.16]
    wire [31:0]     _GEN_408; // @[ISA_functions.scala 120:398:@3544.14]
    wire [31:0]     _GEN_409; // @[ISA_functions.scala 117:313:@3512.12]
    wire            _T_5782; // @[ISA_functions.scala 463:224:@4225.12]
    wire            _T_5787; // @[ISA_functions.scala 463:274:@4228.12]
    wire [31:0]     _T_5789; // @[ISA_functions.scala 464:48:@4230.14]
    wire [31:0]     _T_5792; // @[ISA_functions.scala 464:70:@4232.14]
    wire [31:0]     _GEN_410; // @[ISA_functions.scala 463:325:@4229.12]
    wire            _T_5797; // @[ISA_functions.scala 485:28:@4239.12]
    wire            _T_5802; // @[ISA_functions.scala 488:28:@4245.14]
    wire            _T_5804; // @[ISA_functions.scala 488:57:@4246.14]
    wire            _T_5805; // @[ISA_functions.scala 488:49:@4247.14]
    wire            _T_5813; // @[ISA_functions.scala 491:52:@4255.16]
    wire            _T_5814; // @[ISA_functions.scala 491:49:@4256.16]
    wire            _T_5816; // @[ISA_functions.scala 491:81:@4257.16]
    wire            _T_5817; // @[ISA_functions.scala 491:73:@4258.16]
    wire            _T_5830; // @[ISA_functions.scala 494:76:@4269.18]
    wire            _T_5831; // @[ISA_functions.scala 494:73:@4270.18]
    wire            _T_5833; // @[ISA_functions.scala 494:105:@4271.18]
    wire            _T_5834; // @[ISA_functions.scala 494:97:@4272.18]
    wire            _T_5852; // @[ISA_functions.scala 497:100:@4286.20]
    wire            _T_5853; // @[ISA_functions.scala 497:97:@4287.20]
    wire            _T_5855; // @[ISA_functions.scala 497:129:@4288.20]
    wire            _T_5856; // @[ISA_functions.scala 497:121:@4289.20]
    wire            _T_5879; // @[ISA_functions.scala 500:124:@4306.22]
    wire            _T_5880; // @[ISA_functions.scala 500:121:@4307.22]
    wire            _T_5882; // @[ISA_functions.scala 500:153:@4308.22]
    wire            _T_5883; // @[ISA_functions.scala 500:145:@4309.22]
    wire            _T_5911; // @[ISA_functions.scala 503:148:@4329.24]
    wire            _T_5912; // @[ISA_functions.scala 503:145:@4330.24]
    wire            _T_5914; // @[ISA_functions.scala 503:177:@4331.24]
    wire            _T_5915; // @[ISA_functions.scala 503:169:@4332.24]
    wire            _T_5948; // @[ISA_functions.scala 506:172:@4355.26]
    wire            _T_5949; // @[ISA_functions.scala 506:169:@4356.26]
    wire            _T_5951; // @[ISA_functions.scala 506:201:@4357.26]
    wire            _T_5952; // @[ISA_functions.scala 506:193:@4358.26]
    wire            _T_5990; // @[ISA_functions.scala 509:196:@4384.28]
    wire            _T_5991; // @[ISA_functions.scala 509:193:@4385.28]
    wire            _T_5993; // @[ISA_functions.scala 509:225:@4386.28]
    wire            _T_5994; // @[ISA_functions.scala 509:217:@4387.28]
    wire            _T_6037; // @[ISA_functions.scala 512:220:@4416.30]
    wire            _T_6038; // @[ISA_functions.scala 512:217:@4417.30]
    wire            _T_6040; // @[ISA_functions.scala 512:249:@4418.30]
    wire            _T_6041; // @[ISA_functions.scala 512:241:@4419.30]
    wire            _T_6089; // @[ISA_functions.scala 515:244:@4451.32]
    wire            _T_6090; // @[ISA_functions.scala 515:241:@4452.32]
    wire            _T_6092; // @[ISA_functions.scala 515:273:@4453.32]
    wire            _T_6093; // @[ISA_functions.scala 515:265:@4454.32]
    wire            _T_6146; // @[ISA_functions.scala 518:268:@4489.34]
    wire            _T_6147; // @[ISA_functions.scala 518:265:@4490.34]
    wire            _T_6149; // @[ISA_functions.scala 518:298:@4491.34]
    wire            _T_6150; // @[ISA_functions.scala 518:290:@4492.34]
    wire            _T_6208; // @[ISA_functions.scala 521:293:@4530.36]
    wire            _T_6209; // @[ISA_functions.scala 521:290:@4531.36]
    wire            _T_6211; // @[ISA_functions.scala 521:323:@4532.36]
    wire            _T_6212; // @[ISA_functions.scala 521:315:@4533.36]
    wire            _T_6275; // @[ISA_functions.scala 524:318:@4574.38]
    wire            _T_6276; // @[ISA_functions.scala 524:315:@4575.38]
    wire            _T_6278; // @[ISA_functions.scala 524:348:@4576.38]
    wire            _T_6279; // @[ISA_functions.scala 524:340:@4577.38]
    wire            _T_6347; // @[ISA_functions.scala 527:343:@4621.40]
    wire            _T_6348; // @[ISA_functions.scala 527:340:@4622.40]
    wire            _T_6350; // @[ISA_functions.scala 527:373:@4623.40]
    wire            _T_6351; // @[ISA_functions.scala 527:365:@4624.40]
    wire            _T_6424; // @[ISA_functions.scala 530:368:@4671.42]
    wire            _T_6425; // @[ISA_functions.scala 530:365:@4672.42]
    wire            _T_6427; // @[ISA_functions.scala 530:398:@4673.42]
    wire            _T_6428; // @[ISA_functions.scala 530:390:@4674.42]
    wire            _T_6506; // @[ISA_functions.scala 533:393:@4724.44]
    wire            _T_6507; // @[ISA_functions.scala 533:390:@4725.44]
    wire            _T_6509; // @[ISA_functions.scala 533:423:@4726.44]
    wire            _T_6510; // @[ISA_functions.scala 533:415:@4727.44]
    wire            _T_6593; // @[ISA_functions.scala 536:418:@4780.46]
    wire            _T_6594; // @[ISA_functions.scala 536:415:@4781.46]
    wire            _T_6596; // @[ISA_functions.scala 536:448:@4782.46]
    wire            _T_6597; // @[ISA_functions.scala 536:440:@4783.46]
    wire            _T_6685; // @[ISA_functions.scala 539:443:@4839.48]
    wire            _T_6686; // @[ISA_functions.scala 539:440:@4840.48]
    wire            _T_6688; // @[ISA_functions.scala 539:473:@4841.48]
    wire            _T_6689; // @[ISA_functions.scala 539:465:@4842.48]
    wire            _T_6782; // @[ISA_functions.scala 542:468:@4901.50]
    wire            _T_6783; // @[ISA_functions.scala 542:465:@4902.50]
    wire            _T_6785; // @[ISA_functions.scala 542:498:@4903.50]
    wire            _T_6786; // @[ISA_functions.scala 542:490:@4904.50]
    wire            _T_6884; // @[ISA_functions.scala 545:493:@4966.52]
    wire            _T_6885; // @[ISA_functions.scala 545:490:@4967.52]
    wire            _T_6887; // @[ISA_functions.scala 545:523:@4968.52]
    wire            _T_6888; // @[ISA_functions.scala 545:515:@4969.52]
    wire            _T_6991; // @[ISA_functions.scala 548:518:@5034.54]
    wire            _T_6992; // @[ISA_functions.scala 548:515:@5035.54]
    wire            _T_6994; // @[ISA_functions.scala 548:548:@5036.54]
    wire            _T_6995; // @[ISA_functions.scala 548:540:@5037.54]
    wire            _T_7103; // @[ISA_functions.scala 551:543:@5105.56]
    wire            _T_7104; // @[ISA_functions.scala 551:540:@5106.56]
    wire            _T_7106; // @[ISA_functions.scala 551:573:@5107.56]
    wire            _T_7107; // @[ISA_functions.scala 551:565:@5108.56]
    wire            _T_7220; // @[ISA_functions.scala 554:568:@5179.58]
    wire            _T_7221; // @[ISA_functions.scala 554:565:@5180.58]
    wire            _T_7223; // @[ISA_functions.scala 554:598:@5181.58]
    wire            _T_7224; // @[ISA_functions.scala 554:590:@5182.58]
    wire            _T_7342; // @[ISA_functions.scala 557:593:@5256.60]
    wire            _T_7343; // @[ISA_functions.scala 557:590:@5257.60]
    wire            _T_7345; // @[ISA_functions.scala 557:623:@5258.60]
    wire            _T_7346; // @[ISA_functions.scala 557:615:@5259.60]
    wire            _T_7469; // @[ISA_functions.scala 560:618:@5336.62]
    wire            _T_7470; // @[ISA_functions.scala 560:615:@5337.62]
    wire            _T_7472; // @[ISA_functions.scala 560:648:@5338.62]
    wire            _T_7473; // @[ISA_functions.scala 560:640:@5339.62]
    wire            _T_7601; // @[ISA_functions.scala 563:643:@5419.64]
    wire            _T_7602; // @[ISA_functions.scala 563:640:@5420.64]
    wire            _T_7604; // @[ISA_functions.scala 563:673:@5421.64]
    wire            _T_7605; // @[ISA_functions.scala 563:665:@5422.64]
    wire            _T_7738; // @[ISA_functions.scala 566:668:@5505.66]
    wire            _T_7739; // @[ISA_functions.scala 566:665:@5506.66]
    wire            _T_7741; // @[ISA_functions.scala 566:698:@5507.66]
    wire            _T_7742; // @[ISA_functions.scala 566:690:@5508.66]
    wire            _T_7880; // @[ISA_functions.scala 569:693:@5594.68]
    wire            _T_7881; // @[ISA_functions.scala 569:690:@5595.68]
    wire            _T_7883; // @[ISA_functions.scala 569:723:@5596.68]
    wire            _T_7884; // @[ISA_functions.scala 569:715:@5597.68]
    wire            _T_8027; // @[ISA_functions.scala 572:718:@5686.70]
    wire            _T_8028; // @[ISA_functions.scala 572:715:@5687.70]
    wire            _T_8030; // @[ISA_functions.scala 572:748:@5688.70]
    wire            _T_8031; // @[ISA_functions.scala 572:740:@5689.70]
    wire            _T_8179; // @[ISA_functions.scala 575:743:@5781.72]
    wire            _T_8180; // @[ISA_functions.scala 575:740:@5782.72]
    wire            _T_8182; // @[ISA_functions.scala 575:773:@5783.72]
    wire            _T_8183; // @[ISA_functions.scala 575:765:@5784.72]
    wire [31:0]     _GEN_411; // @[ISA_functions.scala 575:790:@5785.72]
    wire [31:0]     _GEN_412; // @[ISA_functions.scala 572:765:@5690.70]
    wire [31:0]     _GEN_413; // @[ISA_functions.scala 569:740:@5598.68]
    wire [31:0]     _GEN_414; // @[ISA_functions.scala 566:715:@5509.66]
    wire [31:0]     _GEN_415; // @[ISA_functions.scala 563:690:@5423.64]
    wire [31:0]     _GEN_416; // @[ISA_functions.scala 560:665:@5340.62]
    wire [31:0]     _GEN_417; // @[ISA_functions.scala 557:640:@5260.60]
    wire [31:0]     _GEN_418; // @[ISA_functions.scala 554:615:@5183.58]
    wire [31:0]     _GEN_419; // @[ISA_functions.scala 551:590:@5109.56]
    wire [31:0]     _GEN_420; // @[ISA_functions.scala 548:565:@5038.54]
    wire [31:0]     _GEN_421; // @[ISA_functions.scala 545:540:@4970.52]
    wire [31:0]     _GEN_422; // @[ISA_functions.scala 542:515:@4905.50]
    wire [31:0]     _GEN_423; // @[ISA_functions.scala 539:490:@4843.48]
    wire [31:0]     _GEN_424; // @[ISA_functions.scala 536:465:@4784.46]
    wire [31:0]     _GEN_425; // @[ISA_functions.scala 533:440:@4728.44]
    wire [31:0]     _GEN_426; // @[ISA_functions.scala 530:415:@4675.42]
    wire [31:0]     _GEN_427; // @[ISA_functions.scala 527:390:@4625.40]
    wire [31:0]     _GEN_428; // @[ISA_functions.scala 524:365:@4578.38]
    wire [31:0]     _GEN_429; // @[ISA_functions.scala 521:340:@4534.36]
    wire [31:0]     _GEN_430; // @[ISA_functions.scala 518:315:@4493.34]
    wire [31:0]     _GEN_431; // @[ISA_functions.scala 515:290:@4455.32]
    wire [31:0]     _GEN_432; // @[ISA_functions.scala 512:265:@4420.30]
    wire [31:0]     _GEN_433; // @[ISA_functions.scala 509:241:@4388.28]
    wire [31:0]     _GEN_434; // @[ISA_functions.scala 506:217:@4359.26]
    wire [31:0]     _GEN_435; // @[ISA_functions.scala 503:193:@4333.24]
    wire [31:0]     _GEN_436; // @[ISA_functions.scala 500:169:@4310.22]
    wire [31:0]     _GEN_437; // @[ISA_functions.scala 497:145:@4290.20]
    wire [31:0]     _GEN_438; // @[ISA_functions.scala 494:121:@4273.18]
    wire [31:0]     _GEN_439; // @[ISA_functions.scala 491:97:@4259.16]
    wire [31:0]     _GEN_440; // @[ISA_functions.scala 488:73:@4248.14]
    wire [31:0]     _GEN_441; // @[ISA_functions.scala 485:44:@4240.12]
    wire            _T_8194; // @[ISA_functions.scala 474:71:@5796.12]
    wire            _T_8199; // @[ISA_functions.scala 474:121:@5799.12]
    wire [31:0]     _T_8201; // @[ISA_functions.scala 475:48:@5801.14]
    wire [31:0]     _T_8204; // @[ISA_functions.scala 475:70:@5803.14]
    wire [31:0]     _GEN_442; // @[ISA_functions.scala 474:172:@5800.12]
    wire            _T_8209; // @[ISA_functions.scala 485:28:@5810.12]
    wire            _T_8214; // @[ISA_functions.scala 488:28:@5816.14]
    wire            _T_8216; // @[ISA_functions.scala 488:57:@5817.14]
    wire            _T_8217; // @[ISA_functions.scala 488:49:@5818.14]
    wire            _T_8225; // @[ISA_functions.scala 491:52:@5826.16]
    wire            _T_8226; // @[ISA_functions.scala 491:49:@5827.16]
    wire            _T_8228; // @[ISA_functions.scala 491:81:@5828.16]
    wire            _T_8229; // @[ISA_functions.scala 491:73:@5829.16]
    wire            _T_8242; // @[ISA_functions.scala 494:76:@5840.18]
    wire            _T_8243; // @[ISA_functions.scala 494:73:@5841.18]
    wire            _T_8245; // @[ISA_functions.scala 494:105:@5842.18]
    wire            _T_8246; // @[ISA_functions.scala 494:97:@5843.18]
    wire            _T_8264; // @[ISA_functions.scala 497:100:@5857.20]
    wire            _T_8265; // @[ISA_functions.scala 497:97:@5858.20]
    wire            _T_8267; // @[ISA_functions.scala 497:129:@5859.20]
    wire            _T_8268; // @[ISA_functions.scala 497:121:@5860.20]
    wire            _T_8291; // @[ISA_functions.scala 500:124:@5877.22]
    wire            _T_8292; // @[ISA_functions.scala 500:121:@5878.22]
    wire            _T_8294; // @[ISA_functions.scala 500:153:@5879.22]
    wire            _T_8295; // @[ISA_functions.scala 500:145:@5880.22]
    wire            _T_8323; // @[ISA_functions.scala 503:148:@5900.24]
    wire            _T_8324; // @[ISA_functions.scala 503:145:@5901.24]
    wire            _T_8326; // @[ISA_functions.scala 503:177:@5902.24]
    wire            _T_8327; // @[ISA_functions.scala 503:169:@5903.24]
    wire            _T_8360; // @[ISA_functions.scala 506:172:@5926.26]
    wire            _T_8361; // @[ISA_functions.scala 506:169:@5927.26]
    wire            _T_8363; // @[ISA_functions.scala 506:201:@5928.26]
    wire            _T_8364; // @[ISA_functions.scala 506:193:@5929.26]
    wire            _T_8402; // @[ISA_functions.scala 509:196:@5955.28]
    wire            _T_8403; // @[ISA_functions.scala 509:193:@5956.28]
    wire            _T_8405; // @[ISA_functions.scala 509:225:@5957.28]
    wire            _T_8406; // @[ISA_functions.scala 509:217:@5958.28]
    wire            _T_8449; // @[ISA_functions.scala 512:220:@5987.30]
    wire            _T_8450; // @[ISA_functions.scala 512:217:@5988.30]
    wire            _T_8452; // @[ISA_functions.scala 512:249:@5989.30]
    wire            _T_8453; // @[ISA_functions.scala 512:241:@5990.30]
    wire            _T_8501; // @[ISA_functions.scala 515:244:@6022.32]
    wire            _T_8502; // @[ISA_functions.scala 515:241:@6023.32]
    wire            _T_8504; // @[ISA_functions.scala 515:273:@6024.32]
    wire            _T_8505; // @[ISA_functions.scala 515:265:@6025.32]
    wire            _T_8558; // @[ISA_functions.scala 518:268:@6060.34]
    wire            _T_8559; // @[ISA_functions.scala 518:265:@6061.34]
    wire            _T_8561; // @[ISA_functions.scala 518:298:@6062.34]
    wire            _T_8562; // @[ISA_functions.scala 518:290:@6063.34]
    wire            _T_8620; // @[ISA_functions.scala 521:293:@6101.36]
    wire            _T_8621; // @[ISA_functions.scala 521:290:@6102.36]
    wire            _T_8623; // @[ISA_functions.scala 521:323:@6103.36]
    wire            _T_8624; // @[ISA_functions.scala 521:315:@6104.36]
    wire            _T_8687; // @[ISA_functions.scala 524:318:@6145.38]
    wire            _T_8688; // @[ISA_functions.scala 524:315:@6146.38]
    wire            _T_8690; // @[ISA_functions.scala 524:348:@6147.38]
    wire            _T_8691; // @[ISA_functions.scala 524:340:@6148.38]
    wire            _T_8759; // @[ISA_functions.scala 527:343:@6192.40]
    wire            _T_8760; // @[ISA_functions.scala 527:340:@6193.40]
    wire            _T_8762; // @[ISA_functions.scala 527:373:@6194.40]
    wire            _T_8763; // @[ISA_functions.scala 527:365:@6195.40]
    wire            _T_8836; // @[ISA_functions.scala 530:368:@6242.42]
    wire            _T_8837; // @[ISA_functions.scala 530:365:@6243.42]
    wire            _T_8839; // @[ISA_functions.scala 530:398:@6244.42]
    wire            _T_8840; // @[ISA_functions.scala 530:390:@6245.42]
    wire            _T_8918; // @[ISA_functions.scala 533:393:@6295.44]
    wire            _T_8919; // @[ISA_functions.scala 533:390:@6296.44]
    wire            _T_8921; // @[ISA_functions.scala 533:423:@6297.44]
    wire            _T_8922; // @[ISA_functions.scala 533:415:@6298.44]
    wire            _T_9005; // @[ISA_functions.scala 536:418:@6351.46]
    wire            _T_9006; // @[ISA_functions.scala 536:415:@6352.46]
    wire            _T_9008; // @[ISA_functions.scala 536:448:@6353.46]
    wire            _T_9009; // @[ISA_functions.scala 536:440:@6354.46]
    wire            _T_9097; // @[ISA_functions.scala 539:443:@6410.48]
    wire            _T_9098; // @[ISA_functions.scala 539:440:@6411.48]
    wire            _T_9100; // @[ISA_functions.scala 539:473:@6412.48]
    wire            _T_9101; // @[ISA_functions.scala 539:465:@6413.48]
    wire            _T_9194; // @[ISA_functions.scala 542:468:@6472.50]
    wire            _T_9195; // @[ISA_functions.scala 542:465:@6473.50]
    wire            _T_9197; // @[ISA_functions.scala 542:498:@6474.50]
    wire            _T_9198; // @[ISA_functions.scala 542:490:@6475.50]
    wire            _T_9296; // @[ISA_functions.scala 545:493:@6537.52]
    wire            _T_9297; // @[ISA_functions.scala 545:490:@6538.52]
    wire            _T_9299; // @[ISA_functions.scala 545:523:@6539.52]
    wire            _T_9300; // @[ISA_functions.scala 545:515:@6540.52]
    wire            _T_9403; // @[ISA_functions.scala 548:518:@6605.54]
    wire            _T_9404; // @[ISA_functions.scala 548:515:@6606.54]
    wire            _T_9406; // @[ISA_functions.scala 548:548:@6607.54]
    wire            _T_9407; // @[ISA_functions.scala 548:540:@6608.54]
    wire            _T_9515; // @[ISA_functions.scala 551:543:@6676.56]
    wire            _T_9516; // @[ISA_functions.scala 551:540:@6677.56]
    wire            _T_9518; // @[ISA_functions.scala 551:573:@6678.56]
    wire            _T_9519; // @[ISA_functions.scala 551:565:@6679.56]
    wire            _T_9632; // @[ISA_functions.scala 554:568:@6750.58]
    wire            _T_9633; // @[ISA_functions.scala 554:565:@6751.58]
    wire            _T_9635; // @[ISA_functions.scala 554:598:@6752.58]
    wire            _T_9636; // @[ISA_functions.scala 554:590:@6753.58]
    wire            _T_9754; // @[ISA_functions.scala 557:593:@6827.60]
    wire            _T_9755; // @[ISA_functions.scala 557:590:@6828.60]
    wire            _T_9757; // @[ISA_functions.scala 557:623:@6829.60]
    wire            _T_9758; // @[ISA_functions.scala 557:615:@6830.60]
    wire            _T_9881; // @[ISA_functions.scala 560:618:@6907.62]
    wire            _T_9882; // @[ISA_functions.scala 560:615:@6908.62]
    wire            _T_9884; // @[ISA_functions.scala 560:648:@6909.62]
    wire            _T_9885; // @[ISA_functions.scala 560:640:@6910.62]
    wire            _T_10013; // @[ISA_functions.scala 563:643:@6990.64]
    wire            _T_10014; // @[ISA_functions.scala 563:640:@6991.64]
    wire            _T_10016; // @[ISA_functions.scala 563:673:@6992.64]
    wire            _T_10017; // @[ISA_functions.scala 563:665:@6993.64]
    wire            _T_10150; // @[ISA_functions.scala 566:668:@7076.66]
    wire            _T_10151; // @[ISA_functions.scala 566:665:@7077.66]
    wire            _T_10153; // @[ISA_functions.scala 566:698:@7078.66]
    wire            _T_10154; // @[ISA_functions.scala 566:690:@7079.66]
    wire            _T_10292; // @[ISA_functions.scala 569:693:@7165.68]
    wire            _T_10293; // @[ISA_functions.scala 569:690:@7166.68]
    wire            _T_10295; // @[ISA_functions.scala 569:723:@7167.68]
    wire            _T_10296; // @[ISA_functions.scala 569:715:@7168.68]
    wire            _T_10439; // @[ISA_functions.scala 572:718:@7257.70]
    wire            _T_10440; // @[ISA_functions.scala 572:715:@7258.70]
    wire            _T_10442; // @[ISA_functions.scala 572:748:@7259.70]
    wire            _T_10443; // @[ISA_functions.scala 572:740:@7260.70]
    wire            _T_10591; // @[ISA_functions.scala 575:743:@7352.72]
    wire            _T_10592; // @[ISA_functions.scala 575:740:@7353.72]
    wire            _T_10594; // @[ISA_functions.scala 575:773:@7354.72]
    wire            _T_10595; // @[ISA_functions.scala 575:765:@7355.72]
    wire [31:0]     _GEN_443; // @[ISA_functions.scala 575:790:@7356.72]
    wire [31:0]     _GEN_444; // @[ISA_functions.scala 572:765:@7261.70]
    wire [31:0]     _GEN_445; // @[ISA_functions.scala 569:740:@7169.68]
    wire [31:0]     _GEN_446; // @[ISA_functions.scala 566:715:@7080.66]
    wire [31:0]     _GEN_447; // @[ISA_functions.scala 563:690:@6994.64]
    wire [31:0]     _GEN_448; // @[ISA_functions.scala 560:665:@6911.62]
    wire [31:0]     _GEN_449; // @[ISA_functions.scala 557:640:@6831.60]
    wire [31:0]     _GEN_450; // @[ISA_functions.scala 554:615:@6754.58]
    wire [31:0]     _GEN_451; // @[ISA_functions.scala 551:590:@6680.56]
    wire [31:0]     _GEN_452; // @[ISA_functions.scala 548:565:@6609.54]
    wire [31:0]     _GEN_453; // @[ISA_functions.scala 545:540:@6541.52]
    wire [31:0]     _GEN_454; // @[ISA_functions.scala 542:515:@6476.50]
    wire [31:0]     _GEN_455; // @[ISA_functions.scala 539:490:@6414.48]
    wire [31:0]     _GEN_456; // @[ISA_functions.scala 536:465:@6355.46]
    wire [31:0]     _GEN_457; // @[ISA_functions.scala 533:440:@6299.44]
    wire [31:0]     _GEN_458; // @[ISA_functions.scala 530:415:@6246.42]
    wire [31:0]     _GEN_459; // @[ISA_functions.scala 527:390:@6196.40]
    wire [31:0]     _GEN_460; // @[ISA_functions.scala 524:365:@6149.38]
    wire [31:0]     _GEN_461; // @[ISA_functions.scala 521:340:@6105.36]
    wire [31:0]     _GEN_462; // @[ISA_functions.scala 518:315:@6064.34]
    wire [31:0]     _GEN_463; // @[ISA_functions.scala 515:290:@6026.32]
    wire [31:0]     _GEN_464; // @[ISA_functions.scala 512:265:@5991.30]
    wire [31:0]     _GEN_465; // @[ISA_functions.scala 509:241:@5959.28]
    wire [31:0]     _GEN_466; // @[ISA_functions.scala 506:217:@5930.26]
    wire [31:0]     _GEN_467; // @[ISA_functions.scala 503:193:@5904.24]
    wire [31:0]     _GEN_468; // @[ISA_functions.scala 500:169:@5881.22]
    wire [31:0]     _GEN_469; // @[ISA_functions.scala 497:145:@5861.20]
    wire [31:0]     _GEN_470; // @[ISA_functions.scala 494:121:@5844.18]
    wire [31:0]     _GEN_471; // @[ISA_functions.scala 491:97:@5830.16]
    wire [31:0]     _GEN_472; // @[ISA_functions.scala 488:73:@5819.14]
    wire [31:0]     _GEN_473; // @[ISA_functions.scala 485:44:@5811.12]
    wire            _T_10598; // @[ISA_functions.scala 161:36:@7363.12]
    wire [32:0]     _T_10599; // @[ISA_functions.scala 162:43:@7365.14]
    wire [31:0]     _T_10600; // @[ISA_functions.scala 162:43:@7366.14]
    wire            _T_10603; // @[ISA_functions.scala 164:28:@7371.14]
    wire            _T_10604; // @[ISA_functions.scala 164:71:@7372.14]
    wire            _T_10605; // @[ISA_functions.scala 164:55:@7373.14]
    wire [63:0]     _T_10607; // @[ISA_functions.scala 165:55:@7375.16]
    wire [63:0]     _GEN_6225; // @[ISA_functions.scala 165:43:@7376.16]
    wire [64:0]     _T_10608; // @[ISA_functions.scala 165:43:@7376.16]
    wire [63:0]     _T_10609; // @[ISA_functions.scala 165:43:@7377.16]
    wire            _T_10615; // @[ISA_functions.scala 167:58:@7384.16]
    wire            _T_10616; // @[ISA_functions.scala 167:55:@7385.16]
    wire            _T_10617; // @[ISA_functions.scala 167:101:@7386.16]
    wire            _T_10618; // @[ISA_functions.scala 167:85:@7387.16]
    wire [31:0]     _T_10619; // @[ISA_functions.scala 168:43:@7389.18]
    wire            _T_10629; // @[ISA_functions.scala 170:88:@7399.18]
    wire            _T_10630; // @[ISA_functions.scala 170:85:@7400.18]
    wire            _T_10631; // @[ISA_functions.scala 170:131:@7401.18]
    wire            _T_10632; // @[ISA_functions.scala 170:115:@7402.18]
    wire [31:0]     _T_10633; // @[ISA_functions.scala 171:43:@7404.20]
    wire            _T_10647; // @[ISA_functions.scala 173:118:@7417.20]
    wire            _T_10648; // @[ISA_functions.scala 173:115:@7418.20]
    wire            _T_10649; // @[ISA_functions.scala 173:160:@7419.20]
    wire            _T_10650; // @[ISA_functions.scala 173:144:@7420.20]
    wire [31:0]     _T_10651; // @[ISA_functions.scala 174:43:@7422.22]
    wire            _T_10669; // @[ISA_functions.scala 176:147:@7438.22]
    wire            _T_10670; // @[ISA_functions.scala 176:144:@7439.22]
    wire            _T_10671; // @[ISA_functions.scala 176:190:@7440.22]
    wire            _T_10672; // @[ISA_functions.scala 176:174:@7441.22]
    wire [31:0]     _T_10673; // @[ISA_functions.scala 176:217:@7442.22]
    wire [31:0]     _T_10674; // @[ISA_functions.scala 176:237:@7443.22]
    wire            _T_10675; // @[ISA_functions.scala 176:225:@7444.22]
    wire            _T_10676; // @[ISA_functions.scala 176:203:@7445.22]
    wire            _T_10703; // @[ISA_functions.scala 179:206:@7469.24]
    wire            _T_10704; // @[ISA_functions.scala 179:203:@7470.24]
    wire            _T_10727; // @[ISA_functions.scala 182:177:@7490.26]
    wire            _T_10728; // @[ISA_functions.scala 182:174:@7491.26]
    wire            _T_10729; // @[ISA_functions.scala 182:220:@7492.26]
    wire            _T_10730; // @[ISA_functions.scala 182:204:@7493.26]
    wire            _T_10731; // @[ISA_functions.scala 182:247:@7494.26]
    wire            _T_10732; // @[ISA_functions.scala 182:234:@7495.26]
    wire            _T_10761; // @[ISA_functions.scala 185:237:@7520.28]
    wire            _T_10762; // @[ISA_functions.scala 185:234:@7521.28]
    wire            _T_10789; // @[ISA_functions.scala 188:207:@7544.30]
    wire            _T_10790; // @[ISA_functions.scala 188:204:@7545.30]
    wire            _T_10791; // @[ISA_functions.scala 188:251:@7546.30]
    wire            _T_10792; // @[ISA_functions.scala 188:235:@7547.30]
    wire [18:0]     _T_10793; // @[ISA_functions.scala 189:55:@7549.32]
    wire [18:0]     _T_10795; // @[ISA_functions.scala 189:62:@7550.32]
    wire [524318:0] _GEN_6226; // @[ISA_functions.scala 189:43:@7551.32]
    wire [524318:0] _T_10796; // @[ISA_functions.scala 189:43:@7551.32]
    wire [31:0]     _T_10797; // @[ISA_functions.scala 189:76:@7552.32]
    wire            _T_10827; // @[ISA_functions.scala 191:238:@7577.32]
    wire            _T_10828; // @[ISA_functions.scala 191:235:@7578.32]
    wire            _T_10829; // @[ISA_functions.scala 191:281:@7579.32]
    wire            _T_10830; // @[ISA_functions.scala 191:265:@7580.32]
    wire [31:0]     _T_10833; // @[ISA_functions.scala 192:67:@7583.34]
    wire [31:0]     _T_10834; // @[ISA_functions.scala 192:53:@7584.34]
    wire [31:0]     _T_10835; // @[ISA_functions.scala 192:82:@7585.34]
    wire            _T_10869; // @[ISA_functions.scala 194:268:@7613.34]
    wire            _T_10870; // @[ISA_functions.scala 194:265:@7614.34]
    wire            _T_10871; // @[ISA_functions.scala 194:311:@7615.34]
    wire            _T_10872; // @[ISA_functions.scala 194:295:@7616.34]
    wire [31:0]     _T_10875; // @[ISA_functions.scala 195:43:@7619.36]
    wire            _T_10914; // @[ISA_functions.scala 197:298:@7651.36]
    wire            _T_10915; // @[ISA_functions.scala 197:295:@7652.36]
    wire            _T_10916; // @[ISA_functions.scala 197:341:@7653.36]
    wire            _T_10917; // @[ISA_functions.scala 197:325:@7654.36]
    wire [31:0]     _GEN_474; // @[ISA_functions.scala 197:357:@7655.36]
    wire [31:0]     _GEN_475; // @[ISA_functions.scala 194:325:@7617.34]
    wire [31:0]     _GEN_476; // @[ISA_functions.scala 191:295:@7581.32]
    wire [31:0]     _GEN_477; // @[ISA_functions.scala 188:265:@7548.30]
    wire [31:0]     _GEN_478; // @[ISA_functions.scala 185:261:@7522.28]
    wire [31:0]     _GEN_479; // @[ISA_functions.scala 182:260:@7496.26]
    wire [31:0]     _GEN_480; // @[ISA_functions.scala 179:248:@7471.24]
    wire [31:0]     _GEN_481; // @[ISA_functions.scala 176:247:@7446.22]
    wire [31:0]     _GEN_482; // @[ISA_functions.scala 173:174:@7421.20]
    wire [31:0]     _GEN_483; // @[ISA_functions.scala 170:144:@7403.18]
    wire [31:0]     _GEN_484; // @[ISA_functions.scala 167:115:@7388.16]
    wire [63:0]     _GEN_485; // @[ISA_functions.scala 164:85:@7374.14]
    wire [63:0]     _GEN_486; // @[ISA_functions.scala 161:50:@7364.12]
    wire [2:0]      _GEN_622; // @[ISA.scala 227:62:@1715.10]
    wire [31:0]     _GEN_623; // @[ISA.scala 227:62:@1715.10]
    wire [31:0]     _GEN_624; // @[ISA.scala 227:62:@1715.10]
    wire [31:0]     _GEN_625; // @[ISA.scala 227:62:@1715.10]
    wire [31:0]     _GEN_626; // @[ISA.scala 227:62:@1715.10]
    wire [31:0]     _GEN_627; // @[ISA.scala 227:62:@1715.10]
    wire [31:0]     _GEN_628; // @[ISA.scala 227:62:@1715.10]
    wire [63:0]     _GEN_629; // @[ISA.scala 227:62:@1715.10]
    wire [31:0]     _GEN_630; // @[ISA.scala 227:62:@1715.10]
    wire [31:0]     _GEN_631; // @[ISA.scala 227:62:@1715.10]
    wire [31:0]     _GEN_632; // @[ISA.scala 227:62:@1715.10]
    wire [31:0]     _GEN_633; // @[ISA.scala 227:62:@1715.10]
    wire [31:0]     _GEN_634; // @[ISA.scala 227:62:@1715.10]
    wire [63:0]     _GEN_635; // @[ISA.scala 227:62:@1715.10]
    wire            _GEN_636; // @[ISA.scala 227:62:@1715.10]
    wire            _GEN_637; // @[ISA.scala 227:62:@1715.10]
    wire            _GEN_638; // @[ISA.scala 227:62:@1715.10]
    wire [2:0]      _GEN_639; // @[ISA.scala 226:84:@1714.8]
    wire [31:0]     _GEN_640; // @[ISA.scala 226:84:@1714.8]
    wire [31:0]     _GEN_641; // @[ISA.scala 226:84:@1714.8]
    wire [31:0]     _GEN_642; // @[ISA.scala 226:84:@1714.8]
    wire [31:0]     _GEN_643; // @[ISA.scala 226:84:@1714.8]
    wire [31:0]     _GEN_644; // @[ISA.scala 226:84:@1714.8]
    wire [31:0]     _GEN_645; // @[ISA.scala 226:84:@1714.8]
    wire [63:0]     _GEN_646; // @[ISA.scala 226:84:@1714.8]
    wire [31:0]     _GEN_647; // @[ISA.scala 226:84:@1714.8]
    wire [31:0]     _GEN_648; // @[ISA.scala 226:84:@1714.8]
    wire [31:0]     _GEN_649; // @[ISA.scala 226:84:@1714.8]
    wire [31:0]     _GEN_650; // @[ISA.scala 226:84:@1714.8]
    wire [31:0]     _GEN_651; // @[ISA.scala 226:84:@1714.8]
    wire [63:0]     _GEN_652; // @[ISA.scala 226:84:@1714.8]
    wire            _GEN_653; // @[ISA.scala 226:84:@1714.8]
    wire            _GEN_654; // @[ISA.scala 226:84:@1714.8]
    wire            _GEN_655; // @[ISA.scala 226:84:@1714.8]
    wire [2:0]      _GEN_656; // @[ISA.scala 225:44:@1543.6]
    wire [31:0]     _GEN_657; // @[ISA.scala 225:44:@1543.6]
    wire [31:0]     _GEN_658; // @[ISA.scala 225:44:@1543.6]
    wire [31:0]     _GEN_659; // @[ISA.scala 225:44:@1543.6]
    wire [31:0]     _GEN_660; // @[ISA.scala 225:44:@1543.6]
    wire [31:0]     _GEN_661; // @[ISA.scala 225:44:@1543.6]
    wire [31:0]     _GEN_662; // @[ISA.scala 225:44:@1543.6]
    wire [63:0]     _GEN_663; // @[ISA.scala 225:44:@1543.6]
    wire [31:0]     _GEN_664; // @[ISA.scala 225:44:@1543.6]
    wire [31:0]     _GEN_665; // @[ISA.scala 225:44:@1543.6]
    wire [31:0]     _GEN_666; // @[ISA.scala 225:44:@1543.6]
    wire [31:0]     _GEN_667; // @[ISA.scala 225:44:@1543.6]
    wire [31:0]     _GEN_668; // @[ISA.scala 225:44:@1543.6]
    wire [63:0]     _GEN_669; // @[ISA.scala 225:44:@1543.6]
    wire            _GEN_670; // @[ISA.scala 225:44:@1543.6]
    wire            _GEN_671; // @[ISA.scala 225:44:@1543.6]
    wire            _GEN_672; // @[ISA.scala 225:44:@1543.6]
    wire            _T_31159; // @[ISA_functions.scala 91:81:@21596.14]
    wire            _T_31160; // @[ISA_functions.scala 91:67:@21597.14]
    wire            _T_31171; // @[ISA_functions.scala 251:71:@21604.16]
    wire            _T_31176; // @[ISA_functions.scala 251:120:@21607.16]
    wire [31:0]     _T_31178; // @[ISA_functions.scala 251:190:@21608.16]
    wire [31:0]     _T_31181; // @[ISA_functions.scala 251:212:@21610.16]
    wire            _T_31183; // @[ISA_functions.scala 251:225:@21611.16]
    wire            _T_31184; // @[ISA_functions.scala 251:171:@21612.16]
    wire            _T_31210; // @[ISA_functions.scala 254:179:@21631.18]
    wire            _T_31211; // @[ISA_functions.scala 254:176:@21632.18]
    wire [31:0]     _T_31217; // @[ISA_functions.scala 255:57:@21637.20]
    wire            _T_31233; // @[ISA_functions.scala 257:28:@21649.20]
    wire            _T_31238; // @[ISA_functions.scala 257:177:@21652.20]
    wire            _T_31246; // @[ISA_functions.scala 257:226:@21657.20]
    wire [31:0]     _T_31251; // @[ISA_functions.scala 258:71:@21661.22]
    wire [31:0]     _T_31257; // @[ISA_functions.scala 258:87:@21665.22]
    wire            _T_31288; // @[ISA_functions.scala 260:226:@21686.22]
    wire [31:0]     _T_31302; // @[ISA_functions.scala 261:57:@21696.24]
    wire            _T_31325; // @[ISA_functions.scala 263:177:@21712.24]
    wire            _T_31330; // @[ISA_functions.scala 263:227:@21715.24]
    wire            _T_31338; // @[ISA_functions.scala 263:276:@21720.24]
    wire [524318:0] _GEN_6231; // @[ISA_functions.scala 264:50:@21722.26]
    wire [524318:0] _T_31340; // @[ISA_functions.scala 264:50:@21722.26]
    wire [31:0]     _T_31341; // @[ISA_functions.scala 264:63:@21723.26]
    wire [31:0]     _T_31343; // @[ISA_functions.scala 264:71:@21724.26]
    wire [31:0]     _T_31348; // @[ISA_functions.scala 264:126:@21727.26]
    wire [31:0]     _T_31349; // @[ISA_functions.scala 264:87:@21728.26]
    wire [31:0]     _T_31354; // @[ISA_functions.scala 264:181:@21731.26]
    wire [31:0]     _T_31355; // @[ISA_functions.scala 264:143:@21732.26]
    wire            _T_31393; // @[ISA_functions.scala 266:276:@21757.26]
    wire [31:0]     _T_31413; // @[ISA_functions.scala 267:57:@21771.28]
    wire            _T_31443; // @[ISA_functions.scala 269:227:@21791.28]
    wire            _T_31453; // @[ISA_functions.scala 269:277:@21797.28]
    wire [31:0]     _T_31456; // @[ISA_functions.scala 270:47:@21800.30]
    wire            _T_31498; // @[ISA_functions.scala 272:277:@21827.30]
    wire            _T_31503; // @[ISA_functions.scala 272:378:@21830.30]
    wire            _T_31511; // @[ISA_functions.scala 272:428:@21835.30]
    wire [31:0]     _T_31513; // @[ISA_functions.scala 273:49:@21837.32]
    wire [31:0]     _T_31515; // @[ISA_functions.scala 273:85:@21838.32]
    wire [31:0]     _T_31518; // @[ISA_functions.scala 273:106:@21840.32]
    wire [31:0]     _T_31519; // @[ISA_functions.scala 273:68:@21841.32]
    wire [31:0]     _T_31524; // @[ISA_functions.scala 273:162:@21844.32]
    wire [31:0]     _T_31525; // @[ISA_functions.scala 273:123:@21845.32]
    wire            _T_31582; // @[ISA_functions.scala 275:428:@21881.32]
    wire [31:0]     _T_31599; // @[ISA_functions.scala 276:60:@21893.34]
    wire [31:0]     _GEN_868; // @[ISA_functions.scala 275:499:@21882.32]
    wire [31:0]     _GEN_869; // @[ISA_functions.scala 272:498:@21836.30]
    wire [31:0]     _GEN_870; // @[ISA_functions.scala 269:378:@21798.28]
    wire [31:0]     _GEN_871; // @[ISA_functions.scala 266:347:@21758.26]
    wire [31:0]     _GEN_872; // @[ISA_functions.scala 263:346:@21721.24]
    wire [31:0]     _GEN_873; // @[ISA_functions.scala 260:297:@21687.22]
    wire [31:0]     _GEN_874; // @[ISA_functions.scala 257:296:@21658.20]
    wire [31:0]     _GEN_875; // @[ISA_functions.scala 254:247:@21633.18]
    wire [31:0]     _GEN_876; // @[ISA_functions.scala 251:241:@21613.16]
    wire [32:0]     _T_31601; // @[ISA_functions.scala 92:40:@21899.16]
    wire [31:0]     _T_31602; // @[ISA_functions.scala 92:40:@21900.16]
    wire            _T_34242; // @[ISA_functions.scala 94:28:@23640.16]
    wire            _T_36879; // @[ISA_functions.scala 94:164:@25375.16]
    wire            _T_36880; // @[ISA_functions.scala 94:150:@25376.16]
    wire            _T_36881; // @[ISA_functions.scala 94:103:@25377.16]
    wire            _T_42603; // @[ISA_functions.scala 97:106:@29157.18]
    wire            _T_42604; // @[ISA_functions.scala 97:103:@29158.18]
    wire            _T_45241; // @[ISA_functions.scala 97:242:@30893.18]
    wire            _T_45242; // @[ISA_functions.scala 97:228:@30894.18]
    wire            _T_45243; // @[ISA_functions.scala 97:181:@30895.18]
    wire            _T_53606; // @[ISA_functions.scala 100:184:@36413.20]
    wire            _T_53607; // @[ISA_functions.scala 100:181:@36414.20]
    wire            _T_56245; // @[ISA_functions.scala 100:306:@38150.20]
    wire            _T_56246; // @[ISA_functions.scala 100:259:@38151.20]
    wire            _T_67250; // @[ISA_functions.scala 103:262:@45407.22]
    wire            _T_67251; // @[ISA_functions.scala 103:259:@45408.22]
    wire            _T_69889; // @[ISA_functions.scala 103:385:@47144.22]
    wire            _T_69890; // @[ISA_functions.scala 103:337:@47145.22]
    wire            _T_83535; // @[ISA_functions.scala 106:340:@56139.24]
    wire            _T_83536; // @[ISA_functions.scala 106:337:@56140.24]
    wire            _T_86174; // @[ISA_functions.scala 106:464:@57876.24]
    wire            _T_86175; // @[ISA_functions.scala 106:416:@57877.24]
    wire [32:0]     _T_86619; // @[ISA_functions.scala 110:40:@58184.26]
    wire [31:0]     _T_86620; // @[ISA_functions.scala 110:40:@58185.26]
    wire [31:0]     _GEN_1822; // @[ISA_functions.scala 106:495:@57878.24]
    wire [31:0]     _GEN_1823; // @[ISA_functions.scala 103:416:@47146.22]
    wire [31:0]     _GEN_1824; // @[ISA_functions.scala 100:337:@38152.20]
    wire [31:0]     _GEN_1825; // @[ISA_functions.scala 97:259:@30896.18]
    wire [31:0]     _GEN_1826; // @[ISA_functions.scala 94:181:@25378.16]
    wire [31:0]     _GEN_1827; // @[ISA_functions.scala 91:98:@21598.14]
    wire [2:0]      _GEN_4106; // @[ISA.scala 251:70:@13955.12]
    wire [31:0]     _GEN_4107; // @[ISA.scala 251:70:@13955.12]
    wire [31:0]     _GEN_4108; // @[ISA.scala 251:70:@13955.12]
    wire [31:0]     _GEN_4109; // @[ISA.scala 251:70:@13955.12]
    wire [31:0]     _GEN_4110; // @[ISA.scala 251:70:@13955.12]
    wire [31:0]     _GEN_4111; // @[ISA.scala 251:70:@13955.12]
    wire [31:0]     _GEN_4112; // @[ISA.scala 251:70:@13955.12]
    wire [63:0]     _GEN_4113; // @[ISA.scala 251:70:@13955.12]
    wire [31:0]     _GEN_4114; // @[ISA.scala 251:70:@13955.12]
    wire [31:0]     _GEN_4115; // @[ISA.scala 251:70:@13955.12]
    wire [31:0]     _GEN_4116; // @[ISA.scala 251:70:@13955.12]
    wire [31:0]     _GEN_4117; // @[ISA.scala 251:70:@13955.12]
    wire            _GEN_4118; // @[ISA.scala 251:70:@13955.12]
    wire            _GEN_4119; // @[ISA.scala 251:70:@13955.12]
    wire            _GEN_4120; // @[ISA.scala 251:70:@13955.12]
    wire [2:0]      _GEN_4121; // @[ISA.scala 250:92:@13954.10]
    wire [31:0]     _GEN_4122; // @[ISA.scala 250:92:@13954.10]
    wire [31:0]     _GEN_4123; // @[ISA.scala 250:92:@13954.10]
    wire [31:0]     _GEN_4124; // @[ISA.scala 250:92:@13954.10]
    wire [31:0]     _GEN_4125; // @[ISA.scala 250:92:@13954.10]
    wire [31:0]     _GEN_4126; // @[ISA.scala 250:92:@13954.10]
    wire [31:0]     _GEN_4127; // @[ISA.scala 250:92:@13954.10]
    wire [63:0]     _GEN_4128; // @[ISA.scala 250:92:@13954.10]
    wire [31:0]     _GEN_4129; // @[ISA.scala 250:92:@13954.10]
    wire [31:0]     _GEN_4130; // @[ISA.scala 250:92:@13954.10]
    wire [31:0]     _GEN_4131; // @[ISA.scala 250:92:@13954.10]
    wire [31:0]     _GEN_4132; // @[ISA.scala 250:92:@13954.10]
    wire            _GEN_4133; // @[ISA.scala 250:92:@13954.10]
    wire            _GEN_4134; // @[ISA.scala 250:92:@13954.10]
    wire            _GEN_4135; // @[ISA.scala 250:92:@13954.10]
    wire [2:0]      _GEN_4136; // @[ISA.scala 249:85:@13783.8]
    wire [31:0]     _GEN_4137; // @[ISA.scala 249:85:@13783.8]
    wire [31:0]     _GEN_4138; // @[ISA.scala 249:85:@13783.8]
    wire [31:0]     _GEN_4139; // @[ISA.scala 249:85:@13783.8]
    wire [31:0]     _GEN_4140; // @[ISA.scala 249:85:@13783.8]
    wire [31:0]     _GEN_4141; // @[ISA.scala 249:85:@13783.8]
    wire [31:0]     _GEN_4142; // @[ISA.scala 249:85:@13783.8]
    wire [63:0]     _GEN_4143; // @[ISA.scala 249:85:@13783.8]
    wire [31:0]     _GEN_4144; // @[ISA.scala 249:85:@13783.8]
    wire [31:0]     _GEN_4145; // @[ISA.scala 249:85:@13783.8]
    wire [31:0]     _GEN_4146; // @[ISA.scala 249:85:@13783.8]
    wire [31:0]     _GEN_4147; // @[ISA.scala 249:85:@13783.8]
    wire            _GEN_4148; // @[ISA.scala 249:85:@13783.8]
    wire            _GEN_4149; // @[ISA.scala 249:85:@13783.8]
    wire            _GEN_4150; // @[ISA.scala 249:85:@13783.8]
    wire [2:0]      _GEN_4151; // @[ISA.scala 248:44:@13611.6]
    wire [31:0]     _GEN_4152; // @[ISA.scala 248:44:@13611.6]
    wire [31:0]     _GEN_4153; // @[ISA.scala 248:44:@13611.6]
    wire [31:0]     _GEN_4154; // @[ISA.scala 248:44:@13611.6]
    wire [31:0]     _GEN_4155; // @[ISA.scala 248:44:@13611.6]
    wire [31:0]     _GEN_4156; // @[ISA.scala 248:44:@13611.6]
    wire [31:0]     _GEN_4157; // @[ISA.scala 248:44:@13611.6]
    wire [63:0]     _GEN_4158; // @[ISA.scala 248:44:@13611.6]
    wire [31:0]     _GEN_4159; // @[ISA.scala 248:44:@13611.6]
    wire [31:0]     _GEN_4160; // @[ISA.scala 248:44:@13611.6]
    wire [31:0]     _GEN_4161; // @[ISA.scala 248:44:@13611.6]
    wire [31:0]     _GEN_4162; // @[ISA.scala 248:44:@13611.6]
    wire            _GEN_4163; // @[ISA.scala 248:44:@13611.6]
    wire            _GEN_4164; // @[ISA.scala 248:44:@13611.6]
    wire            _GEN_4165; // @[ISA.scala 248:44:@13611.6]
    wire [32:0]     _T_223492; // @[ISA_functions.scala 162:43:@149070.18]
    wire [31:0]     _T_223493; // @[ISA_functions.scala 162:43:@149071.18]
    wire [63:0]     _T_223500; // @[ISA_functions.scala 165:55:@149080.20]
    wire [64:0]     _T_223501; // @[ISA_functions.scala 165:43:@149081.20]
    wire [63:0]     _T_223502; // @[ISA_functions.scala 165:43:@149082.20]
    wire [31:0]     _T_223512; // @[ISA_functions.scala 168:43:@149094.22]
    wire [31:0]     _T_223526; // @[ISA_functions.scala 171:43:@149109.24]
    wire [31:0]     _T_223544; // @[ISA_functions.scala 174:43:@149127.26]
    wire [31:0]     _T_223567; // @[ISA_functions.scala 176:237:@149148.26]
    wire            _T_223568; // @[ISA_functions.scala 176:225:@149149.26]
    wire            _T_223596; // @[ISA_functions.scala 179:206:@149174.28]
    wire            _T_223624; // @[ISA_functions.scala 182:247:@149199.30]
    wire            _T_223654; // @[ISA_functions.scala 185:237:@149225.32]
    wire [18:0]     _T_223686; // @[ISA_functions.scala 189:55:@149254.36]
    wire [18:0]     _T_223688; // @[ISA_functions.scala 189:62:@149255.36]
    wire [524318:0] _T_223689; // @[ISA_functions.scala 189:43:@149256.36]
    wire [31:0]     _T_223690; // @[ISA_functions.scala 189:76:@149257.36]
    wire [31:0]     _T_223726; // @[ISA_functions.scala 192:67:@149288.38]
    wire [31:0]     _T_223727; // @[ISA_functions.scala 192:53:@149289.38]
    wire [31:0]     _T_223728; // @[ISA_functions.scala 192:82:@149290.38]
    wire [31:0]     _T_223768; // @[ISA_functions.scala 195:43:@149324.40]
    wire [63:0]     _GEN_4243; // @[ISA_functions.scala 161:50:@149069.16]
    wire            _T_228862; // @[ISA_functions.scala 429:45:@152675.16]
    wire            _T_228873; // @[ISA_functions.scala 432:28:@152683.18]
    wire            _T_228876; // @[ISA_functions.scala 432:101:@152686.18]
    wire            _T_228877; // @[ISA_functions.scala 432:76:@152687.18]
    wire            _T_228887; // @[ISA_functions.scala 435:79:@152699.20]
    wire            _T_228888; // @[ISA_functions.scala 435:76:@152700.20]
    wire            _T_228891; // @[ISA_functions.scala 435:152:@152703.20]
    wire            _T_228892; // @[ISA_functions.scala 435:127:@152704.20]
    wire            _T_228908; // @[ISA_functions.scala 438:130:@152721.22]
    wire            _T_228909; // @[ISA_functions.scala 438:127:@152722.22]
    wire            _T_228911; // @[ISA_functions.scala 438:178:@152724.22]
    wire            _T_228931; // @[ISA_functions.scala 441:181:@152744.24]
    wire            _T_228932; // @[ISA_functions.scala 441:178:@152745.24]
    wire            _T_228934; // @[ISA_functions.scala 441:204:@152747.24]
    wire [31:0]     _GEN_4321; // @[ISA_functions.scala 441:230:@152748.24]
    wire [31:0]     _GEN_4322; // @[ISA_functions.scala 438:204:@152725.22]
    wire [31:0]     _GEN_4323; // @[ISA_functions.scala 435:178:@152705.20]
    wire [31:0]     _GEN_4324; // @[ISA_functions.scala 432:127:@152688.18]
    wire [31:0]     _GEN_4325; // @[ISA_functions.scala 429:71:@152676.16]
    wire [2:0]      _GEN_4462; // @[ISA.scala 275:78:@147185.14]
    wire [63:0]     _GEN_4463; // @[ISA.scala 275:78:@147185.14]
    wire [31:0]     _GEN_4464; // @[ISA.scala 275:78:@147185.14]
    wire [31:0]     _GEN_4465; // @[ISA.scala 275:78:@147185.14]
    wire [31:0]     _GEN_4466; // @[ISA.scala 275:78:@147185.14]
    wire [31:0]     _GEN_4467; // @[ISA.scala 275:78:@147185.14]
    wire [31:0]     _GEN_4468; // @[ISA.scala 275:78:@147185.14]
    wire [63:0]     _GEN_4469; // @[ISA.scala 275:78:@147185.14]
    wire [63:0]     _GEN_4470; // @[ISA.scala 275:78:@147185.14]
    wire [31:0]     _GEN_4471; // @[ISA.scala 275:78:@147185.14]
    wire [31:0]     _GEN_4472; // @[ISA.scala 275:78:@147185.14]
    wire [31:0]     _GEN_4473; // @[ISA.scala 275:78:@147185.14]
    wire            _GEN_4474; // @[ISA.scala 275:78:@147185.14]
    wire            _GEN_4475; // @[ISA.scala 275:78:@147185.14]
    wire            _GEN_4476; // @[ISA.scala 275:78:@147185.14]
    wire [2:0]      _GEN_4477; // @[ISA.scala 274:100:@147184.12]
    wire [63:0]     _GEN_4478; // @[ISA.scala 274:100:@147184.12]
    wire [31:0]     _GEN_4479; // @[ISA.scala 274:100:@147184.12]
    wire [31:0]     _GEN_4480; // @[ISA.scala 274:100:@147184.12]
    wire [31:0]     _GEN_4481; // @[ISA.scala 274:100:@147184.12]
    wire [31:0]     _GEN_4482; // @[ISA.scala 274:100:@147184.12]
    wire [31:0]     _GEN_4483; // @[ISA.scala 274:100:@147184.12]
    wire [63:0]     _GEN_4484; // @[ISA.scala 274:100:@147184.12]
    wire [63:0]     _GEN_4485; // @[ISA.scala 274:100:@147184.12]
    wire [31:0]     _GEN_4486; // @[ISA.scala 274:100:@147184.12]
    wire [31:0]     _GEN_4487; // @[ISA.scala 274:100:@147184.12]
    wire [31:0]     _GEN_4488; // @[ISA.scala 274:100:@147184.12]
    wire            _GEN_4489; // @[ISA.scala 274:100:@147184.12]
    wire            _GEN_4490; // @[ISA.scala 274:100:@147184.12]
    wire            _GEN_4491; // @[ISA.scala 274:100:@147184.12]
    wire [2:0]      _GEN_4492; // @[ISA.scala 273:93:@147013.10]
    wire [63:0]     _GEN_4493; // @[ISA.scala 273:93:@147013.10]
    wire [31:0]     _GEN_4494; // @[ISA.scala 273:93:@147013.10]
    wire [31:0]     _GEN_4495; // @[ISA.scala 273:93:@147013.10]
    wire [31:0]     _GEN_4496; // @[ISA.scala 273:93:@147013.10]
    wire [31:0]     _GEN_4497; // @[ISA.scala 273:93:@147013.10]
    wire [31:0]     _GEN_4498; // @[ISA.scala 273:93:@147013.10]
    wire [63:0]     _GEN_4499; // @[ISA.scala 273:93:@147013.10]
    wire [63:0]     _GEN_4500; // @[ISA.scala 273:93:@147013.10]
    wire [31:0]     _GEN_4501; // @[ISA.scala 273:93:@147013.10]
    wire [31:0]     _GEN_4502; // @[ISA.scala 273:93:@147013.10]
    wire [31:0]     _GEN_4503; // @[ISA.scala 273:93:@147013.10]
    wire            _GEN_4504; // @[ISA.scala 273:93:@147013.10]
    wire            _GEN_4505; // @[ISA.scala 273:93:@147013.10]
    wire            _GEN_4506; // @[ISA.scala 273:93:@147013.10]
    wire [2:0]      _GEN_4507; // @[ISA.scala 272:85:@146841.8]
    wire [63:0]     _GEN_4508; // @[ISA.scala 272:85:@146841.8]
    wire [31:0]     _GEN_4509; // @[ISA.scala 272:85:@146841.8]
    wire [31:0]     _GEN_4510; // @[ISA.scala 272:85:@146841.8]
    wire [31:0]     _GEN_4511; // @[ISA.scala 272:85:@146841.8]
    wire [31:0]     _GEN_4512; // @[ISA.scala 272:85:@146841.8]
    wire [31:0]     _GEN_4513; // @[ISA.scala 272:85:@146841.8]
    wire [63:0]     _GEN_4514; // @[ISA.scala 272:85:@146841.8]
    wire [63:0]     _GEN_4515; // @[ISA.scala 272:85:@146841.8]
    wire [31:0]     _GEN_4516; // @[ISA.scala 272:85:@146841.8]
    wire [31:0]     _GEN_4517; // @[ISA.scala 272:85:@146841.8]
    wire [31:0]     _GEN_4518; // @[ISA.scala 272:85:@146841.8]
    wire            _GEN_4519; // @[ISA.scala 272:85:@146841.8]
    wire            _GEN_4520; // @[ISA.scala 272:85:@146841.8]
    wire            _GEN_4521; // @[ISA.scala 272:85:@146841.8]
    wire [2:0]      _GEN_4522; // @[ISA.scala 271:44:@146669.6]
    wire [63:0]     _GEN_4523; // @[ISA.scala 271:44:@146669.6]
    wire [31:0]     _GEN_4524; // @[ISA.scala 271:44:@146669.6]
    wire [31:0]     _GEN_4525; // @[ISA.scala 271:44:@146669.6]
    wire [31:0]     _GEN_4526; // @[ISA.scala 271:44:@146669.6]
    wire [31:0]     _GEN_4527; // @[ISA.scala 271:44:@146669.6]
    wire [31:0]     _GEN_4528; // @[ISA.scala 271:44:@146669.6]
    wire [63:0]     _GEN_4529; // @[ISA.scala 271:44:@146669.6]
    wire [63:0]     _GEN_4530; // @[ISA.scala 271:44:@146669.6]
    wire [31:0]     _GEN_4531; // @[ISA.scala 271:44:@146669.6]
    wire [31:0]     _GEN_4532; // @[ISA.scala 271:44:@146669.6]
    wire [31:0]     _GEN_4533; // @[ISA.scala 271:44:@146669.6]
    wire            _GEN_4534; // @[ISA.scala 271:44:@146669.6]
    wire            _GEN_4535; // @[ISA.scala 271:44:@146669.6]
    wire            _GEN_4536; // @[ISA.scala 271:44:@146669.6]
    wire [63:0]     _GEN_6281; // @[ISA_functions.scala 165:43:@161117.24]
    wire [63:0]     _GEN_4658; // @[ISA_functions.scala 161:50:@161706.20]
    wire [63:0]     _GEN_4659; // @[ISA_functions.scala 240:67:@160802.18]
    wire [2:0]      _GEN_4751; // @[ISA.scala 301:86:@159025.16]
    wire [63:0]     _GEN_4752; // @[ISA.scala 301:86:@159025.16]
    wire [31:0]     _GEN_4753; // @[ISA.scala 301:86:@159025.16]
    wire [31:0]     _GEN_4754; // @[ISA.scala 301:86:@159025.16]
    wire [31:0]     _GEN_4755; // @[ISA.scala 301:86:@159025.16]
    wire [31:0]     _GEN_4756; // @[ISA.scala 301:86:@159025.16]
    wire [31:0]     _GEN_4757; // @[ISA.scala 301:86:@159025.16]
    wire [63:0]     _GEN_4758; // @[ISA.scala 301:86:@159025.16]
    wire [63:0]     _GEN_4759; // @[ISA.scala 301:86:@159025.16]
    wire [31:0]     _GEN_4760; // @[ISA.scala 301:86:@159025.16]
    wire [31:0]     _GEN_4761; // @[ISA.scala 301:86:@159025.16]
    wire [31:0]     _GEN_4762; // @[ISA.scala 301:86:@159025.16]
    wire [31:0]     _GEN_4763; // @[ISA.scala 301:86:@159025.16]
    wire [63:0]     _GEN_4764; // @[ISA.scala 301:86:@159025.16]
    wire            _GEN_4765; // @[ISA.scala 301:86:@159025.16]
    wire            _GEN_4766; // @[ISA.scala 301:86:@159025.16]
    wire            _GEN_4767; // @[ISA.scala 301:86:@159025.16]
    wire [2:0]      _GEN_4768; // @[ISA.scala 300:108:@159024.14]
    wire [63:0]     _GEN_4769; // @[ISA.scala 300:108:@159024.14]
    wire [31:0]     _GEN_4770; // @[ISA.scala 300:108:@159024.14]
    wire [31:0]     _GEN_4771; // @[ISA.scala 300:108:@159024.14]
    wire [31:0]     _GEN_4772; // @[ISA.scala 300:108:@159024.14]
    wire [31:0]     _GEN_4773; // @[ISA.scala 300:108:@159024.14]
    wire [31:0]     _GEN_4774; // @[ISA.scala 300:108:@159024.14]
    wire [63:0]     _GEN_4775; // @[ISA.scala 300:108:@159024.14]
    wire [63:0]     _GEN_4776; // @[ISA.scala 300:108:@159024.14]
    wire [31:0]     _GEN_4777; // @[ISA.scala 300:108:@159024.14]
    wire [31:0]     _GEN_4778; // @[ISA.scala 300:108:@159024.14]
    wire [31:0]     _GEN_4779; // @[ISA.scala 300:108:@159024.14]
    wire [31:0]     _GEN_4780; // @[ISA.scala 300:108:@159024.14]
    wire [63:0]     _GEN_4781; // @[ISA.scala 300:108:@159024.14]
    wire            _GEN_4782; // @[ISA.scala 300:108:@159024.14]
    wire            _GEN_4783; // @[ISA.scala 300:108:@159024.14]
    wire            _GEN_4784; // @[ISA.scala 300:108:@159024.14]
    wire [2:0]      _GEN_4785; // @[ISA.scala 299:101:@158853.12]
    wire [63:0]     _GEN_4786; // @[ISA.scala 299:101:@158853.12]
    wire [31:0]     _GEN_4787; // @[ISA.scala 299:101:@158853.12]
    wire [31:0]     _GEN_4788; // @[ISA.scala 299:101:@158853.12]
    wire [31:0]     _GEN_4789; // @[ISA.scala 299:101:@158853.12]
    wire [31:0]     _GEN_4790; // @[ISA.scala 299:101:@158853.12]
    wire [31:0]     _GEN_4791; // @[ISA.scala 299:101:@158853.12]
    wire [63:0]     _GEN_4792; // @[ISA.scala 299:101:@158853.12]
    wire [63:0]     _GEN_4793; // @[ISA.scala 299:101:@158853.12]
    wire [31:0]     _GEN_4794; // @[ISA.scala 299:101:@158853.12]
    wire [31:0]     _GEN_4795; // @[ISA.scala 299:101:@158853.12]
    wire [31:0]     _GEN_4796; // @[ISA.scala 299:101:@158853.12]
    wire [31:0]     _GEN_4797; // @[ISA.scala 299:101:@158853.12]
    wire [63:0]     _GEN_4798; // @[ISA.scala 299:101:@158853.12]
    wire            _GEN_4799; // @[ISA.scala 299:101:@158853.12]
    wire            _GEN_4800; // @[ISA.scala 299:101:@158853.12]
    wire            _GEN_4801; // @[ISA.scala 299:101:@158853.12]
    wire [2:0]      _GEN_4802; // @[ISA.scala 298:93:@158681.10]
    wire [63:0]     _GEN_4803; // @[ISA.scala 298:93:@158681.10]
    wire [31:0]     _GEN_4804; // @[ISA.scala 298:93:@158681.10]
    wire [31:0]     _GEN_4805; // @[ISA.scala 298:93:@158681.10]
    wire [31:0]     _GEN_4806; // @[ISA.scala 298:93:@158681.10]
    wire [31:0]     _GEN_4807; // @[ISA.scala 298:93:@158681.10]
    wire [31:0]     _GEN_4808; // @[ISA.scala 298:93:@158681.10]
    wire [63:0]     _GEN_4809; // @[ISA.scala 298:93:@158681.10]
    wire [63:0]     _GEN_4810; // @[ISA.scala 298:93:@158681.10]
    wire [31:0]     _GEN_4811; // @[ISA.scala 298:93:@158681.10]
    wire [31:0]     _GEN_4812; // @[ISA.scala 298:93:@158681.10]
    wire [31:0]     _GEN_4813; // @[ISA.scala 298:93:@158681.10]
    wire [31:0]     _GEN_4814; // @[ISA.scala 298:93:@158681.10]
    wire [63:0]     _GEN_4815; // @[ISA.scala 298:93:@158681.10]
    wire            _GEN_4816; // @[ISA.scala 298:93:@158681.10]
    wire            _GEN_4817; // @[ISA.scala 298:93:@158681.10]
    wire            _GEN_4818; // @[ISA.scala 298:93:@158681.10]
    wire [2:0]      _GEN_4819; // @[ISA.scala 297:85:@158509.8]
    wire [63:0]     _GEN_4820; // @[ISA.scala 297:85:@158509.8]
    wire [31:0]     _GEN_4821; // @[ISA.scala 297:85:@158509.8]
    wire [31:0]     _GEN_4822; // @[ISA.scala 297:85:@158509.8]
    wire [31:0]     _GEN_4823; // @[ISA.scala 297:85:@158509.8]
    wire [31:0]     _GEN_4824; // @[ISA.scala 297:85:@158509.8]
    wire [31:0]     _GEN_4825; // @[ISA.scala 297:85:@158509.8]
    wire [63:0]     _GEN_4826; // @[ISA.scala 297:85:@158509.8]
    wire [63:0]     _GEN_4827; // @[ISA.scala 297:85:@158509.8]
    wire [31:0]     _GEN_4828; // @[ISA.scala 297:85:@158509.8]
    wire [31:0]     _GEN_4829; // @[ISA.scala 297:85:@158509.8]
    wire [31:0]     _GEN_4830; // @[ISA.scala 297:85:@158509.8]
    wire [31:0]     _GEN_4831; // @[ISA.scala 297:85:@158509.8]
    wire [63:0]     _GEN_4832; // @[ISA.scala 297:85:@158509.8]
    wire            _GEN_4833; // @[ISA.scala 297:85:@158509.8]
    wire            _GEN_4834; // @[ISA.scala 297:85:@158509.8]
    wire            _GEN_4835; // @[ISA.scala 297:85:@158509.8]
    wire [2:0]      _GEN_4836; // @[ISA.scala 296:44:@158337.6]
    wire [63:0]     _GEN_4837; // @[ISA.scala 296:44:@158337.6]
    wire [31:0]     _GEN_4838; // @[ISA.scala 296:44:@158337.6]
    wire [31:0]     _GEN_4839; // @[ISA.scala 296:44:@158337.6]
    wire [31:0]     _GEN_4840; // @[ISA.scala 296:44:@158337.6]
    wire [31:0]     _GEN_4841; // @[ISA.scala 296:44:@158337.6]
    wire [31:0]     _GEN_4842; // @[ISA.scala 296:44:@158337.6]
    wire [63:0]     _GEN_4843; // @[ISA.scala 296:44:@158337.6]
    wire [63:0]     _GEN_4844; // @[ISA.scala 296:44:@158337.6]
    wire [31:0]     _GEN_4845; // @[ISA.scala 296:44:@158337.6]
    wire [31:0]     _GEN_4846; // @[ISA.scala 296:44:@158337.6]
    wire [31:0]     _GEN_4847; // @[ISA.scala 296:44:@158337.6]
    wire [31:0]     _GEN_4848; // @[ISA.scala 296:44:@158337.6]
    wire [63:0]     _GEN_4849; // @[ISA.scala 296:44:@158337.6]
    wire            _GEN_4850; // @[ISA.scala 296:44:@158337.6]
    wire            _GEN_4851; // @[ISA.scala 296:44:@158337.6]
    wire            _GEN_4852; // @[ISA.scala 296:44:@158337.6]
    wire [2:0]      _GEN_4922; // @[ISA.scala 331:94:@165852.18]
    wire [63:0]     _GEN_4923; // @[ISA.scala 331:94:@165852.18]
    wire [31:0]     _GEN_4924; // @[ISA.scala 331:94:@165852.18]
    wire [31:0]     _GEN_4925; // @[ISA.scala 331:94:@165852.18]
    wire [31:0]     _GEN_4926; // @[ISA.scala 331:94:@165852.18]
    wire [31:0]     _GEN_4927; // @[ISA.scala 331:94:@165852.18]
    wire [31:0]     _GEN_4928; // @[ISA.scala 331:94:@165852.18]
    wire [63:0]     _GEN_4929; // @[ISA.scala 331:94:@165852.18]
    wire [63:0]     _GEN_4930; // @[ISA.scala 331:94:@165852.18]
    wire [31:0]     _GEN_4931; // @[ISA.scala 331:94:@165852.18]
    wire [31:0]     _GEN_4932; // @[ISA.scala 331:94:@165852.18]
    wire [31:0]     _GEN_4933; // @[ISA.scala 331:94:@165852.18]
    wire [31:0]     _GEN_4934; // @[ISA.scala 331:94:@165852.18]
    wire [63:0]     _GEN_4935; // @[ISA.scala 331:94:@165852.18]
    wire            _GEN_4936; // @[ISA.scala 331:94:@165852.18]
    wire            _GEN_4937; // @[ISA.scala 331:94:@165852.18]
    wire            _GEN_4938; // @[ISA.scala 331:94:@165852.18]
    wire [2:0]      _GEN_4939; // @[ISA.scala 330:116:@165851.16]
    wire [63:0]     _GEN_4940; // @[ISA.scala 330:116:@165851.16]
    wire [31:0]     _GEN_4941; // @[ISA.scala 330:116:@165851.16]
    wire [31:0]     _GEN_4942; // @[ISA.scala 330:116:@165851.16]
    wire [31:0]     _GEN_4943; // @[ISA.scala 330:116:@165851.16]
    wire [31:0]     _GEN_4944; // @[ISA.scala 330:116:@165851.16]
    wire [31:0]     _GEN_4945; // @[ISA.scala 330:116:@165851.16]
    wire [63:0]     _GEN_4946; // @[ISA.scala 330:116:@165851.16]
    wire [63:0]     _GEN_4947; // @[ISA.scala 330:116:@165851.16]
    wire [31:0]     _GEN_4948; // @[ISA.scala 330:116:@165851.16]
    wire [31:0]     _GEN_4949; // @[ISA.scala 330:116:@165851.16]
    wire [31:0]     _GEN_4950; // @[ISA.scala 330:116:@165851.16]
    wire [31:0]     _GEN_4951; // @[ISA.scala 330:116:@165851.16]
    wire [63:0]     _GEN_4952; // @[ISA.scala 330:116:@165851.16]
    wire            _GEN_4953; // @[ISA.scala 330:116:@165851.16]
    wire            _GEN_4954; // @[ISA.scala 330:116:@165851.16]
    wire            _GEN_4955; // @[ISA.scala 330:116:@165851.16]
    wire [2:0]      _GEN_4956; // @[ISA.scala 329:109:@165680.14]
    wire [63:0]     _GEN_4957; // @[ISA.scala 329:109:@165680.14]
    wire [31:0]     _GEN_4958; // @[ISA.scala 329:109:@165680.14]
    wire [31:0]     _GEN_4959; // @[ISA.scala 329:109:@165680.14]
    wire [31:0]     _GEN_4960; // @[ISA.scala 329:109:@165680.14]
    wire [31:0]     _GEN_4961; // @[ISA.scala 329:109:@165680.14]
    wire [31:0]     _GEN_4962; // @[ISA.scala 329:109:@165680.14]
    wire [63:0]     _GEN_4963; // @[ISA.scala 329:109:@165680.14]
    wire [63:0]     _GEN_4964; // @[ISA.scala 329:109:@165680.14]
    wire [31:0]     _GEN_4965; // @[ISA.scala 329:109:@165680.14]
    wire [31:0]     _GEN_4966; // @[ISA.scala 329:109:@165680.14]
    wire [31:0]     _GEN_4967; // @[ISA.scala 329:109:@165680.14]
    wire [31:0]     _GEN_4968; // @[ISA.scala 329:109:@165680.14]
    wire [63:0]     _GEN_4969; // @[ISA.scala 329:109:@165680.14]
    wire            _GEN_4970; // @[ISA.scala 329:109:@165680.14]
    wire            _GEN_4971; // @[ISA.scala 329:109:@165680.14]
    wire            _GEN_4972; // @[ISA.scala 329:109:@165680.14]
    wire [2:0]      _GEN_4973; // @[ISA.scala 328:101:@165508.12]
    wire [63:0]     _GEN_4974; // @[ISA.scala 328:101:@165508.12]
    wire [31:0]     _GEN_4975; // @[ISA.scala 328:101:@165508.12]
    wire [31:0]     _GEN_4976; // @[ISA.scala 328:101:@165508.12]
    wire [31:0]     _GEN_4977; // @[ISA.scala 328:101:@165508.12]
    wire [31:0]     _GEN_4978; // @[ISA.scala 328:101:@165508.12]
    wire [31:0]     _GEN_4979; // @[ISA.scala 328:101:@165508.12]
    wire [63:0]     _GEN_4980; // @[ISA.scala 328:101:@165508.12]
    wire [63:0]     _GEN_4981; // @[ISA.scala 328:101:@165508.12]
    wire [31:0]     _GEN_4982; // @[ISA.scala 328:101:@165508.12]
    wire [31:0]     _GEN_4983; // @[ISA.scala 328:101:@165508.12]
    wire [31:0]     _GEN_4984; // @[ISA.scala 328:101:@165508.12]
    wire [31:0]     _GEN_4985; // @[ISA.scala 328:101:@165508.12]
    wire [63:0]     _GEN_4986; // @[ISA.scala 328:101:@165508.12]
    wire            _GEN_4987; // @[ISA.scala 328:101:@165508.12]
    wire            _GEN_4988; // @[ISA.scala 328:101:@165508.12]
    wire            _GEN_4989; // @[ISA.scala 328:101:@165508.12]
    wire [2:0]      _GEN_4990; // @[ISA.scala 327:93:@165336.10]
    wire [63:0]     _GEN_4991; // @[ISA.scala 327:93:@165336.10]
    wire [31:0]     _GEN_4992; // @[ISA.scala 327:93:@165336.10]
    wire [31:0]     _GEN_4993; // @[ISA.scala 327:93:@165336.10]
    wire [31:0]     _GEN_4994; // @[ISA.scala 327:93:@165336.10]
    wire [31:0]     _GEN_4995; // @[ISA.scala 327:93:@165336.10]
    wire [31:0]     _GEN_4996; // @[ISA.scala 327:93:@165336.10]
    wire [63:0]     _GEN_4997; // @[ISA.scala 327:93:@165336.10]
    wire [63:0]     _GEN_4998; // @[ISA.scala 327:93:@165336.10]
    wire [31:0]     _GEN_4999; // @[ISA.scala 327:93:@165336.10]
    wire [31:0]     _GEN_5000; // @[ISA.scala 327:93:@165336.10]
    wire [31:0]     _GEN_5001; // @[ISA.scala 327:93:@165336.10]
    wire [31:0]     _GEN_5002; // @[ISA.scala 327:93:@165336.10]
    wire [63:0]     _GEN_5003; // @[ISA.scala 327:93:@165336.10]
    wire            _GEN_5004; // @[ISA.scala 327:93:@165336.10]
    wire            _GEN_5005; // @[ISA.scala 327:93:@165336.10]
    wire            _GEN_5006; // @[ISA.scala 327:93:@165336.10]
    wire [2:0]      _GEN_5007; // @[ISA.scala 326:85:@165164.8]
    wire [63:0]     _GEN_5008; // @[ISA.scala 326:85:@165164.8]
    wire [31:0]     _GEN_5009; // @[ISA.scala 326:85:@165164.8]
    wire [31:0]     _GEN_5010; // @[ISA.scala 326:85:@165164.8]
    wire [31:0]     _GEN_5011; // @[ISA.scala 326:85:@165164.8]
    wire [31:0]     _GEN_5012; // @[ISA.scala 326:85:@165164.8]
    wire [31:0]     _GEN_5013; // @[ISA.scala 326:85:@165164.8]
    wire [63:0]     _GEN_5014; // @[ISA.scala 326:85:@165164.8]
    wire [63:0]     _GEN_5015; // @[ISA.scala 326:85:@165164.8]
    wire [31:0]     _GEN_5016; // @[ISA.scala 326:85:@165164.8]
    wire [31:0]     _GEN_5017; // @[ISA.scala 326:85:@165164.8]
    wire [31:0]     _GEN_5018; // @[ISA.scala 326:85:@165164.8]
    wire [31:0]     _GEN_5019; // @[ISA.scala 326:85:@165164.8]
    wire [63:0]     _GEN_5020; // @[ISA.scala 326:85:@165164.8]
    wire            _GEN_5021; // @[ISA.scala 326:85:@165164.8]
    wire            _GEN_5022; // @[ISA.scala 326:85:@165164.8]
    wire            _GEN_5023; // @[ISA.scala 326:85:@165164.8]
    wire [2:0]      _GEN_5024; // @[ISA.scala 325:44:@164992.6]
    wire [63:0]     _GEN_5025; // @[ISA.scala 325:44:@164992.6]
    wire [31:0]     _GEN_5026; // @[ISA.scala 325:44:@164992.6]
    wire [31:0]     _GEN_5027; // @[ISA.scala 325:44:@164992.6]
    wire [31:0]     _GEN_5028; // @[ISA.scala 325:44:@164992.6]
    wire [31:0]     _GEN_5029; // @[ISA.scala 325:44:@164992.6]
    wire [31:0]     _GEN_5030; // @[ISA.scala 325:44:@164992.6]
    wire [63:0]     _GEN_5031; // @[ISA.scala 325:44:@164992.6]
    wire [63:0]     _GEN_5032; // @[ISA.scala 325:44:@164992.6]
    wire [31:0]     _GEN_5033; // @[ISA.scala 325:44:@164992.6]
    wire [31:0]     _GEN_5034; // @[ISA.scala 325:44:@164992.6]
    wire [31:0]     _GEN_5035; // @[ISA.scala 325:44:@164992.6]
    wire [31:0]     _GEN_5036; // @[ISA.scala 325:44:@164992.6]
    wire [63:0]     _GEN_5037; // @[ISA.scala 325:44:@164992.6]
    wire            _GEN_5038; // @[ISA.scala 325:44:@164992.6]
    wire            _GEN_5039; // @[ISA.scala 325:44:@164992.6]
    wire            _GEN_5040; // @[ISA.scala 325:44:@164992.6]
    wire            _T_257102; // @[ISA_functions.scala 176:203:@172339.32]
    wire            _T_257130; // @[ISA_functions.scala 179:203:@172364.34]
    wire            _T_257158; // @[ISA_functions.scala 182:234:@172389.36]
    wire            _T_257188; // @[ISA_functions.scala 185:234:@172415.38]
    wire [31:0]     _GEN_5189; // @[ISA_functions.scala 194:325:@172511.44]
    wire [31:0]     _GEN_5190; // @[ISA_functions.scala 191:295:@172475.42]
    wire [31:0]     _GEN_5191; // @[ISA_functions.scala 188:265:@172442.40]
    wire [31:0]     _GEN_5192; // @[ISA_functions.scala 185:261:@172416.38]
    wire [31:0]     _GEN_5193; // @[ISA_functions.scala 182:260:@172390.36]
    wire [31:0]     _GEN_5194; // @[ISA_functions.scala 179:248:@172365.34]
    wire [31:0]     _GEN_5195; // @[ISA_functions.scala 176:247:@172340.32]
    wire [31:0]     _GEN_5196; // @[ISA_functions.scala 173:174:@172315.30]
    wire [31:0]     _GEN_5197; // @[ISA_functions.scala 170:144:@172297.28]
    wire [31:0]     _GEN_5198; // @[ISA_functions.scala 167:115:@172282.26]
    wire [63:0]     _GEN_5199; // @[ISA_functions.scala 164:85:@172268.24]
    wire [63:0]     _GEN_5200; // @[ISA_functions.scala 161:50:@172258.22]
    wire [2:0]      _GEN_5313; // @[ISA.scala 363:102:@167880.20]
    wire [63:0]     _GEN_5314; // @[ISA.scala 363:102:@167880.20]
    wire [31:0]     _GEN_5315; // @[ISA.scala 363:102:@167880.20]
    wire [31:0]     _GEN_5316; // @[ISA.scala 363:102:@167880.20]
    wire [31:0]     _GEN_5317; // @[ISA.scala 363:102:@167880.20]
    wire [31:0]     _GEN_5318; // @[ISA.scala 363:102:@167880.20]
    wire [31:0]     _GEN_5319; // @[ISA.scala 363:102:@167880.20]
    wire [63:0]     _GEN_5320; // @[ISA.scala 363:102:@167880.20]
    wire [63:0]     _GEN_5321; // @[ISA.scala 363:102:@167880.20]
    wire [31:0]     _GEN_5322; // @[ISA.scala 363:102:@167880.20]
    wire [31:0]     _GEN_5323; // @[ISA.scala 363:102:@167880.20]
    wire [31:0]     _GEN_5324; // @[ISA.scala 363:102:@167880.20]
    wire [31:0]     _GEN_5325; // @[ISA.scala 363:102:@167880.20]
    wire [63:0]     _GEN_5326; // @[ISA.scala 363:102:@167880.20]
    wire            _GEN_5327; // @[ISA.scala 363:102:@167880.20]
    wire            _GEN_5328; // @[ISA.scala 363:102:@167880.20]
    wire            _GEN_5329; // @[ISA.scala 363:102:@167880.20]
    wire [2:0]      _GEN_5330; // @[ISA.scala 362:126:@167879.18]
    wire [63:0]     _GEN_5331; // @[ISA.scala 362:126:@167879.18]
    wire [31:0]     _GEN_5332; // @[ISA.scala 362:126:@167879.18]
    wire [31:0]     _GEN_5333; // @[ISA.scala 362:126:@167879.18]
    wire [31:0]     _GEN_5334; // @[ISA.scala 362:126:@167879.18]
    wire [31:0]     _GEN_5335; // @[ISA.scala 362:126:@167879.18]
    wire [31:0]     _GEN_5336; // @[ISA.scala 362:126:@167879.18]
    wire [63:0]     _GEN_5337; // @[ISA.scala 362:126:@167879.18]
    wire [63:0]     _GEN_5338; // @[ISA.scala 362:126:@167879.18]
    wire [31:0]     _GEN_5339; // @[ISA.scala 362:126:@167879.18]
    wire [31:0]     _GEN_5340; // @[ISA.scala 362:126:@167879.18]
    wire [31:0]     _GEN_5341; // @[ISA.scala 362:126:@167879.18]
    wire [31:0]     _GEN_5342; // @[ISA.scala 362:126:@167879.18]
    wire [63:0]     _GEN_5343; // @[ISA.scala 362:126:@167879.18]
    wire            _GEN_5344; // @[ISA.scala 362:126:@167879.18]
    wire            _GEN_5345; // @[ISA.scala 362:126:@167879.18]
    wire            _GEN_5346; // @[ISA.scala 362:126:@167879.18]
    wire [2:0]      _GEN_5347; // @[ISA.scala 361:117:@167708.16]
    wire [63:0]     _GEN_5348; // @[ISA.scala 361:117:@167708.16]
    wire [31:0]     _GEN_5349; // @[ISA.scala 361:117:@167708.16]
    wire [31:0]     _GEN_5350; // @[ISA.scala 361:117:@167708.16]
    wire [31:0]     _GEN_5351; // @[ISA.scala 361:117:@167708.16]
    wire [31:0]     _GEN_5352; // @[ISA.scala 361:117:@167708.16]
    wire [31:0]     _GEN_5353; // @[ISA.scala 361:117:@167708.16]
    wire [63:0]     _GEN_5354; // @[ISA.scala 361:117:@167708.16]
    wire [63:0]     _GEN_5355; // @[ISA.scala 361:117:@167708.16]
    wire [31:0]     _GEN_5356; // @[ISA.scala 361:117:@167708.16]
    wire [31:0]     _GEN_5357; // @[ISA.scala 361:117:@167708.16]
    wire [31:0]     _GEN_5358; // @[ISA.scala 361:117:@167708.16]
    wire [31:0]     _GEN_5359; // @[ISA.scala 361:117:@167708.16]
    wire [63:0]     _GEN_5360; // @[ISA.scala 361:117:@167708.16]
    wire            _GEN_5361; // @[ISA.scala 361:117:@167708.16]
    wire            _GEN_5362; // @[ISA.scala 361:117:@167708.16]
    wire            _GEN_5363; // @[ISA.scala 361:117:@167708.16]
    wire [2:0]      _GEN_5364; // @[ISA.scala 360:109:@167536.14]
    wire [63:0]     _GEN_5365; // @[ISA.scala 360:109:@167536.14]
    wire [31:0]     _GEN_5366; // @[ISA.scala 360:109:@167536.14]
    wire [31:0]     _GEN_5367; // @[ISA.scala 360:109:@167536.14]
    wire [31:0]     _GEN_5368; // @[ISA.scala 360:109:@167536.14]
    wire [31:0]     _GEN_5369; // @[ISA.scala 360:109:@167536.14]
    wire [31:0]     _GEN_5370; // @[ISA.scala 360:109:@167536.14]
    wire [63:0]     _GEN_5371; // @[ISA.scala 360:109:@167536.14]
    wire [63:0]     _GEN_5372; // @[ISA.scala 360:109:@167536.14]
    wire [31:0]     _GEN_5373; // @[ISA.scala 360:109:@167536.14]
    wire [31:0]     _GEN_5374; // @[ISA.scala 360:109:@167536.14]
    wire [31:0]     _GEN_5375; // @[ISA.scala 360:109:@167536.14]
    wire [31:0]     _GEN_5376; // @[ISA.scala 360:109:@167536.14]
    wire [63:0]     _GEN_5377; // @[ISA.scala 360:109:@167536.14]
    wire            _GEN_5378; // @[ISA.scala 360:109:@167536.14]
    wire            _GEN_5379; // @[ISA.scala 360:109:@167536.14]
    wire            _GEN_5380; // @[ISA.scala 360:109:@167536.14]
    wire [2:0]      _GEN_5381; // @[ISA.scala 359:101:@167364.12]
    wire [63:0]     _GEN_5382; // @[ISA.scala 359:101:@167364.12]
    wire [31:0]     _GEN_5383; // @[ISA.scala 359:101:@167364.12]
    wire [31:0]     _GEN_5384; // @[ISA.scala 359:101:@167364.12]
    wire [31:0]     _GEN_5385; // @[ISA.scala 359:101:@167364.12]
    wire [31:0]     _GEN_5386; // @[ISA.scala 359:101:@167364.12]
    wire [31:0]     _GEN_5387; // @[ISA.scala 359:101:@167364.12]
    wire [63:0]     _GEN_5388; // @[ISA.scala 359:101:@167364.12]
    wire [63:0]     _GEN_5389; // @[ISA.scala 359:101:@167364.12]
    wire [31:0]     _GEN_5390; // @[ISA.scala 359:101:@167364.12]
    wire [31:0]     _GEN_5391; // @[ISA.scala 359:101:@167364.12]
    wire [31:0]     _GEN_5392; // @[ISA.scala 359:101:@167364.12]
    wire [31:0]     _GEN_5393; // @[ISA.scala 359:101:@167364.12]
    wire [63:0]     _GEN_5394; // @[ISA.scala 359:101:@167364.12]
    wire            _GEN_5395; // @[ISA.scala 359:101:@167364.12]
    wire            _GEN_5396; // @[ISA.scala 359:101:@167364.12]
    wire            _GEN_5397; // @[ISA.scala 359:101:@167364.12]
    wire [2:0]      _GEN_5398; // @[ISA.scala 358:93:@167192.10]
    wire [63:0]     _GEN_5399; // @[ISA.scala 358:93:@167192.10]
    wire [31:0]     _GEN_5400; // @[ISA.scala 358:93:@167192.10]
    wire [31:0]     _GEN_5401; // @[ISA.scala 358:93:@167192.10]
    wire [31:0]     _GEN_5402; // @[ISA.scala 358:93:@167192.10]
    wire [31:0]     _GEN_5403; // @[ISA.scala 358:93:@167192.10]
    wire [31:0]     _GEN_5404; // @[ISA.scala 358:93:@167192.10]
    wire [63:0]     _GEN_5405; // @[ISA.scala 358:93:@167192.10]
    wire [63:0]     _GEN_5406; // @[ISA.scala 358:93:@167192.10]
    wire [31:0]     _GEN_5407; // @[ISA.scala 358:93:@167192.10]
    wire [31:0]     _GEN_5408; // @[ISA.scala 358:93:@167192.10]
    wire [31:0]     _GEN_5409; // @[ISA.scala 358:93:@167192.10]
    wire [31:0]     _GEN_5410; // @[ISA.scala 358:93:@167192.10]
    wire [63:0]     _GEN_5411; // @[ISA.scala 358:93:@167192.10]
    wire            _GEN_5412; // @[ISA.scala 358:93:@167192.10]
    wire            _GEN_5413; // @[ISA.scala 358:93:@167192.10]
    wire            _GEN_5414; // @[ISA.scala 358:93:@167192.10]
    wire [2:0]      _GEN_5415; // @[ISA.scala 357:85:@167020.8]
    wire [63:0]     _GEN_5416; // @[ISA.scala 357:85:@167020.8]
    wire [31:0]     _GEN_5417; // @[ISA.scala 357:85:@167020.8]
    wire [31:0]     _GEN_5418; // @[ISA.scala 357:85:@167020.8]
    wire [31:0]     _GEN_5419; // @[ISA.scala 357:85:@167020.8]
    wire [31:0]     _GEN_5420; // @[ISA.scala 357:85:@167020.8]
    wire [31:0]     _GEN_5421; // @[ISA.scala 357:85:@167020.8]
    wire [63:0]     _GEN_5422; // @[ISA.scala 357:85:@167020.8]
    wire [63:0]     _GEN_5423; // @[ISA.scala 357:85:@167020.8]
    wire [31:0]     _GEN_5424; // @[ISA.scala 357:85:@167020.8]
    wire [31:0]     _GEN_5425; // @[ISA.scala 357:85:@167020.8]
    wire [31:0]     _GEN_5426; // @[ISA.scala 357:85:@167020.8]
    wire [31:0]     _GEN_5427; // @[ISA.scala 357:85:@167020.8]
    wire [63:0]     _GEN_5428; // @[ISA.scala 357:85:@167020.8]
    wire            _GEN_5429; // @[ISA.scala 357:85:@167020.8]
    wire            _GEN_5430; // @[ISA.scala 357:85:@167020.8]
    wire            _GEN_5431; // @[ISA.scala 357:85:@167020.8]
    wire [2:0]      _GEN_5432; // @[ISA.scala 356:44:@166848.6]
    wire [63:0]     _GEN_5433; // @[ISA.scala 356:44:@166848.6]
    wire [31:0]     _GEN_5434; // @[ISA.scala 356:44:@166848.6]
    wire [31:0]     _GEN_5435; // @[ISA.scala 356:44:@166848.6]
    wire [31:0]     _GEN_5436; // @[ISA.scala 356:44:@166848.6]
    wire [31:0]     _GEN_5437; // @[ISA.scala 356:44:@166848.6]
    wire [31:0]     _GEN_5438; // @[ISA.scala 356:44:@166848.6]
    wire [63:0]     _GEN_5439; // @[ISA.scala 356:44:@166848.6]
    wire [63:0]     _GEN_5440; // @[ISA.scala 356:44:@166848.6]
    wire [31:0]     _GEN_5441; // @[ISA.scala 356:44:@166848.6]
    wire [31:0]     _GEN_5442; // @[ISA.scala 356:44:@166848.6]
    wire [31:0]     _GEN_5443; // @[ISA.scala 356:44:@166848.6]
    wire [31:0]     _GEN_5444; // @[ISA.scala 356:44:@166848.6]
    wire [63:0]     _GEN_5445; // @[ISA.scala 356:44:@166848.6]
    wire            _GEN_5446; // @[ISA.scala 356:44:@166848.6]
    wire            _GEN_5447; // @[ISA.scala 356:44:@166848.6]
    wire            _GEN_5448; // @[ISA.scala 356:44:@166848.6]
    wire [2:0]      _GEN_5714; // @[ISA.scala 397:110:@178443.22]
    wire [63:0]     _GEN_5715; // @[ISA.scala 397:110:@178443.22]
    wire [31:0]     _GEN_5716; // @[ISA.scala 397:110:@178443.22]
    wire [31:0]     _GEN_5717; // @[ISA.scala 397:110:@178443.22]
    wire [31:0]     _GEN_5718; // @[ISA.scala 397:110:@178443.22]
    wire [31:0]     _GEN_5719; // @[ISA.scala 397:110:@178443.22]
    wire [31:0]     _GEN_5720; // @[ISA.scala 397:110:@178443.22]
    wire [63:0]     _GEN_5721; // @[ISA.scala 397:110:@178443.22]
    wire [63:0]     _GEN_5722; // @[ISA.scala 397:110:@178443.22]
    wire [31:0]     _GEN_5723; // @[ISA.scala 397:110:@178443.22]
    wire [31:0]     _GEN_5724; // @[ISA.scala 397:110:@178443.22]
    wire [31:0]     _GEN_5725; // @[ISA.scala 397:110:@178443.22]
    wire            _GEN_5726; // @[ISA.scala 397:110:@178443.22]
    wire            _GEN_5727; // @[ISA.scala 397:110:@178443.22]
    wire            _GEN_5728; // @[ISA.scala 397:110:@178443.22]
    wire [2:0]      _GEN_5729; // @[ISA.scala 396:134:@178442.20]
    wire [63:0]     _GEN_5730; // @[ISA.scala 396:134:@178442.20]
    wire [31:0]     _GEN_5731; // @[ISA.scala 396:134:@178442.20]
    wire [31:0]     _GEN_5732; // @[ISA.scala 396:134:@178442.20]
    wire [31:0]     _GEN_5733; // @[ISA.scala 396:134:@178442.20]
    wire [31:0]     _GEN_5734; // @[ISA.scala 396:134:@178442.20]
    wire [31:0]     _GEN_5735; // @[ISA.scala 396:134:@178442.20]
    wire [63:0]     _GEN_5736; // @[ISA.scala 396:134:@178442.20]
    wire [63:0]     _GEN_5737; // @[ISA.scala 396:134:@178442.20]
    wire [31:0]     _GEN_5738; // @[ISA.scala 396:134:@178442.20]
    wire [31:0]     _GEN_5739; // @[ISA.scala 396:134:@178442.20]
    wire [31:0]     _GEN_5740; // @[ISA.scala 396:134:@178442.20]
    wire            _GEN_5741; // @[ISA.scala 396:134:@178442.20]
    wire            _GEN_5742; // @[ISA.scala 396:134:@178442.20]
    wire            _GEN_5743; // @[ISA.scala 396:134:@178442.20]
    wire [2:0]      _GEN_5744; // @[ISA.scala 395:127:@178271.18]
    wire [63:0]     _GEN_5745; // @[ISA.scala 395:127:@178271.18]
    wire [31:0]     _GEN_5746; // @[ISA.scala 395:127:@178271.18]
    wire [31:0]     _GEN_5747; // @[ISA.scala 395:127:@178271.18]
    wire [31:0]     _GEN_5748; // @[ISA.scala 395:127:@178271.18]
    wire [31:0]     _GEN_5749; // @[ISA.scala 395:127:@178271.18]
    wire [31:0]     _GEN_5750; // @[ISA.scala 395:127:@178271.18]
    wire [63:0]     _GEN_5751; // @[ISA.scala 395:127:@178271.18]
    wire [63:0]     _GEN_5752; // @[ISA.scala 395:127:@178271.18]
    wire [31:0]     _GEN_5753; // @[ISA.scala 395:127:@178271.18]
    wire [31:0]     _GEN_5754; // @[ISA.scala 395:127:@178271.18]
    wire [31:0]     _GEN_5755; // @[ISA.scala 395:127:@178271.18]
    wire            _GEN_5756; // @[ISA.scala 395:127:@178271.18]
    wire            _GEN_5757; // @[ISA.scala 395:127:@178271.18]
    wire            _GEN_5758; // @[ISA.scala 395:127:@178271.18]
    wire [2:0]      _GEN_5759; // @[ISA.scala 394:117:@178099.16]
    wire [63:0]     _GEN_5760; // @[ISA.scala 394:117:@178099.16]
    wire [31:0]     _GEN_5761; // @[ISA.scala 394:117:@178099.16]
    wire [31:0]     _GEN_5762; // @[ISA.scala 394:117:@178099.16]
    wire [31:0]     _GEN_5763; // @[ISA.scala 394:117:@178099.16]
    wire [31:0]     _GEN_5764; // @[ISA.scala 394:117:@178099.16]
    wire [31:0]     _GEN_5765; // @[ISA.scala 394:117:@178099.16]
    wire [63:0]     _GEN_5766; // @[ISA.scala 394:117:@178099.16]
    wire [63:0]     _GEN_5767; // @[ISA.scala 394:117:@178099.16]
    wire [31:0]     _GEN_5768; // @[ISA.scala 394:117:@178099.16]
    wire [31:0]     _GEN_5769; // @[ISA.scala 394:117:@178099.16]
    wire [31:0]     _GEN_5770; // @[ISA.scala 394:117:@178099.16]
    wire            _GEN_5771; // @[ISA.scala 394:117:@178099.16]
    wire            _GEN_5772; // @[ISA.scala 394:117:@178099.16]
    wire            _GEN_5773; // @[ISA.scala 394:117:@178099.16]
    wire [2:0]      _GEN_5774; // @[ISA.scala 393:109:@177927.14]
    wire [63:0]     _GEN_5775; // @[ISA.scala 393:109:@177927.14]
    wire [31:0]     _GEN_5776; // @[ISA.scala 393:109:@177927.14]
    wire [31:0]     _GEN_5777; // @[ISA.scala 393:109:@177927.14]
    wire [31:0]     _GEN_5778; // @[ISA.scala 393:109:@177927.14]
    wire [31:0]     _GEN_5779; // @[ISA.scala 393:109:@177927.14]
    wire [31:0]     _GEN_5780; // @[ISA.scala 393:109:@177927.14]
    wire [63:0]     _GEN_5781; // @[ISA.scala 393:109:@177927.14]
    wire [63:0]     _GEN_5782; // @[ISA.scala 393:109:@177927.14]
    wire [31:0]     _GEN_5783; // @[ISA.scala 393:109:@177927.14]
    wire [31:0]     _GEN_5784; // @[ISA.scala 393:109:@177927.14]
    wire [31:0]     _GEN_5785; // @[ISA.scala 393:109:@177927.14]
    wire            _GEN_5786; // @[ISA.scala 393:109:@177927.14]
    wire            _GEN_5787; // @[ISA.scala 393:109:@177927.14]
    wire            _GEN_5788; // @[ISA.scala 393:109:@177927.14]
    wire [2:0]      _GEN_5789; // @[ISA.scala 392:101:@177755.12]
    wire [63:0]     _GEN_5790; // @[ISA.scala 392:101:@177755.12]
    wire [31:0]     _GEN_5791; // @[ISA.scala 392:101:@177755.12]
    wire [31:0]     _GEN_5792; // @[ISA.scala 392:101:@177755.12]
    wire [31:0]     _GEN_5793; // @[ISA.scala 392:101:@177755.12]
    wire [31:0]     _GEN_5794; // @[ISA.scala 392:101:@177755.12]
    wire [31:0]     _GEN_5795; // @[ISA.scala 392:101:@177755.12]
    wire [63:0]     _GEN_5796; // @[ISA.scala 392:101:@177755.12]
    wire [63:0]     _GEN_5797; // @[ISA.scala 392:101:@177755.12]
    wire [31:0]     _GEN_5798; // @[ISA.scala 392:101:@177755.12]
    wire [31:0]     _GEN_5799; // @[ISA.scala 392:101:@177755.12]
    wire [31:0]     _GEN_5800; // @[ISA.scala 392:101:@177755.12]
    wire            _GEN_5801; // @[ISA.scala 392:101:@177755.12]
    wire            _GEN_5802; // @[ISA.scala 392:101:@177755.12]
    wire            _GEN_5803; // @[ISA.scala 392:101:@177755.12]
    wire [2:0]      _GEN_5804; // @[ISA.scala 391:93:@177583.10]
    wire [63:0]     _GEN_5805; // @[ISA.scala 391:93:@177583.10]
    wire [31:0]     _GEN_5806; // @[ISA.scala 391:93:@177583.10]
    wire [31:0]     _GEN_5807; // @[ISA.scala 391:93:@177583.10]
    wire [31:0]     _GEN_5808; // @[ISA.scala 391:93:@177583.10]
    wire [31:0]     _GEN_5809; // @[ISA.scala 391:93:@177583.10]
    wire [31:0]     _GEN_5810; // @[ISA.scala 391:93:@177583.10]
    wire [63:0]     _GEN_5811; // @[ISA.scala 391:93:@177583.10]
    wire [63:0]     _GEN_5812; // @[ISA.scala 391:93:@177583.10]
    wire [31:0]     _GEN_5813; // @[ISA.scala 391:93:@177583.10]
    wire [31:0]     _GEN_5814; // @[ISA.scala 391:93:@177583.10]
    wire [31:0]     _GEN_5815; // @[ISA.scala 391:93:@177583.10]
    wire            _GEN_5816; // @[ISA.scala 391:93:@177583.10]
    wire            _GEN_5817; // @[ISA.scala 391:93:@177583.10]
    wire            _GEN_5818; // @[ISA.scala 391:93:@177583.10]
    wire [2:0]      _GEN_5819; // @[ISA.scala 390:85:@177411.8]
    wire [63:0]     _GEN_5820; // @[ISA.scala 390:85:@177411.8]
    wire [31:0]     _GEN_5821; // @[ISA.scala 390:85:@177411.8]
    wire [31:0]     _GEN_5822; // @[ISA.scala 390:85:@177411.8]
    wire [31:0]     _GEN_5823; // @[ISA.scala 390:85:@177411.8]
    wire [31:0]     _GEN_5824; // @[ISA.scala 390:85:@177411.8]
    wire [31:0]     _GEN_5825; // @[ISA.scala 390:85:@177411.8]
    wire [63:0]     _GEN_5826; // @[ISA.scala 390:85:@177411.8]
    wire [63:0]     _GEN_5827; // @[ISA.scala 390:85:@177411.8]
    wire [31:0]     _GEN_5828; // @[ISA.scala 390:85:@177411.8]
    wire [31:0]     _GEN_5829; // @[ISA.scala 390:85:@177411.8]
    wire [31:0]     _GEN_5830; // @[ISA.scala 390:85:@177411.8]
    wire            _GEN_5831; // @[ISA.scala 390:85:@177411.8]
    wire            _GEN_5832; // @[ISA.scala 390:85:@177411.8]
    wire            _GEN_5833; // @[ISA.scala 390:85:@177411.8]
    wire [2:0]      _GEN_5834; // @[ISA.scala 389:44:@177239.6]
    wire [63:0]     _GEN_5835; // @[ISA.scala 389:44:@177239.6]
    wire [31:0]     _GEN_5836; // @[ISA.scala 389:44:@177239.6]
    wire [31:0]     _GEN_5837; // @[ISA.scala 389:44:@177239.6]
    wire [31:0]     _GEN_5838; // @[ISA.scala 389:44:@177239.6]
    wire [31:0]     _GEN_5839; // @[ISA.scala 389:44:@177239.6]
    wire [31:0]     _GEN_5840; // @[ISA.scala 389:44:@177239.6]
    wire [63:0]     _GEN_5841; // @[ISA.scala 389:44:@177239.6]
    wire [63:0]     _GEN_5842; // @[ISA.scala 389:44:@177239.6]
    wire [31:0]     _GEN_5843; // @[ISA.scala 389:44:@177239.6]
    wire [31:0]     _GEN_5844; // @[ISA.scala 389:44:@177239.6]
    wire [31:0]     _GEN_5845; // @[ISA.scala 389:44:@177239.6]
    wire            _GEN_5846; // @[ISA.scala 389:44:@177239.6]
    wire            _GEN_5847; // @[ISA.scala 389:44:@177239.6]
    wire            _GEN_5848; // @[ISA.scala 389:44:@177239.6]
    wire [2:0]      _GEN_6038; // @[ISA.scala 431:118:@187863.24]
    wire [63:0]     _GEN_6039; // @[ISA.scala 431:118:@187863.24]
    wire [31:0]     _GEN_6040; // @[ISA.scala 431:118:@187863.24]
    wire [31:0]     _GEN_6041; // @[ISA.scala 431:118:@187863.24]
    wire [31:0]     _GEN_6042; // @[ISA.scala 431:118:@187863.24]
    wire [31:0]     _GEN_6043; // @[ISA.scala 431:118:@187863.24]
    wire [31:0]     _GEN_6044; // @[ISA.scala 431:118:@187863.24]
    wire [63:0]     _GEN_6045; // @[ISA.scala 431:118:@187863.24]
    wire [63:0]     _GEN_6046; // @[ISA.scala 431:118:@187863.24]
    wire [31:0]     _GEN_6047; // @[ISA.scala 431:118:@187863.24]
    wire [31:0]     _GEN_6048; // @[ISA.scala 431:118:@187863.24]
    wire [31:0]     _GEN_6049; // @[ISA.scala 431:118:@187863.24]
    wire [31:0]     _GEN_6050; // @[ISA.scala 431:118:@187863.24]
    wire [63:0]     _GEN_6051; // @[ISA.scala 431:118:@187863.24]
    wire            _GEN_6052; // @[ISA.scala 431:118:@187863.24]
    wire            _GEN_6053; // @[ISA.scala 431:118:@187863.24]
    wire            _GEN_6054; // @[ISA.scala 431:118:@187863.24]
    wire [2:0]      _GEN_6055; // @[ISA.scala 430:142:@187862.22]
    wire [63:0]     _GEN_6056; // @[ISA.scala 430:142:@187862.22]
    wire [31:0]     _GEN_6057; // @[ISA.scala 430:142:@187862.22]
    wire [31:0]     _GEN_6058; // @[ISA.scala 430:142:@187862.22]
    wire [31:0]     _GEN_6059; // @[ISA.scala 430:142:@187862.22]
    wire [31:0]     _GEN_6060; // @[ISA.scala 430:142:@187862.22]
    wire [31:0]     _GEN_6061; // @[ISA.scala 430:142:@187862.22]
    wire [63:0]     _GEN_6062; // @[ISA.scala 430:142:@187862.22]
    wire [63:0]     _GEN_6063; // @[ISA.scala 430:142:@187862.22]
    wire [31:0]     _GEN_6064; // @[ISA.scala 430:142:@187862.22]
    wire [31:0]     _GEN_6065; // @[ISA.scala 430:142:@187862.22]
    wire [31:0]     _GEN_6066; // @[ISA.scala 430:142:@187862.22]
    wire [31:0]     _GEN_6067; // @[ISA.scala 430:142:@187862.22]
    wire [63:0]     _GEN_6068; // @[ISA.scala 430:142:@187862.22]
    wire            _GEN_6069; // @[ISA.scala 430:142:@187862.22]
    wire            _GEN_6070; // @[ISA.scala 430:142:@187862.22]
    wire            _GEN_6071; // @[ISA.scala 430:142:@187862.22]
    wire [2:0]      _GEN_6072; // @[ISA.scala 429:135:@187691.20]
    wire [63:0]     _GEN_6073; // @[ISA.scala 429:135:@187691.20]
    wire [31:0]     _GEN_6074; // @[ISA.scala 429:135:@187691.20]
    wire [31:0]     _GEN_6075; // @[ISA.scala 429:135:@187691.20]
    wire [31:0]     _GEN_6076; // @[ISA.scala 429:135:@187691.20]
    wire [31:0]     _GEN_6077; // @[ISA.scala 429:135:@187691.20]
    wire [31:0]     _GEN_6078; // @[ISA.scala 429:135:@187691.20]
    wire [63:0]     _GEN_6079; // @[ISA.scala 429:135:@187691.20]
    wire [63:0]     _GEN_6080; // @[ISA.scala 429:135:@187691.20]
    wire [31:0]     _GEN_6081; // @[ISA.scala 429:135:@187691.20]
    wire [31:0]     _GEN_6082; // @[ISA.scala 429:135:@187691.20]
    wire [31:0]     _GEN_6083; // @[ISA.scala 429:135:@187691.20]
    wire [31:0]     _GEN_6084; // @[ISA.scala 429:135:@187691.20]
    wire [63:0]     _GEN_6085; // @[ISA.scala 429:135:@187691.20]
    wire            _GEN_6086; // @[ISA.scala 429:135:@187691.20]
    wire            _GEN_6087; // @[ISA.scala 429:135:@187691.20]
    wire            _GEN_6088; // @[ISA.scala 429:135:@187691.20]
    wire [2:0]      _GEN_6089; // @[ISA.scala 428:127:@187519.18]
    wire [63:0]     _GEN_6090; // @[ISA.scala 428:127:@187519.18]
    wire [31:0]     _GEN_6091; // @[ISA.scala 428:127:@187519.18]
    wire [31:0]     _GEN_6092; // @[ISA.scala 428:127:@187519.18]
    wire [31:0]     _GEN_6093; // @[ISA.scala 428:127:@187519.18]
    wire [31:0]     _GEN_6094; // @[ISA.scala 428:127:@187519.18]
    wire [31:0]     _GEN_6095; // @[ISA.scala 428:127:@187519.18]
    wire [63:0]     _GEN_6096; // @[ISA.scala 428:127:@187519.18]
    wire [63:0]     _GEN_6097; // @[ISA.scala 428:127:@187519.18]
    wire [31:0]     _GEN_6098; // @[ISA.scala 428:127:@187519.18]
    wire [31:0]     _GEN_6099; // @[ISA.scala 428:127:@187519.18]
    wire [31:0]     _GEN_6100; // @[ISA.scala 428:127:@187519.18]
    wire [31:0]     _GEN_6101; // @[ISA.scala 428:127:@187519.18]
    wire [63:0]     _GEN_6102; // @[ISA.scala 428:127:@187519.18]
    wire            _GEN_6103; // @[ISA.scala 428:127:@187519.18]
    wire            _GEN_6104; // @[ISA.scala 428:127:@187519.18]
    wire            _GEN_6105; // @[ISA.scala 428:127:@187519.18]
    wire [2:0]      _GEN_6106; // @[ISA.scala 427:117:@187347.16]
    wire [63:0]     _GEN_6107; // @[ISA.scala 427:117:@187347.16]
    wire [31:0]     _GEN_6108; // @[ISA.scala 427:117:@187347.16]
    wire [31:0]     _GEN_6109; // @[ISA.scala 427:117:@187347.16]
    wire [31:0]     _GEN_6110; // @[ISA.scala 427:117:@187347.16]
    wire [31:0]     _GEN_6111; // @[ISA.scala 427:117:@187347.16]
    wire [31:0]     _GEN_6112; // @[ISA.scala 427:117:@187347.16]
    wire [63:0]     _GEN_6113; // @[ISA.scala 427:117:@187347.16]
    wire [63:0]     _GEN_6114; // @[ISA.scala 427:117:@187347.16]
    wire [31:0]     _GEN_6115; // @[ISA.scala 427:117:@187347.16]
    wire [31:0]     _GEN_6116; // @[ISA.scala 427:117:@187347.16]
    wire [31:0]     _GEN_6117; // @[ISA.scala 427:117:@187347.16]
    wire [31:0]     _GEN_6118; // @[ISA.scala 427:117:@187347.16]
    wire [63:0]     _GEN_6119; // @[ISA.scala 427:117:@187347.16]
    wire            _GEN_6120; // @[ISA.scala 427:117:@187347.16]
    wire            _GEN_6121; // @[ISA.scala 427:117:@187347.16]
    wire            _GEN_6122; // @[ISA.scala 427:117:@187347.16]
    wire [2:0]      _GEN_6123; // @[ISA.scala 426:109:@187175.14]
    wire [63:0]     _GEN_6124; // @[ISA.scala 426:109:@187175.14]
    wire [31:0]     _GEN_6125; // @[ISA.scala 426:109:@187175.14]
    wire [31:0]     _GEN_6126; // @[ISA.scala 426:109:@187175.14]
    wire [31:0]     _GEN_6127; // @[ISA.scala 426:109:@187175.14]
    wire [31:0]     _GEN_6128; // @[ISA.scala 426:109:@187175.14]
    wire [31:0]     _GEN_6129; // @[ISA.scala 426:109:@187175.14]
    wire [63:0]     _GEN_6130; // @[ISA.scala 426:109:@187175.14]
    wire [63:0]     _GEN_6131; // @[ISA.scala 426:109:@187175.14]
    wire [31:0]     _GEN_6132; // @[ISA.scala 426:109:@187175.14]
    wire [31:0]     _GEN_6133; // @[ISA.scala 426:109:@187175.14]
    wire [31:0]     _GEN_6134; // @[ISA.scala 426:109:@187175.14]
    wire [31:0]     _GEN_6135; // @[ISA.scala 426:109:@187175.14]
    wire [63:0]     _GEN_6136; // @[ISA.scala 426:109:@187175.14]
    wire            _GEN_6137; // @[ISA.scala 426:109:@187175.14]
    wire            _GEN_6138; // @[ISA.scala 426:109:@187175.14]
    wire            _GEN_6139; // @[ISA.scala 426:109:@187175.14]
    wire [2:0]      _GEN_6140; // @[ISA.scala 425:101:@187003.12]
    wire [63:0]     _GEN_6141; // @[ISA.scala 425:101:@187003.12]
    wire [31:0]     _GEN_6142; // @[ISA.scala 425:101:@187003.12]
    wire [31:0]     _GEN_6143; // @[ISA.scala 425:101:@187003.12]
    wire [31:0]     _GEN_6144; // @[ISA.scala 425:101:@187003.12]
    wire [31:0]     _GEN_6145; // @[ISA.scala 425:101:@187003.12]
    wire [31:0]     _GEN_6146; // @[ISA.scala 425:101:@187003.12]
    wire [63:0]     _GEN_6147; // @[ISA.scala 425:101:@187003.12]
    wire [63:0]     _GEN_6148; // @[ISA.scala 425:101:@187003.12]
    wire [31:0]     _GEN_6149; // @[ISA.scala 425:101:@187003.12]
    wire [31:0]     _GEN_6150; // @[ISA.scala 425:101:@187003.12]
    wire [31:0]     _GEN_6151; // @[ISA.scala 425:101:@187003.12]
    wire [31:0]     _GEN_6152; // @[ISA.scala 425:101:@187003.12]
    wire [63:0]     _GEN_6153; // @[ISA.scala 425:101:@187003.12]
    wire            _GEN_6154; // @[ISA.scala 425:101:@187003.12]
    wire            _GEN_6155; // @[ISA.scala 425:101:@187003.12]
    wire            _GEN_6156; // @[ISA.scala 425:101:@187003.12]
    wire [2:0]      _GEN_6157; // @[ISA.scala 424:93:@186831.10]
    wire [63:0]     _GEN_6158; // @[ISA.scala 424:93:@186831.10]
    wire [31:0]     _GEN_6159; // @[ISA.scala 424:93:@186831.10]
    wire [31:0]     _GEN_6160; // @[ISA.scala 424:93:@186831.10]
    wire [31:0]     _GEN_6161; // @[ISA.scala 424:93:@186831.10]
    wire [31:0]     _GEN_6162; // @[ISA.scala 424:93:@186831.10]
    wire [31:0]     _GEN_6163; // @[ISA.scala 424:93:@186831.10]
    wire [63:0]     _GEN_6164; // @[ISA.scala 424:93:@186831.10]
    wire [63:0]     _GEN_6165; // @[ISA.scala 424:93:@186831.10]
    wire [31:0]     _GEN_6166; // @[ISA.scala 424:93:@186831.10]
    wire [31:0]     _GEN_6167; // @[ISA.scala 424:93:@186831.10]
    wire [31:0]     _GEN_6168; // @[ISA.scala 424:93:@186831.10]
    wire [31:0]     _GEN_6169; // @[ISA.scala 424:93:@186831.10]
    wire [63:0]     _GEN_6170; // @[ISA.scala 424:93:@186831.10]
    wire            _GEN_6171; // @[ISA.scala 424:93:@186831.10]
    wire            _GEN_6172; // @[ISA.scala 424:93:@186831.10]
    wire            _GEN_6173; // @[ISA.scala 424:93:@186831.10]
    wire [2:0]      _GEN_6174; // @[ISA.scala 423:85:@186659.8]
    wire [63:0]     _GEN_6175; // @[ISA.scala 423:85:@186659.8]
    wire [31:0]     _GEN_6176; // @[ISA.scala 423:85:@186659.8]
    wire [31:0]     _GEN_6177; // @[ISA.scala 423:85:@186659.8]
    wire [31:0]     _GEN_6178; // @[ISA.scala 423:85:@186659.8]
    wire [31:0]     _GEN_6179; // @[ISA.scala 423:85:@186659.8]
    wire [31:0]     _GEN_6180; // @[ISA.scala 423:85:@186659.8]
    wire [63:0]     _GEN_6181; // @[ISA.scala 423:85:@186659.8]
    wire [63:0]     _GEN_6182; // @[ISA.scala 423:85:@186659.8]
    wire [31:0]     _GEN_6183; // @[ISA.scala 423:85:@186659.8]
    wire [31:0]     _GEN_6184; // @[ISA.scala 423:85:@186659.8]
    wire [31:0]     _GEN_6185; // @[ISA.scala 423:85:@186659.8]
    wire [31:0]     _GEN_6186; // @[ISA.scala 423:85:@186659.8]
    wire [63:0]     _GEN_6187; // @[ISA.scala 423:85:@186659.8]
    wire            _GEN_6188; // @[ISA.scala 423:85:@186659.8]
    wire            _GEN_6189; // @[ISA.scala 423:85:@186659.8]
    wire            _GEN_6190; // @[ISA.scala 423:85:@186659.8]
    wire [2:0]      _GEN_6191; // @[ISA.scala 422:44:@186487.6]
    wire [63:0]     _GEN_6192; // @[ISA.scala 422:44:@186487.6]
    wire [31:0]     _GEN_6193; // @[ISA.scala 422:44:@186487.6]
    wire [31:0]     _GEN_6194; // @[ISA.scala 422:44:@186487.6]
    wire [31:0]     _GEN_6195; // @[ISA.scala 422:44:@186487.6]
    wire [31:0]     _GEN_6196; // @[ISA.scala 422:44:@186487.6]
    wire [31:0]     _GEN_6197; // @[ISA.scala 422:44:@186487.6]
    wire [63:0]     _GEN_6198; // @[ISA.scala 422:44:@186487.6]
    wire [63:0]     _GEN_6199; // @[ISA.scala 422:44:@186487.6]
    wire [31:0]     _GEN_6200; // @[ISA.scala 422:44:@186487.6]
    wire [31:0]     _GEN_6201; // @[ISA.scala 422:44:@186487.6]
    wire [31:0]     _GEN_6202; // @[ISA.scala 422:44:@186487.6]
    wire [31:0]     _GEN_6203; // @[ISA.scala 422:44:@186487.6]
    wire [63:0]     _GEN_6204; // @[ISA.scala 422:44:@186487.6]
    wire            _GEN_6205; // @[ISA.scala 422:44:@186487.6]
    wire            _GEN_6206; // @[ISA.scala 422:44:@186487.6]
    wire            _GEN_6207; // @[ISA.scala 422:44:@186487.6]
    wire [63:0]     _GEN_6209; // @[ISA.scala 87:28:@18.4]
    wire [63:0]     _GEN_6215; // @[ISA.scala 87:28:@18.4]
    wire [63:0]     _GEN_6216; // @[ISA.scala 87:28:@18.4]
    wire [63:0]     _GEN_6224; // @[ISA.scala 87:28:@18.4]
    assign _T_43 = state_r == 3'h0; // @[ISA.scala 105:30:@36.6]
    assign _GEN_0 = io_toMemoryPort_sync ? 3'h1 : state_r; // @[ISA.scala 106:52:@38.8]
    assign _GEN_8 = io_toMemoryPort_sync ? 1'h1 : fromMemoryPort_notify_r; // @[ISA.scala 106:52:@38.8]
    assign _GEN_9 = io_toMemoryPort_sync ? 1'h0 : toMemoryPort_notify_r; // @[ISA.scala 106:52:@38.8]
    assign _GEN_10 = io_toMemoryPort_sync ? 1'h0 : toRegsPort_notify_r; // @[ISA.scala 106:52:@38.8]
    assign _GEN_11 = _T_43 ? _GEN_0 : state_r; // @[ISA.scala 105:45:@37.6]
    assign _GEN_19 = _T_43 ? _GEN_8 : fromMemoryPort_notify_r; // @[ISA.scala 105:45:@37.6]
    assign _GEN_20 = _T_43 ? _GEN_9 : toMemoryPort_notify_r; // @[ISA.scala 105:45:@37.6]
    assign _GEN_21 = _T_43 ? _GEN_10 : toRegsPort_notify_r; // @[ISA.scala 105:45:@37.6]
    assign _T_47 = state_r == 3'h1; // @[ISA.scala 120:30:@52.6]
    assign _T_49 = 32'h4 + pcReg_signal_r; // @[ISA.scala 123:76:@56.10]
    assign _T_50 = 32'h4 + pcReg_signal_r; // @[ISA.scala 123:76:@57.10]
    assign _GEN_22 = io_fromMemoryPort_sync ? 3'h4 : _GEN_11; // @[ISA.scala 121:54:@54.8]
    assign _GEN_23 = io_fromMemoryPort_sync ? _T_50 : memoryAccess_signal_r_addrIn; // @[ISA.scala 121:54:@54.8]
    assign _GEN_24 = io_fromMemoryPort_sync ? 32'h0 : memoryAccess_signal_r_dataIn; // @[ISA.scala 121:54:@54.8]
    assign _GEN_25 = io_fromMemoryPort_sync ? 32'h1 : memoryAccess_signal_r_mask; // @[ISA.scala 121:54:@54.8]
    assign _GEN_26 = io_fromMemoryPort_sync ? 32'h1 : memoryAccess_signal_r_req; // @[ISA.scala 121:54:@54.8]
    assign _GEN_27 = io_fromMemoryPort_sync ? _T_50 : pcReg_signal_r; // @[ISA.scala 121:54:@54.8]
    assign _GEN_30 = io_fromMemoryPort_sync ? _T_50 : toMemoryPort_r_addrIn; // @[ISA.scala 121:54:@54.8]
    assign _GEN_31 = io_fromMemoryPort_sync ? 32'h0 : toMemoryPort_r_dataIn; // @[ISA.scala 121:54:@54.8]
    assign _GEN_32 = io_fromMemoryPort_sync ? 32'h1 : toMemoryPort_r_mask; // @[ISA.scala 121:54:@54.8]
    assign _GEN_33 = io_fromMemoryPort_sync ? 32'h1 : toMemoryPort_r_req; // @[ISA.scala 121:54:@54.8]
    assign _GEN_34 = io_fromMemoryPort_sync ? 1'h0 : _GEN_19; // @[ISA.scala 121:54:@54.8]
    assign _GEN_35 = io_fromMemoryPort_sync ? 1'h1 : _GEN_20; // @[ISA.scala 121:54:@54.8]
    assign _GEN_36 = io_fromMemoryPort_sync ? 1'h0 : _GEN_21; // @[ISA.scala 121:54:@54.8]
    assign _GEN_37 = _T_47 ? _GEN_22 : _GEN_11; // @[ISA.scala 120:45:@53.6]
    assign _GEN_38 = _T_47 ? _GEN_23 : memoryAccess_signal_r_addrIn; // @[ISA.scala 120:45:@53.6]
    assign _GEN_39 = _T_47 ? _GEN_24 : memoryAccess_signal_r_dataIn; // @[ISA.scala 120:45:@53.6]
    assign _GEN_40 = _T_47 ? _GEN_25 : memoryAccess_signal_r_mask; // @[ISA.scala 120:45:@53.6]
    assign _GEN_41 = _T_47 ? _GEN_26 : memoryAccess_signal_r_req; // @[ISA.scala 120:45:@53.6]
    assign _GEN_42 = _T_47 ? _GEN_27 : pcReg_signal_r; // @[ISA.scala 120:45:@53.6]
    assign _GEN_45 = _T_47 ? _GEN_30 : toMemoryPort_r_addrIn; // @[ISA.scala 120:45:@53.6]
    assign _GEN_46 = _T_47 ? _GEN_31 : toMemoryPort_r_dataIn; // @[ISA.scala 120:45:@53.6]
    assign _GEN_47 = _T_47 ? _GEN_32 : toMemoryPort_r_mask; // @[ISA.scala 120:45:@53.6]
    assign _GEN_48 = _T_47 ? _GEN_33 : toMemoryPort_r_req; // @[ISA.scala 120:45:@53.6]
    assign _GEN_49 = _T_47 ? _GEN_34 : _GEN_19; // @[ISA.scala 120:45:@53.6]
    assign _GEN_50 = _T_47 ? _GEN_35 : _GEN_20; // @[ISA.scala 120:45:@53.6]
    assign _GEN_51 = _T_47 ? _GEN_36 : _GEN_21; // @[ISA.scala 120:45:@53.6]
    assign _T_62 = state_r == 3'h2; // @[ISA.scala 139:30:@78.6]
    assign _GEN_52 = io_toMemoryPort_sync ? 3'h3 : _GEN_37; // @[ISA.scala 140:52:@80.8]
    assign _GEN_53 = io_toMemoryPort_sync ? memoryAccess_signal_r_addrIn : _GEN_38; // @[ISA.scala 140:52:@80.8]
    assign _GEN_54 = io_toMemoryPort_sync ? memoryAccess_signal_r_dataIn : _GEN_39; // @[ISA.scala 140:52:@80.8]
    assign _GEN_55 = io_toMemoryPort_sync ? memoryAccess_signal_r_mask : _GEN_40; // @[ISA.scala 140:52:@80.8]
    assign _GEN_56 = io_toMemoryPort_sync ? memoryAccess_signal_r_req : _GEN_41; // @[ISA.scala 140:52:@80.8]
    assign _GEN_57 = io_toMemoryPort_sync ? pcReg_signal_r : _GEN_42; // @[ISA.scala 140:52:@80.8]
    assign _GEN_60 = io_toMemoryPort_sync ? 1'h1 : _GEN_49; // @[ISA.scala 140:52:@80.8]
    assign _GEN_61 = io_toMemoryPort_sync ? 1'h0 : _GEN_50; // @[ISA.scala 140:52:@80.8]
    assign _GEN_62 = io_toMemoryPort_sync ? 1'h0 : _GEN_51; // @[ISA.scala 140:52:@80.8]
    assign _GEN_63 = _T_62 ? _GEN_52 : _GEN_37; // @[ISA.scala 139:46:@79.6]
    assign _GEN_64 = _T_62 ? _GEN_53 : _GEN_38; // @[ISA.scala 139:46:@79.6]
    assign _GEN_65 = _T_62 ? _GEN_54 : _GEN_39; // @[ISA.scala 139:46:@79.6]
    assign _GEN_66 = _T_62 ? _GEN_55 : _GEN_40; // @[ISA.scala 139:46:@79.6]
    assign _GEN_67 = _T_62 ? _GEN_56 : _GEN_41; // @[ISA.scala 139:46:@79.6]
    assign _GEN_68 = _T_62 ? _GEN_57 : _GEN_42; // @[ISA.scala 139:46:@79.6]
    assign _GEN_71 = _T_62 ? _GEN_60 : _GEN_49; // @[ISA.scala 139:46:@79.6]
    assign _GEN_72 = _T_62 ? _GEN_61 : _GEN_50; // @[ISA.scala 139:46:@79.6]
    assign _GEN_73 = _T_62 ? _GEN_62 : _GEN_51; // @[ISA.scala 139:46:@79.6]
    assign _T_66 = state_r == 3'h3; // @[ISA.scala 154:30:@94.6]
    assign _GEN_74 = io_fromMemoryPort_sync ? 3'h4 : _GEN_63; // @[ISA.scala 155:54:@96.8]
    assign _GEN_75 = io_fromMemoryPort_sync ? _T_50 : _GEN_64; // @[ISA.scala 155:54:@96.8]
    assign _GEN_76 = io_fromMemoryPort_sync ? 32'h0 : _GEN_65; // @[ISA.scala 155:54:@96.8]
    assign _GEN_77 = io_fromMemoryPort_sync ? 32'h1 : _GEN_66; // @[ISA.scala 155:54:@96.8]
    assign _GEN_78 = io_fromMemoryPort_sync ? 32'h1 : _GEN_67; // @[ISA.scala 155:54:@96.8]
    assign _GEN_79 = io_fromMemoryPort_sync ? _T_50 : _GEN_68; // @[ISA.scala 155:54:@96.8]
    assign _GEN_81 = io_fromMemoryPort_sync ? io_fromMemoryPort_loadedData : regfileWrite_signal_r_dstData; // @[ISA.scala 155:54:@96.8]
    assign _GEN_82 = io_fromMemoryPort_sync ? _T_50 : _GEN_45; // @[ISA.scala 155:54:@96.8]
    assign _GEN_83 = io_fromMemoryPort_sync ? 32'h0 : _GEN_46; // @[ISA.scala 155:54:@96.8]
    assign _GEN_84 = io_fromMemoryPort_sync ? 32'h1 : _GEN_47; // @[ISA.scala 155:54:@96.8]
    assign _GEN_85 = io_fromMemoryPort_sync ? 32'h1 : _GEN_48; // @[ISA.scala 155:54:@96.8]
    assign _GEN_86 = io_fromMemoryPort_sync ? regfileWrite_signal_r_dst : toRegsPort_r_dst; // @[ISA.scala 155:54:@96.8]
    assign _GEN_87 = io_fromMemoryPort_sync ? io_fromMemoryPort_loadedData : toRegsPort_r_dstData; // @[ISA.scala 155:54:@96.8]
    assign _GEN_88 = io_fromMemoryPort_sync ? 1'h0 : _GEN_71; // @[ISA.scala 155:54:@96.8]
    assign _GEN_89 = io_fromMemoryPort_sync ? 1'h1 : _GEN_72; // @[ISA.scala 155:54:@96.8]
    assign _GEN_90 = io_fromMemoryPort_sync ? 1'h1 : _GEN_73; // @[ISA.scala 155:54:@96.8]
    assign _GEN_91 = _T_66 ? _GEN_74 : _GEN_63; // @[ISA.scala 154:46:@95.6]
    assign _GEN_92 = _T_66 ? _GEN_75 : _GEN_64; // @[ISA.scala 154:46:@95.6]
    assign _GEN_93 = _T_66 ? _GEN_76 : _GEN_65; // @[ISA.scala 154:46:@95.6]
    assign _GEN_94 = _T_66 ? _GEN_77 : _GEN_66; // @[ISA.scala 154:46:@95.6]
    assign _GEN_95 = _T_66 ? _GEN_78 : _GEN_67; // @[ISA.scala 154:46:@95.6]
    assign _GEN_96 = _T_66 ? _GEN_79 : _GEN_68; // @[ISA.scala 154:46:@95.6]
    assign _GEN_98 = _T_66 ? _GEN_81 : regfileWrite_signal_r_dstData; // @[ISA.scala 154:46:@95.6]
    assign _GEN_99 = _T_66 ? _GEN_82 : _GEN_45; // @[ISA.scala 154:46:@95.6]
    assign _GEN_100 = _T_66 ? _GEN_83 : _GEN_46; // @[ISA.scala 154:46:@95.6]
    assign _GEN_101 = _T_66 ? _GEN_84 : _GEN_47; // @[ISA.scala 154:46:@95.6]
    assign _GEN_102 = _T_66 ? _GEN_85 : _GEN_48; // @[ISA.scala 154:46:@95.6]
    assign _GEN_103 = _T_66 ? _GEN_86 : toRegsPort_r_dst; // @[ISA.scala 154:46:@95.6]
    assign _GEN_104 = _T_66 ? _GEN_87 : toRegsPort_r_dstData; // @[ISA.scala 154:46:@95.6]
    assign _GEN_105 = _T_66 ? _GEN_88 : _GEN_71; // @[ISA.scala 154:46:@95.6]
    assign _GEN_106 = _T_66 ? _GEN_89 : _GEN_72; // @[ISA.scala 154:46:@95.6]
    assign _GEN_107 = _T_66 ? _GEN_90 : _GEN_73; // @[ISA.scala 154:46:@95.6]
    assign _T_81 = state_r == 3'h4; // @[ISA.scala 175:30:@122.6]
    assign _GEN_108 = io_toMemoryPort_sync ? 3'h5 : _GEN_91; // @[ISA.scala 176:52:@124.8]
    assign _GEN_109 = io_toMemoryPort_sync ? memoryAccess_signal_r_addrIn : _GEN_92; // @[ISA.scala 176:52:@124.8]
    assign _GEN_110 = io_toMemoryPort_sync ? memoryAccess_signal_r_dataIn : _GEN_93; // @[ISA.scala 176:52:@124.8]
    assign _GEN_111 = io_toMemoryPort_sync ? memoryAccess_signal_r_mask : _GEN_94; // @[ISA.scala 176:52:@124.8]
    assign _GEN_112 = io_toMemoryPort_sync ? memoryAccess_signal_r_req : _GEN_95; // @[ISA.scala 176:52:@124.8]
    assign _GEN_113 = io_toMemoryPort_sync ? pcReg_signal_r : _GEN_96; // @[ISA.scala 176:52:@124.8]
    assign _GEN_115 = io_toMemoryPort_sync ? regfileWrite_signal_r_dstData : _GEN_98; // @[ISA.scala 176:52:@124.8]
    assign _GEN_116 = io_toMemoryPort_sync ? 1'h1 : _GEN_105; // @[ISA.scala 176:52:@124.8]
    assign _GEN_117 = io_toMemoryPort_sync ? 1'h0 : _GEN_106; // @[ISA.scala 176:52:@124.8]
    assign _GEN_118 = io_toMemoryPort_sync ? 1'h0 : _GEN_107; // @[ISA.scala 176:52:@124.8]
    assign _GEN_119 = _T_81 ? _GEN_108 : _GEN_91; // @[ISA.scala 175:44:@123.6]
    assign _GEN_120 = _T_81 ? _GEN_109 : _GEN_92; // @[ISA.scala 175:44:@123.6]
    assign _GEN_121 = _T_81 ? _GEN_110 : _GEN_93; // @[ISA.scala 175:44:@123.6]
    assign _GEN_122 = _T_81 ? _GEN_111 : _GEN_94; // @[ISA.scala 175:44:@123.6]
    assign _GEN_123 = _T_81 ? _GEN_112 : _GEN_95; // @[ISA.scala 175:44:@123.6]
    assign _GEN_124 = _T_81 ? _GEN_113 : _GEN_96; // @[ISA.scala 175:44:@123.6]
    assign _GEN_126 = _T_81 ? _GEN_115 : _GEN_98; // @[ISA.scala 175:44:@123.6]
    assign _GEN_127 = _T_81 ? _GEN_116 : _GEN_105; // @[ISA.scala 175:44:@123.6]
    assign _GEN_128 = _T_81 ? _GEN_117 : _GEN_106; // @[ISA.scala 175:44:@123.6]
    assign _GEN_129 = _T_81 ? _GEN_118 : _GEN_107; // @[ISA.scala 175:44:@123.6]
    assign _T_85 = state_r == 3'h5; // @[ISA.scala 190:30:@138.6]
    assign _T_89 = io_fromMemoryPort_loadedData & 32'h7f; // @[ISA_functions.scala 208:38:@141.8]
    assign _T_91 = _T_89 == 32'h33; // @[ISA_functions.scala 208:53:@142.8]
    assign _T_106 = _T_91 == 1'h0; // @[ISA_functions.scala 211:28:@149.10]
    assign _T_110 = _T_89 == 32'h13; // @[ISA_functions.scala 211:108:@151.10]
    assign _T_111 = _T_106 & _T_110; // @[ISA_functions.scala 211:75:@152.10]
    assign _T_123 = _T_110 == 1'h0; // @[ISA_functions.scala 214:78:@162.12]
    assign _T_124 = _T_106 & _T_123; // @[ISA_functions.scala 214:75:@163.12]
    assign _T_128 = _T_89 == 32'h3; // @[ISA_functions.scala 214:158:@165.12]
    assign _T_129 = _T_124 & _T_128; // @[ISA_functions.scala 214:125:@166.12]
    assign _T_148 = _T_128 == 1'h0; // @[ISA_functions.scala 217:128:@180.14]
    assign _T_149 = _T_124 & _T_148; // @[ISA_functions.scala 217:125:@181.14]
    assign _T_153 = _T_89 == 32'h67; // @[ISA_functions.scala 217:207:@183.14]
    assign _T_154 = _T_149 & _T_153; // @[ISA_functions.scala 217:174:@184.14]
    assign _T_180 = _T_153 == 1'h0; // @[ISA_functions.scala 220:177:@202.16]
    assign _T_181 = _T_149 & _T_180; // @[ISA_functions.scala 220:174:@203.16]
    assign _T_185 = _T_89 == 32'h23; // @[ISA_functions.scala 220:258:@205.16]
    assign _T_186 = _T_181 & _T_185; // @[ISA_functions.scala 220:225:@206.16]
    assign _T_219 = _T_185 == 1'h0; // @[ISA_functions.scala 223:228:@228.18]
    assign _T_220 = _T_181 & _T_219; // @[ISA_functions.scala 223:225:@229.18]
    assign _T_224 = _T_89 == 32'h63; // @[ISA_functions.scala 223:308:@231.18]
    assign _T_225 = _T_220 & _T_224; // @[ISA_functions.scala 223:275:@232.18]
    assign _T_265 = _T_224 == 1'h0; // @[ISA_functions.scala 226:278:@258.20]
    assign _T_266 = _T_220 & _T_265; // @[ISA_functions.scala 226:275:@259.20]
    assign _T_270 = _T_89 == 32'h37; // @[ISA_functions.scala 226:359:@261.20]
    assign _T_274 = _T_89 == 32'h17; // @[ISA_functions.scala 226:408:@263.20]
    assign _T_275 = _T_270 | _T_274; // @[ISA_functions.scala 226:375:@264.20]
    assign _T_276 = _T_266 & _T_275; // @[ISA_functions.scala 226:325:@265.20]
    assign _T_328 = _T_275 == 1'h0; // @[ISA_functions.scala 229:328:@298.22]
    assign _T_329 = _T_266 & _T_328; // @[ISA_functions.scala 229:325:@299.22]
    assign _T_333 = _T_89 == 32'h6f; // @[ISA_functions.scala 229:459:@301.22]
    assign _T_334 = _T_329 & _T_333; // @[ISA_functions.scala 229:426:@302.22]
    assign _GEN_130 = _T_334 ? 32'h7 : 32'h8; // @[ISA_functions.scala 229:477:@303.22]
    assign _GEN_131 = _T_276 ? 32'h6 : _GEN_130; // @[ISA_functions.scala 226:426:@266.20]
    assign _GEN_132 = _T_225 ? 32'h5 : _GEN_131; // @[ISA_functions.scala 223:325:@233.18]
    assign _GEN_133 = _T_186 ? 32'h4 : _GEN_132; // @[ISA_functions.scala 220:275:@207.16]
    assign _GEN_134 = _T_154 ? 32'h3 : _GEN_133; // @[ISA_functions.scala 217:225:@185.14]
    assign _GEN_135 = _T_129 ? 32'h2 : _GEN_134; // @[ISA_functions.scala 214:174:@167.12]
    assign _GEN_136 = _T_111 ? 32'h1 : _GEN_135; // @[ISA_functions.scala 211:125:@153.10]
    assign _GEN_137 = _T_91 ? 32'h0 : _GEN_136; // @[ISA_functions.scala 208:70:@143.8]
    assign _T_335 = _GEN_137 == 32'h0; // @[ISA.scala 191:73:@309.8]
    assign _T_337 = _T_335 == 1'h0; // @[ISA.scala 191:30:@310.8]
    assign _T_578 = _GEN_137 == 32'h5; // @[ISA.scala 192:81:@481.10]
    assign _T_580 = _T_578 == 1'h0; // @[ISA.scala 192:38:@482.10]
    assign _T_821 = _GEN_137 == 32'h4; // @[ISA.scala 193:89:@653.12]
    assign _T_823 = _T_821 == 1'h0; // @[ISA.scala 193:46:@654.12]
    assign _T_1064 = _GEN_137 == 32'h6; // @[ISA.scala 194:97:@825.14]
    assign _T_1066 = _T_1064 == 1'h0; // @[ISA.scala 194:54:@826.14]
    assign _T_1307 = _GEN_137 == 32'h7; // @[ISA.scala 195:105:@997.16]
    assign _T_1309 = _T_1307 == 1'h0; // @[ISA.scala 195:62:@998.16]
    assign _T_1550 = _GEN_137 == 32'h1; // @[ISA.scala 196:113:@1169.18]
    assign _T_1552 = _T_1550 == 1'h0; // @[ISA.scala 196:70:@1170.18]
    assign _T_1793 = _GEN_137 == 32'h2; // @[ISA.scala 197:121:@1341.20]
    assign _T_1795 = _T_1793 == 1'h0; // @[ISA.scala 197:78:@1342.20]
    assign _T_2036 = _GEN_137 == 32'h3; // @[ISA.scala 198:129:@1513.22]
    assign _T_2038 = _T_2036 == 1'h0; // @[ISA.scala 198:86:@1514.22]
    assign _GEN_194 = io_fromMemoryPort_sync ? 3'h4 : _GEN_119; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_195 = io_fromMemoryPort_sync ? pcReg_signal_r : _GEN_120; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_196 = io_fromMemoryPort_sync ? 32'h0 : _GEN_121; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_197 = io_fromMemoryPort_sync ? 32'h1 : _GEN_122; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_198 = io_fromMemoryPort_sync ? 32'h1 : _GEN_123; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_199 = io_fromMemoryPort_sync ? pcReg_signal_r : _GEN_124; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_201 = io_fromMemoryPort_sync ? regfileWrite_signal_r_dstData : _GEN_126; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_202 = io_fromMemoryPort_sync ? pcReg_signal_r : _GEN_99; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_203 = io_fromMemoryPort_sync ? 32'h0 : _GEN_100; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_204 = io_fromMemoryPort_sync ? 32'h1 : _GEN_101; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_205 = io_fromMemoryPort_sync ? 32'h1 : _GEN_102; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_206 = io_fromMemoryPort_sync ? 1'h0 : _GEN_127; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_207 = io_fromMemoryPort_sync ? 1'h1 : _GEN_128; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_208 = io_fromMemoryPort_sync ? 1'h0 : _GEN_129; // @[ISA.scala 199:118:@1516.24]
    assign _GEN_209 = _T_2038 ? _GEN_194 : _GEN_119; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_210 = _T_2038 ? _GEN_195 : _GEN_120; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_211 = _T_2038 ? _GEN_196 : _GEN_121; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_212 = _T_2038 ? _GEN_197 : _GEN_122; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_213 = _T_2038 ? _GEN_198 : _GEN_123; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_214 = _T_2038 ? _GEN_199 : _GEN_124; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_216 = _T_2038 ? _GEN_201 : _GEN_126; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_217 = _T_2038 ? _GEN_202 : _GEN_99; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_218 = _T_2038 ? _GEN_203 : _GEN_100; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_219 = _T_2038 ? _GEN_204 : _GEN_101; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_220 = _T_2038 ? _GEN_205 : _GEN_102; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_221 = _T_2038 ? _GEN_206 : _GEN_127; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_222 = _T_2038 ? _GEN_207 : _GEN_128; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_223 = _T_2038 ? _GEN_208 : _GEN_129; // @[ISA.scala 198:143:@1515.22]
    assign _GEN_224 = _T_1795 ? _GEN_209 : _GEN_119; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_225 = _T_1795 ? _GEN_210 : _GEN_120; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_226 = _T_1795 ? _GEN_211 : _GEN_121; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_227 = _T_1795 ? _GEN_212 : _GEN_122; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_228 = _T_1795 ? _GEN_213 : _GEN_123; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_229 = _T_1795 ? _GEN_214 : _GEN_124; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_231 = _T_1795 ? _GEN_216 : _GEN_126; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_232 = _T_1795 ? _GEN_217 : _GEN_99; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_233 = _T_1795 ? _GEN_218 : _GEN_100; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_234 = _T_1795 ? _GEN_219 : _GEN_101; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_235 = _T_1795 ? _GEN_220 : _GEN_102; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_236 = _T_1795 ? _GEN_221 : _GEN_127; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_237 = _T_1795 ? _GEN_222 : _GEN_128; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_238 = _T_1795 ? _GEN_223 : _GEN_129; // @[ISA.scala 197:135:@1343.20]
    assign _GEN_239 = _T_1552 ? _GEN_224 : _GEN_119; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_240 = _T_1552 ? _GEN_225 : _GEN_120; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_241 = _T_1552 ? _GEN_226 : _GEN_121; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_242 = _T_1552 ? _GEN_227 : _GEN_122; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_243 = _T_1552 ? _GEN_228 : _GEN_123; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_244 = _T_1552 ? _GEN_229 : _GEN_124; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_246 = _T_1552 ? _GEN_231 : _GEN_126; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_247 = _T_1552 ? _GEN_232 : _GEN_99; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_248 = _T_1552 ? _GEN_233 : _GEN_100; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_249 = _T_1552 ? _GEN_234 : _GEN_101; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_250 = _T_1552 ? _GEN_235 : _GEN_102; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_251 = _T_1552 ? _GEN_236 : _GEN_127; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_252 = _T_1552 ? _GEN_237 : _GEN_128; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_253 = _T_1552 ? _GEN_238 : _GEN_129; // @[ISA.scala 196:127:@1171.18]
    assign _GEN_254 = _T_1309 ? _GEN_239 : _GEN_119; // @[ISA.scala 195:117:@999.16]
    assign _GEN_255 = _T_1309 ? _GEN_240 : _GEN_120; // @[ISA.scala 195:117:@999.16]
    assign _GEN_256 = _T_1309 ? _GEN_241 : _GEN_121; // @[ISA.scala 195:117:@999.16]
    assign _GEN_257 = _T_1309 ? _GEN_242 : _GEN_122; // @[ISA.scala 195:117:@999.16]
    assign _GEN_258 = _T_1309 ? _GEN_243 : _GEN_123; // @[ISA.scala 195:117:@999.16]
    assign _GEN_259 = _T_1309 ? _GEN_244 : _GEN_124; // @[ISA.scala 195:117:@999.16]
    assign _GEN_261 = _T_1309 ? _GEN_246 : _GEN_126; // @[ISA.scala 195:117:@999.16]
    assign _GEN_262 = _T_1309 ? _GEN_247 : _GEN_99; // @[ISA.scala 195:117:@999.16]
    assign _GEN_263 = _T_1309 ? _GEN_248 : _GEN_100; // @[ISA.scala 195:117:@999.16]
    assign _GEN_264 = _T_1309 ? _GEN_249 : _GEN_101; // @[ISA.scala 195:117:@999.16]
    assign _GEN_265 = _T_1309 ? _GEN_250 : _GEN_102; // @[ISA.scala 195:117:@999.16]
    assign _GEN_266 = _T_1309 ? _GEN_251 : _GEN_127; // @[ISA.scala 195:117:@999.16]
    assign _GEN_267 = _T_1309 ? _GEN_252 : _GEN_128; // @[ISA.scala 195:117:@999.16]
    assign _GEN_268 = _T_1309 ? _GEN_253 : _GEN_129; // @[ISA.scala 195:117:@999.16]
    assign _GEN_269 = _T_1066 ? _GEN_254 : _GEN_119; // @[ISA.scala 194:109:@827.14]
    assign _GEN_270 = _T_1066 ? _GEN_255 : _GEN_120; // @[ISA.scala 194:109:@827.14]
    assign _GEN_271 = _T_1066 ? _GEN_256 : _GEN_121; // @[ISA.scala 194:109:@827.14]
    assign _GEN_272 = _T_1066 ? _GEN_257 : _GEN_122; // @[ISA.scala 194:109:@827.14]
    assign _GEN_273 = _T_1066 ? _GEN_258 : _GEN_123; // @[ISA.scala 194:109:@827.14]
    assign _GEN_274 = _T_1066 ? _GEN_259 : _GEN_124; // @[ISA.scala 194:109:@827.14]
    assign _GEN_276 = _T_1066 ? _GEN_261 : _GEN_126; // @[ISA.scala 194:109:@827.14]
    assign _GEN_277 = _T_1066 ? _GEN_262 : _GEN_99; // @[ISA.scala 194:109:@827.14]
    assign _GEN_278 = _T_1066 ? _GEN_263 : _GEN_100; // @[ISA.scala 194:109:@827.14]
    assign _GEN_279 = _T_1066 ? _GEN_264 : _GEN_101; // @[ISA.scala 194:109:@827.14]
    assign _GEN_280 = _T_1066 ? _GEN_265 : _GEN_102; // @[ISA.scala 194:109:@827.14]
    assign _GEN_281 = _T_1066 ? _GEN_266 : _GEN_127; // @[ISA.scala 194:109:@827.14]
    assign _GEN_282 = _T_1066 ? _GEN_267 : _GEN_128; // @[ISA.scala 194:109:@827.14]
    assign _GEN_283 = _T_1066 ? _GEN_268 : _GEN_129; // @[ISA.scala 194:109:@827.14]
    assign _GEN_284 = _T_823 ? _GEN_269 : _GEN_119; // @[ISA.scala 193:101:@655.12]
    assign _GEN_285 = _T_823 ? _GEN_270 : _GEN_120; // @[ISA.scala 193:101:@655.12]
    assign _GEN_286 = _T_823 ? _GEN_271 : _GEN_121; // @[ISA.scala 193:101:@655.12]
    assign _GEN_287 = _T_823 ? _GEN_272 : _GEN_122; // @[ISA.scala 193:101:@655.12]
    assign _GEN_288 = _T_823 ? _GEN_273 : _GEN_123; // @[ISA.scala 193:101:@655.12]
    assign _GEN_289 = _T_823 ? _GEN_274 : _GEN_124; // @[ISA.scala 193:101:@655.12]
    assign _GEN_291 = _T_823 ? _GEN_276 : _GEN_126; // @[ISA.scala 193:101:@655.12]
    assign _GEN_292 = _T_823 ? _GEN_277 : _GEN_99; // @[ISA.scala 193:101:@655.12]
    assign _GEN_293 = _T_823 ? _GEN_278 : _GEN_100; // @[ISA.scala 193:101:@655.12]
    assign _GEN_294 = _T_823 ? _GEN_279 : _GEN_101; // @[ISA.scala 193:101:@655.12]
    assign _GEN_295 = _T_823 ? _GEN_280 : _GEN_102; // @[ISA.scala 193:101:@655.12]
    assign _GEN_296 = _T_823 ? _GEN_281 : _GEN_127; // @[ISA.scala 193:101:@655.12]
    assign _GEN_297 = _T_823 ? _GEN_282 : _GEN_128; // @[ISA.scala 193:101:@655.12]
    assign _GEN_298 = _T_823 ? _GEN_283 : _GEN_129; // @[ISA.scala 193:101:@655.12]
    assign _GEN_299 = _T_580 ? _GEN_284 : _GEN_119; // @[ISA.scala 192:93:@483.10]
    assign _GEN_300 = _T_580 ? _GEN_285 : _GEN_120; // @[ISA.scala 192:93:@483.10]
    assign _GEN_301 = _T_580 ? _GEN_286 : _GEN_121; // @[ISA.scala 192:93:@483.10]
    assign _GEN_302 = _T_580 ? _GEN_287 : _GEN_122; // @[ISA.scala 192:93:@483.10]
    assign _GEN_303 = _T_580 ? _GEN_288 : _GEN_123; // @[ISA.scala 192:93:@483.10]
    assign _GEN_304 = _T_580 ? _GEN_289 : _GEN_124; // @[ISA.scala 192:93:@483.10]
    assign _GEN_306 = _T_580 ? _GEN_291 : _GEN_126; // @[ISA.scala 192:93:@483.10]
    assign _GEN_307 = _T_580 ? _GEN_292 : _GEN_99; // @[ISA.scala 192:93:@483.10]
    assign _GEN_308 = _T_580 ? _GEN_293 : _GEN_100; // @[ISA.scala 192:93:@483.10]
    assign _GEN_309 = _T_580 ? _GEN_294 : _GEN_101; // @[ISA.scala 192:93:@483.10]
    assign _GEN_310 = _T_580 ? _GEN_295 : _GEN_102; // @[ISA.scala 192:93:@483.10]
    assign _GEN_311 = _T_580 ? _GEN_296 : _GEN_127; // @[ISA.scala 192:93:@483.10]
    assign _GEN_312 = _T_580 ? _GEN_297 : _GEN_128; // @[ISA.scala 192:93:@483.10]
    assign _GEN_313 = _T_580 ? _GEN_298 : _GEN_129; // @[ISA.scala 192:93:@483.10]
    assign _GEN_314 = _T_337 ? _GEN_299 : _GEN_119; // @[ISA.scala 191:85:@311.8]
    assign _GEN_315 = _T_337 ? _GEN_300 : _GEN_120; // @[ISA.scala 191:85:@311.8]
    assign _GEN_316 = _T_337 ? _GEN_301 : _GEN_121; // @[ISA.scala 191:85:@311.8]
    assign _GEN_317 = _T_337 ? _GEN_302 : _GEN_122; // @[ISA.scala 191:85:@311.8]
    assign _GEN_318 = _T_337 ? _GEN_303 : _GEN_123; // @[ISA.scala 191:85:@311.8]
    assign _GEN_319 = _T_337 ? _GEN_304 : _GEN_124; // @[ISA.scala 191:85:@311.8]
    assign _GEN_321 = _T_337 ? _GEN_306 : _GEN_126; // @[ISA.scala 191:85:@311.8]
    assign _GEN_322 = _T_337 ? _GEN_307 : _GEN_99; // @[ISA.scala 191:85:@311.8]
    assign _GEN_323 = _T_337 ? _GEN_308 : _GEN_100; // @[ISA.scala 191:85:@311.8]
    assign _GEN_324 = _T_337 ? _GEN_309 : _GEN_101; // @[ISA.scala 191:85:@311.8]
    assign _GEN_325 = _T_337 ? _GEN_310 : _GEN_102; // @[ISA.scala 191:85:@311.8]
    assign _GEN_326 = _T_337 ? _GEN_311 : _GEN_127; // @[ISA.scala 191:85:@311.8]
    assign _GEN_327 = _T_337 ? _GEN_312 : _GEN_128; // @[ISA.scala 191:85:@311.8]
    assign _GEN_328 = _T_337 ? _GEN_313 : _GEN_129; // @[ISA.scala 191:85:@311.8]
    assign _GEN_329 = _T_85 ? _GEN_314 : _GEN_119; // @[ISA.scala 190:44:@139.6]
    assign _GEN_330 = _T_85 ? _GEN_315 : _GEN_120; // @[ISA.scala 190:44:@139.6]
    assign _GEN_331 = _T_85 ? _GEN_316 : _GEN_121; // @[ISA.scala 190:44:@139.6]
    assign _GEN_332 = _T_85 ? _GEN_317 : _GEN_122; // @[ISA.scala 190:44:@139.6]
    assign _GEN_333 = _T_85 ? _GEN_318 : _GEN_123; // @[ISA.scala 190:44:@139.6]
    assign _GEN_334 = _T_85 ? _GEN_319 : _GEN_124; // @[ISA.scala 190:44:@139.6]
    assign _GEN_336 = _T_85 ? _GEN_321 : _GEN_126; // @[ISA.scala 190:44:@139.6]
    assign _GEN_337 = _T_85 ? _GEN_322 : _GEN_99; // @[ISA.scala 190:44:@139.6]
    assign _GEN_338 = _T_85 ? _GEN_323 : _GEN_100; // @[ISA.scala 190:44:@139.6]
    assign _GEN_339 = _T_85 ? _GEN_324 : _GEN_101; // @[ISA.scala 190:44:@139.6]
    assign _GEN_340 = _T_85 ? _GEN_325 : _GEN_102; // @[ISA.scala 190:44:@139.6]
    assign _GEN_341 = _T_85 ? _GEN_326 : _GEN_127; // @[ISA.scala 190:44:@139.6]
    assign _GEN_342 = _T_85 ? _GEN_327 : _GEN_128; // @[ISA.scala 190:44:@139.6]
    assign _GEN_343 = _T_85 ? _GEN_328 : _GEN_129; // @[ISA.scala 190:44:@139.6]
    assign _T_2303 = _T_91 | _T_110; // @[ISA_functions.scala 452:75:@1731.12]
    assign _T_2308 = _T_2303 | _T_128; // @[ISA_functions.scala 452:125:@1734.12]
    assign _T_2313 = _T_2308 | _T_153; // @[ISA_functions.scala 452:174:@1737.12]
    assign _T_2318 = _T_2313 | _T_270; // @[ISA_functions.scala 452:225:@1740.12]
    assign _T_2323 = _T_2318 | _T_274; // @[ISA_functions.scala 452:275:@1743.12]
    assign _T_2328 = _T_2323 | _T_333; // @[ISA_functions.scala 452:325:@1746.12]
    assign _T_2330 = io_fromMemoryPort_loadedData >> 32'h7; // @[ISA_functions.scala 453:48:@1748.14]
    assign _T_2333 = _T_2330 & 32'h1f; // @[ISA_functions.scala 453:69:@1750.14]
    assign _GEN_352 = _T_2328 ? _T_2333 : 32'h0; // @[ISA_functions.scala 452:377:@1747.12]
    assign _T_2342 = io_fromMemoryPort_loadedData >> 32'hc; // @[ISA_functions.scala 286:88:@1760.12]
    assign _T_2345 = _T_2342 & 32'h7; // @[ISA_functions.scala 286:110:@1762.12]
    assign _T_2347 = _T_2345 == 32'h0; // @[ISA_functions.scala 286:123:@1763.12]
    assign _T_2348 = _T_91 & _T_2347; // @[ISA_functions.scala 286:69:@1764.12]
    assign _T_2350 = io_fromMemoryPort_loadedData >> 32'h19; // @[ISA_functions.scala 286:157:@1765.12]
    assign _T_2353 = _T_2350 & 32'h7f; // @[ISA_functions.scala 286:179:@1767.12]
    assign _T_2355 = _T_2353 == 32'h0; // @[ISA_functions.scala 286:194:@1768.12]
    assign _T_2356 = _T_2348 & _T_2355; // @[ISA_functions.scala 286:138:@1769.12]
    assign _T_2415 = _T_2355 == 1'h0; // @[ISA_functions.scala 289:146:@1785.14]
    assign _T_2416 = _T_2348 & _T_2415; // @[ISA_functions.scala 289:143:@1786.14]
    assign _T_2423 = _T_2353 == 32'h20; // @[ISA_functions.scala 289:271:@1790.14]
    assign _T_2424 = _T_2416 & _T_2423; // @[ISA_functions.scala 289:215:@1791.14]
    assign _T_2455 = _T_2423 == 1'h0; // @[ISA_functions.scala 292:218:@1813.16]
    assign _T_2456 = _T_2416 & _T_2455; // @[ISA_functions.scala 292:215:@1814.16]
    assign _T_2469 = _T_2347 == 1'h0; // @[ISA_functions.scala 295:77:@1825.18]
    assign _T_2470 = _T_91 & _T_2469; // @[ISA_functions.scala 295:74:@1826.18]
    assign _T_2477 = _T_2345 == 32'h1; // @[ISA_functions.scala 295:198:@1830.18]
    assign _T_2478 = _T_2470 & _T_2477; // @[ISA_functions.scala 295:144:@1831.18]
    assign _T_2501 = _T_2477 == 1'h0; // @[ISA_functions.scala 298:147:@1848.20]
    assign _T_2502 = _T_2470 & _T_2501; // @[ISA_functions.scala 298:144:@1849.20]
    assign _T_2509 = _T_2345 == 32'h2; // @[ISA_functions.scala 298:268:@1853.20]
    assign _T_2510 = _T_2502 & _T_2509; // @[ISA_functions.scala 298:214:@1854.20]
    assign _T_2543 = _T_2509 == 1'h0; // @[ISA_functions.scala 301:217:@1877.22]
    assign _T_2544 = _T_2502 & _T_2543; // @[ISA_functions.scala 301:214:@1878.22]
    assign _T_2551 = _T_2345 == 32'h3; // @[ISA_functions.scala 301:338:@1882.22]
    assign _T_2552 = _T_2544 & _T_2551; // @[ISA_functions.scala 301:284:@1883.22]
    assign _T_2595 = _T_2551 == 1'h0; // @[ISA_functions.scala 304:287:@1912.24]
    assign _T_2596 = _T_2544 & _T_2595; // @[ISA_functions.scala 304:284:@1913.24]
    assign _T_2603 = _T_2345 == 32'h4; // @[ISA_functions.scala 304:408:@1917.24]
    assign _T_2604 = _T_2596 & _T_2603; // @[ISA_functions.scala 304:354:@1918.24]
    assign _T_2657 = _T_2603 == 1'h0; // @[ISA_functions.scala 307:357:@1953.26]
    assign _T_2658 = _T_2596 & _T_2657; // @[ISA_functions.scala 307:354:@1954.26]
    assign _T_2665 = _T_2345 == 32'h5; // @[ISA_functions.scala 307:478:@1958.26]
    assign _T_2666 = _T_2658 & _T_2665; // @[ISA_functions.scala 307:424:@1959.26]
    assign _T_2674 = _T_2666 & _T_2355; // @[ISA_functions.scala 307:493:@1964.26]
    assign _T_2746 = _T_2666 & _T_2415; // @[ISA_functions.scala 310:493:@2011.28]
    assign _T_2754 = _T_2746 & _T_2423; // @[ISA_functions.scala 310:565:@2016.28]
    assign _T_2836 = _T_2746 & _T_2455; // @[ISA_functions.scala 313:565:@2069.30]
    assign _T_2899 = _T_2665 == 1'h0; // @[ISA_functions.scala 316:427:@2110.32]
    assign _T_2900 = _T_2658 & _T_2899; // @[ISA_functions.scala 316:424:@2111.32]
    assign _T_2907 = _T_2345 == 32'h6; // @[ISA_functions.scala 316:548:@2115.32]
    assign _T_2908 = _T_2900 & _T_2907; // @[ISA_functions.scala 316:494:@2116.32]
    assign _T_2981 = _T_2907 == 1'h0; // @[ISA_functions.scala 319:497:@2163.34]
    assign _T_2982 = _T_2900 & _T_2981; // @[ISA_functions.scala 319:494:@2164.34]
    assign _T_2989 = _T_2345 == 32'h7; // @[ISA_functions.scala 319:618:@2168.34]
    assign _T_2990 = _T_2982 & _T_2989; // @[ISA_functions.scala 319:564:@2169.34]
    assign _T_3073 = _T_2989 == 1'h0; // @[ISA_functions.scala 322:567:@2222.36]
    assign _T_3074 = _T_2982 & _T_3073; // @[ISA_functions.scala 322:564:@2223.36]
    assign _T_3093 = _T_111 & _T_2347; // @[ISA_functions.scala 325:124:@2238.38]
    assign _T_3114 = _T_111 & _T_2469; // @[ISA_functions.scala 328:124:@2254.40]
    assign _T_3122 = _T_3114 & _T_2477; // @[ISA_functions.scala 328:194:@2259.40]
    assign _T_3153 = _T_3114 & _T_2501; // @[ISA_functions.scala 331:194:@2281.42]
    assign _T_3161 = _T_3153 & _T_2509; // @[ISA_functions.scala 331:264:@2286.42]
    assign _T_3202 = _T_3153 & _T_2543; // @[ISA_functions.scala 334:264:@2314.44]
    assign _T_3210 = _T_3202 & _T_2551; // @[ISA_functions.scala 334:334:@2319.44]
    assign _T_3261 = _T_3202 & _T_2595; // @[ISA_functions.scala 337:334:@2353.46]
    assign _T_3269 = _T_3261 & _T_2603; // @[ISA_functions.scala 337:404:@2358.46]
    assign _T_3330 = _T_3261 & _T_2657; // @[ISA_functions.scala 340:404:@2398.48]
    assign _T_3338 = _T_3330 & _T_2665; // @[ISA_functions.scala 340:474:@2403.48]
    assign _T_3346 = _T_3338 & _T_2355; // @[ISA_functions.scala 340:543:@2408.48]
    assign _T_3425 = _T_3338 & _T_2415; // @[ISA_functions.scala 343:543:@2459.50]
    assign _T_3433 = _T_3425 & _T_2423; // @[ISA_functions.scala 343:615:@2464.50]
    assign _T_3522 = _T_3425 & _T_2455; // @[ISA_functions.scala 346:615:@2521.52]
    assign _T_3593 = _T_3330 & _T_2899; // @[ISA_functions.scala 349:474:@2567.54]
    assign _T_3601 = _T_3593 & _T_2907; // @[ISA_functions.scala 349:544:@2572.54]
    assign _T_3682 = _T_3593 & _T_2981; // @[ISA_functions.scala 352:544:@2624.56]
    assign _T_3690 = _T_3682 & _T_2989; // @[ISA_functions.scala 352:614:@2629.56]
    assign _T_3781 = _T_3682 & _T_3073; // @[ISA_functions.scala 355:614:@2687.58]
    assign _T_3807 = _T_129 & _T_2347; // @[ISA_functions.scala 358:173:@2706.60]
    assign _T_3835 = _T_129 & _T_2469; // @[ISA_functions.scala 361:173:@2726.62]
    assign _T_3843 = _T_3835 & _T_2477; // @[ISA_functions.scala 361:243:@2731.62]
    assign _T_3881 = _T_3835 & _T_2501; // @[ISA_functions.scala 364:243:@2757.64]
    assign _T_3889 = _T_3881 & _T_2509; // @[ISA_functions.scala 364:313:@2762.64]
    assign _T_3937 = _T_3881 & _T_2543; // @[ISA_functions.scala 367:313:@2794.66]
    assign _T_3945 = _T_3937 & _T_2603; // @[ISA_functions.scala 367:383:@2799.66]
    assign _T_4003 = _T_3937 & _T_2657; // @[ISA_functions.scala 370:383:@2837.68]
    assign _T_4011 = _T_4003 & _T_2665; // @[ISA_functions.scala 370:453:@2842.68]
    assign _T_4079 = _T_4003 & _T_2899; // @[ISA_functions.scala 373:453:@2886.70]
    assign _T_4144 = _T_186 & _T_2347; // @[ISA_functions.scala 379:274:@2931.74]
    assign _T_4186 = _T_186 & _T_2469; // @[ISA_functions.scala 382:274:@2959.76]
    assign _T_4194 = _T_4186 & _T_2477; // @[ISA_functions.scala 382:344:@2964.76]
    assign _T_4246 = _T_4186 & _T_2501; // @[ISA_functions.scala 385:344:@2998.78]
    assign _T_4254 = _T_4246 & _T_2509; // @[ISA_functions.scala 385:414:@3003.78]
    assign _T_4316 = _T_4246 & _T_2543; // @[ISA_functions.scala 388:414:@3043.80]
    assign _T_4363 = _T_225 & _T_2347; // @[ISA_functions.scala 391:324:@3074.82]
    assign _T_4412 = _T_225 & _T_2469; // @[ISA_functions.scala 394:324:@3106.84]
    assign _T_4420 = _T_4412 & _T_2477; // @[ISA_functions.scala 394:394:@3111.84]
    assign _T_4479 = _T_4412 & _T_2501; // @[ISA_functions.scala 397:394:@3149.86]
    assign _T_4487 = _T_4479 & _T_2603; // @[ISA_functions.scala 397:464:@3154.86]
    assign _T_4556 = _T_4479 & _T_2657; // @[ISA_functions.scala 400:464:@3198.88]
    assign _T_4564 = _T_4556 & _T_2665; // @[ISA_functions.scala 400:534:@3203.88]
    assign _T_4643 = _T_4556 & _T_2899; // @[ISA_functions.scala 403:534:@3253.90]
    assign _T_4651 = _T_4643 & _T_2907; // @[ISA_functions.scala 403:604:@3258.90]
    assign _T_4740 = _T_4643 & _T_2981; // @[ISA_functions.scala 406:604:@3314.92]
    assign _T_4748 = _T_4740 & _T_2989; // @[ISA_functions.scala 406:674:@3319.92]
    assign _T_4847 = _T_4740 & _T_3073; // @[ISA_functions.scala 409:674:@3381.94]
    assign _T_4893 = _T_266 & _T_270; // @[ISA_functions.scala 412:325:@3411.96]
    assign _T_4940 = _T_270 == 1'h0; // @[ISA_functions.scala 415:328:@3441.98]
    assign _T_4941 = _T_266 & _T_4940; // @[ISA_functions.scala 415:325:@3442.98]
    assign _T_4946 = _T_4941 & _T_274; // @[ISA_functions.scala 415:375:@3445.98]
    assign _T_5000 = _T_274 == 1'h0; // @[ISA_functions.scala 418:378:@3479.100]
    assign _T_5001 = _T_4941 & _T_5000; // @[ISA_functions.scala 418:375:@3480.100]
    assign _T_5006 = _T_5001 & _T_333; // @[ISA_functions.scala 418:425:@3483.100]
    assign _GEN_353 = _T_5006 ? 32'h25 : 32'h0; // @[ISA_functions.scala 418:476:@3484.100]
    assign _GEN_354 = _T_4946 ? 32'h24 : _GEN_353; // @[ISA_functions.scala 415:425:@3446.98]
    assign _GEN_355 = _T_4893 ? 32'h23 : _GEN_354; // @[ISA_functions.scala 412:375:@3412.96]
    assign _GEN_356 = _T_4847 ? 32'h0 : _GEN_355; // @[ISA_functions.scala 409:745:@3382.94]
    assign _GEN_357 = _T_4748 ? 32'h22 : _GEN_356; // @[ISA_functions.scala 406:744:@3320.92]
    assign _GEN_358 = _T_4651 ? 32'h21 : _GEN_357; // @[ISA_functions.scala 403:674:@3259.90]
    assign _GEN_359 = _T_4564 ? 32'h20 : _GEN_358; // @[ISA_functions.scala 400:604:@3204.88]
    assign _GEN_360 = _T_4487 ? 32'h1f : _GEN_359; // @[ISA_functions.scala 397:534:@3155.86]
    assign _GEN_361 = _T_4420 ? 32'h1e : _GEN_360; // @[ISA_functions.scala 394:464:@3112.84]
    assign _GEN_362 = _T_4363 ? 32'h1d : _GEN_361; // @[ISA_functions.scala 391:394:@3075.82]
    assign _GEN_363 = _T_4316 ? 32'h0 : _GEN_362; // @[ISA_functions.scala 388:485:@3044.80]
    assign _GEN_364 = _T_4254 ? 32'h1c : _GEN_363; // @[ISA_functions.scala 385:484:@3004.78]
    assign _GEN_365 = _T_4194 ? 32'h1b : _GEN_364; // @[ISA_functions.scala 382:414:@2965.76]
    assign _GEN_366 = _T_4144 ? 32'h1a : _GEN_365; // @[ISA_functions.scala 379:344:@2932.74]
    assign _GEN_367 = _T_154 ? 32'h19 : _GEN_366; // @[ISA_functions.scala 376:225:@2905.72]
    assign _GEN_368 = _T_4079 ? 32'h0 : _GEN_367; // @[ISA_functions.scala 373:524:@2887.70]
    assign _GEN_369 = _T_4011 ? 32'h18 : _GEN_368; // @[ISA_functions.scala 370:523:@2843.68]
    assign _GEN_370 = _T_3945 ? 32'h17 : _GEN_369; // @[ISA_functions.scala 367:453:@2800.66]
    assign _GEN_371 = _T_3889 ? 32'h16 : _GEN_370; // @[ISA_functions.scala 364:383:@2763.64]
    assign _GEN_372 = _T_3843 ? 32'h15 : _GEN_371; // @[ISA_functions.scala 361:313:@2732.62]
    assign _GEN_373 = _T_3807 ? 32'h14 : _GEN_372; // @[ISA_functions.scala 358:243:@2707.60]
    assign _GEN_374 = _T_3781 ? 32'h0 : _GEN_373; // @[ISA_functions.scala 355:685:@2688.58]
    assign _GEN_375 = _T_3690 ? 32'h13 : _GEN_374; // @[ISA_functions.scala 352:684:@2630.56]
    assign _GEN_376 = _T_3601 ? 32'h12 : _GEN_375; // @[ISA_functions.scala 349:614:@2573.54]
    assign _GEN_377 = _T_3522 ? 32'h0 : _GEN_376; // @[ISA_functions.scala 346:689:@2522.52]
    assign _GEN_378 = _T_3433 ? 32'h11 : _GEN_377; // @[ISA_functions.scala 343:688:@2465.50]
    assign _GEN_379 = _T_3346 ? 32'h10 : _GEN_378; // @[ISA_functions.scala 340:615:@2409.48]
    assign _GEN_380 = _T_3269 ? 32'hf : _GEN_379; // @[ISA_functions.scala 337:474:@2359.46]
    assign _GEN_381 = _T_3210 ? 32'he : _GEN_380; // @[ISA_functions.scala 334:404:@2320.44]
    assign _GEN_382 = _T_3161 ? 32'hd : _GEN_381; // @[ISA_functions.scala 331:334:@2287.42]
    assign _GEN_383 = _T_3122 ? 32'hc : _GEN_382; // @[ISA_functions.scala 328:264:@2260.40]
    assign _GEN_384 = _T_3093 ? 32'hb : _GEN_383; // @[ISA_functions.scala 325:194:@2239.38]
    assign _GEN_385 = _T_3074 ? 32'h0 : _GEN_384; // @[ISA_functions.scala 322:635:@2224.36]
    assign _GEN_386 = _T_2990 ? 32'ha : _GEN_385; // @[ISA_functions.scala 319:634:@2170.34]
    assign _GEN_387 = _T_2908 ? 32'h9 : _GEN_386; // @[ISA_functions.scala 316:564:@2117.32]
    assign _GEN_388 = _T_2836 ? 32'h0 : _GEN_387; // @[ISA_functions.scala 313:639:@2070.30]
    assign _GEN_389 = _T_2754 ? 32'h8 : _GEN_388; // @[ISA_functions.scala 310:638:@2017.28]
    assign _GEN_390 = _T_2674 ? 32'h7 : _GEN_389; // @[ISA_functions.scala 307:565:@1965.26]
    assign _GEN_391 = _T_2604 ? 32'h6 : _GEN_390; // @[ISA_functions.scala 304:424:@1919.24]
    assign _GEN_392 = _T_2552 ? 32'h5 : _GEN_391; // @[ISA_functions.scala 301:354:@1884.22]
    assign _GEN_393 = _T_2510 ? 32'h4 : _GEN_392; // @[ISA_functions.scala 298:284:@1855.20]
    assign _GEN_394 = _T_2478 ? 32'h3 : _GEN_393; // @[ISA_functions.scala 295:214:@1832.18]
    assign _GEN_395 = _T_2456 ? 32'h0 : _GEN_394; // @[ISA_functions.scala 292:289:@1815.16]
    assign _GEN_396 = _T_2424 ? 32'h2 : _GEN_395; // @[ISA_functions.scala 289:288:@1792.14]
    assign _GEN_397 = _T_2356 ? 32'h1 : _GEN_396; // @[ISA_functions.scala 286:210:@1770.12]
    assign _T_5009 = _GEN_397 == 32'h1; // @[ISA_functions.scala 117:40:@3491.12]
    assign _T_5010 = _GEN_397 == 32'hb; // @[ISA_functions.scala 117:65:@3492.12]
    assign _T_5011 = _T_5009 | _T_5010; // @[ISA_functions.scala 117:55:@3493.12]
    assign _T_5012 = _GEN_397 == 32'h14; // @[ISA_functions.scala 117:92:@3494.12]
    assign _T_5013 = _T_5011 | _T_5012; // @[ISA_functions.scala 117:82:@3495.12]
    assign _T_5014 = _GEN_397 == 32'h15; // @[ISA_functions.scala 117:117:@3496.12]
    assign _T_5015 = _T_5013 | _T_5014; // @[ISA_functions.scala 117:107:@3497.12]
    assign _T_5016 = _GEN_397 == 32'h16; // @[ISA_functions.scala 117:142:@3498.12]
    assign _T_5017 = _T_5015 | _T_5016; // @[ISA_functions.scala 117:132:@3499.12]
    assign _T_5018 = _GEN_397 == 32'h17; // @[ISA_functions.scala 117:167:@3500.12]
    assign _T_5019 = _T_5017 | _T_5018; // @[ISA_functions.scala 117:157:@3501.12]
    assign _T_5020 = _GEN_397 == 32'h18; // @[ISA_functions.scala 117:193:@3502.12]
    assign _T_5021 = _T_5019 | _T_5020; // @[ISA_functions.scala 117:183:@3503.12]
    assign _T_5022 = _GEN_397 == 32'h1a; // @[ISA_functions.scala 117:219:@3504.12]
    assign _T_5023 = _T_5021 | _T_5022; // @[ISA_functions.scala 117:209:@3505.12]
    assign _T_5024 = _GEN_397 == 32'h1b; // @[ISA_functions.scala 117:244:@3506.12]
    assign _T_5025 = _T_5023 | _T_5024; // @[ISA_functions.scala 117:234:@3507.12]
    assign _T_5026 = _GEN_397 == 32'h1c; // @[ISA_functions.scala 117:269:@3508.12]
    assign _T_5027 = _T_5025 | _T_5026; // @[ISA_functions.scala 117:259:@3509.12]
    assign _T_5028 = _GEN_397 == 32'h24; // @[ISA_functions.scala 117:294:@3510.12]
    assign _T_5029 = _T_5027 | _T_5028; // @[ISA_functions.scala 117:284:@3511.12]
    assign _T_5064 = _T_5029 == 1'h0; // @[ISA_functions.scala 120:28:@3537.14]
    assign _T_5065 = _GEN_397 == 32'h2; // @[ISA_functions.scala 120:330:@3538.14]
    assign _T_5066 = _GEN_397 == 32'h1d; // @[ISA_functions.scala 120:355:@3539.14]
    assign _T_5067 = _T_5065 | _T_5066; // @[ISA_functions.scala 120:345:@3540.14]
    assign _T_5068 = _GEN_397 == 32'h1e; // @[ISA_functions.scala 120:381:@3541.14]
    assign _T_5069 = _T_5067 | _T_5068; // @[ISA_functions.scala 120:371:@3542.14]
    assign _T_5070 = _T_5064 & _T_5069; // @[ISA_functions.scala 120:318:@3543.14]
    assign _T_5100 = _T_5069 == 1'h0; // @[ISA_functions.scala 123:321:@3575.16]
    assign _T_5101 = _T_5064 & _T_5100; // @[ISA_functions.scala 123:318:@3576.16]
    assign _T_5102 = _GEN_397 == 32'h3; // @[ISA_functions.scala 123:409:@3577.16]
    assign _T_5103 = _GEN_397 == 32'hc; // @[ISA_functions.scala 123:434:@3578.16]
    assign _T_5104 = _T_5102 | _T_5103; // @[ISA_functions.scala 123:424:@3579.16]
    assign _T_5105 = _T_5101 & _T_5104; // @[ISA_functions.scala 123:398:@3580.16]
    assign _T_5141 = _T_5104 == 1'h0; // @[ISA_functions.scala 126:401:@3617.18]
    assign _T_5142 = _T_5101 & _T_5141; // @[ISA_functions.scala 126:398:@3618.18]
    assign _T_5143 = _GEN_397 == 32'h4; // @[ISA_functions.scala 126:465:@3619.18]
    assign _T_5144 = _GEN_397 == 32'hd; // @[ISA_functions.scala 126:490:@3620.18]
    assign _T_5145 = _T_5143 | _T_5144; // @[ISA_functions.scala 126:480:@3621.18]
    assign _T_5146 = _GEN_397 == 32'h1f; // @[ISA_functions.scala 126:517:@3622.18]
    assign _T_5147 = _T_5145 | _T_5146; // @[ISA_functions.scala 126:507:@3623.18]
    assign _T_5148 = _GEN_397 == 32'h20; // @[ISA_functions.scala 126:543:@3624.18]
    assign _T_5149 = _T_5147 | _T_5148; // @[ISA_functions.scala 126:533:@3625.18]
    assign _T_5150 = _T_5142 & _T_5149; // @[ISA_functions.scala 126:452:@3626.18]
    assign _T_5196 = _T_5149 == 1'h0; // @[ISA_functions.scala 129:455:@3672.20]
    assign _T_5197 = _T_5142 & _T_5196; // @[ISA_functions.scala 129:452:@3673.20]
    assign _T_5198 = _GEN_397 == 32'h5; // @[ISA_functions.scala 129:573:@3674.20]
    assign _T_5199 = _GEN_397 == 32'he; // @[ISA_functions.scala 129:599:@3675.20]
    assign _T_5200 = _T_5198 | _T_5199; // @[ISA_functions.scala 129:589:@3676.20]
    assign _T_5201 = _GEN_397 == 32'h21; // @[ISA_functions.scala 129:627:@3677.20]
    assign _T_5202 = _T_5200 | _T_5201; // @[ISA_functions.scala 129:617:@3678.20]
    assign _T_5203 = _GEN_397 == 32'h22; // @[ISA_functions.scala 129:654:@3679.20]
    assign _T_5204 = _T_5202 | _T_5203; // @[ISA_functions.scala 129:644:@3680.20]
    assign _T_5205 = _T_5197 & _T_5204; // @[ISA_functions.scala 129:560:@3681.20]
    assign _T_5261 = _T_5204 == 1'h0; // @[ISA_functions.scala 132:563:@3736.22]
    assign _T_5262 = _T_5197 & _T_5261; // @[ISA_functions.scala 132:560:@3737.22]
    assign _T_5263 = _GEN_397 == 32'h6; // @[ISA_functions.scala 132:683:@3738.22]
    assign _T_5264 = _GEN_397 == 32'hf; // @[ISA_functions.scala 132:708:@3739.22]
    assign _T_5265 = _T_5263 | _T_5264; // @[ISA_functions.scala 132:698:@3740.22]
    assign _T_5266 = _T_5262 & _T_5265; // @[ISA_functions.scala 132:672:@3741.22]
    assign _T_5328 = _T_5265 == 1'h0; // @[ISA_functions.scala 135:675:@3801.24]
    assign _T_5329 = _T_5262 & _T_5328; // @[ISA_functions.scala 135:672:@3802.24]
    assign _T_5330 = _GEN_397 == 32'h7; // @[ISA_functions.scala 135:737:@3803.24]
    assign _T_5331 = _GEN_397 == 32'h10; // @[ISA_functions.scala 135:762:@3804.24]
    assign _T_5332 = _T_5330 | _T_5331; // @[ISA_functions.scala 135:752:@3805.24]
    assign _T_5333 = _T_5329 & _T_5332; // @[ISA_functions.scala 135:726:@3806.24]
    assign _T_5401 = _T_5332 == 1'h0; // @[ISA_functions.scala 138:729:@3871.26]
    assign _T_5402 = _T_5329 & _T_5401; // @[ISA_functions.scala 138:726:@3872.26]
    assign _T_5403 = _GEN_397 == 32'h8; // @[ISA_functions.scala 138:791:@3873.26]
    assign _T_5404 = _GEN_397 == 32'h11; // @[ISA_functions.scala 138:816:@3874.26]
    assign _T_5405 = _T_5403 | _T_5404; // @[ISA_functions.scala 138:806:@3875.26]
    assign _T_5406 = _T_5402 & _T_5405; // @[ISA_functions.scala 138:780:@3876.26]
    assign _T_5480 = _T_5405 == 1'h0; // @[ISA_functions.scala 141:783:@3946.28]
    assign _T_5481 = _T_5402 & _T_5480; // @[ISA_functions.scala 141:780:@3947.28]
    assign _T_5482 = _GEN_397 == 32'h9; // @[ISA_functions.scala 141:845:@3948.28]
    assign _T_5483 = _GEN_397 == 32'h12; // @[ISA_functions.scala 141:869:@3949.28]
    assign _T_5484 = _T_5482 | _T_5483; // @[ISA_functions.scala 141:859:@3950.28]
    assign _T_5485 = _T_5481 & _T_5484; // @[ISA_functions.scala 141:834:@3951.28]
    assign _T_5565 = _T_5484 == 1'h0; // @[ISA_functions.scala 144:837:@4026.30]
    assign _T_5566 = _T_5481 & _T_5565; // @[ISA_functions.scala 144:834:@4027.30]
    assign _T_5567 = _GEN_397 == 32'ha; // @[ISA_functions.scala 144:897:@4028.30]
    assign _T_5568 = _GEN_397 == 32'h13; // @[ISA_functions.scala 144:922:@4029.30]
    assign _T_5569 = _T_5567 | _T_5568; // @[ISA_functions.scala 144:912:@4030.30]
    assign _T_5570 = _T_5566 & _T_5569; // @[ISA_functions.scala 144:886:@4031.30]
    assign _T_5656 = _T_5569 == 1'h0; // @[ISA_functions.scala 147:889:@4111.32]
    assign _T_5657 = _T_5566 & _T_5656; // @[ISA_functions.scala 147:886:@4112.32]
    assign _T_5658 = _GEN_397 == 32'h19; // @[ISA_functions.scala 147:951:@4113.32]
    assign _T_5659 = _GEN_397 == 32'h25; // @[ISA_functions.scala 147:977:@4114.32]
    assign _T_5660 = _T_5658 | _T_5659; // @[ISA_functions.scala 147:967:@4115.32]
    assign _T_5661 = _T_5657 & _T_5660; // @[ISA_functions.scala 147:940:@4116.32]
    assign _T_5753 = _T_5660 == 1'h0; // @[ISA_functions.scala 150:943:@4201.34]
    assign _T_5754 = _T_5657 & _T_5753; // @[ISA_functions.scala 150:940:@4202.34]
    assign _T_5755 = _GEN_397 == 32'h23; // @[ISA_functions.scala 150:1004:@4203.34]
    assign _T_5756 = _T_5754 & _T_5755; // @[ISA_functions.scala 150:994:@4204.34]
    assign _GEN_398 = _T_5756 ? 32'hb : 32'h0; // @[ISA_functions.scala 150:1020:@4205.34]
    assign _GEN_399 = _T_5661 ? 32'h0 : _GEN_398; // @[ISA_functions.scala 147:994:@4117.32]
    assign _GEN_400 = _T_5570 ? 32'h6 : _GEN_399; // @[ISA_functions.scala 144:940:@4032.30]
    assign _GEN_401 = _T_5485 ? 32'h7 : _GEN_400; // @[ISA_functions.scala 141:886:@3952.28]
    assign _GEN_402 = _T_5406 ? 32'h5 : _GEN_401; // @[ISA_functions.scala 138:834:@3877.26]
    assign _GEN_403 = _T_5333 ? 32'h4 : _GEN_402; // @[ISA_functions.scala 135:780:@3807.24]
    assign _GEN_404 = _T_5266 ? 32'h8 : _GEN_403; // @[ISA_functions.scala 132:726:@3742.22]
    assign _GEN_405 = _T_5205 ? 32'ha : _GEN_404; // @[ISA_functions.scala 129:672:@3682.20]
    assign _GEN_406 = _T_5150 ? 32'h9 : _GEN_405; // @[ISA_functions.scala 126:560:@3627.18]
    assign _GEN_407 = _T_5105 ? 32'h3 : _GEN_406; // @[ISA_functions.scala 123:452:@3581.16]
    assign _GEN_408 = _T_5070 ? 32'h2 : _GEN_407; // @[ISA_functions.scala 120:398:@3544.14]
    assign _GEN_409 = _T_5029 ? 32'h1 : _GEN_408; // @[ISA_functions.scala 117:313:@3512.12]
    assign _T_5782 = _T_2313 | _T_185; // @[ISA_functions.scala 463:224:@4225.12]
    assign _T_5787 = _T_5782 | _T_224; // @[ISA_functions.scala 463:274:@4228.12]
    assign _T_5789 = io_fromMemoryPort_loadedData >> 32'hf; // @[ISA_functions.scala 464:48:@4230.14]
    assign _T_5792 = _T_5789 & 32'h1f; // @[ISA_functions.scala 464:70:@4232.14]
    assign _GEN_410 = _T_5787 ? _T_5792 : 32'h0; // @[ISA_functions.scala 463:325:@4229.12]
    assign _T_5797 = _GEN_410 == 32'h0; // @[ISA_functions.scala 485:28:@4239.12]
    assign _T_5802 = _T_5797 == 1'h0; // @[ISA_functions.scala 488:28:@4245.14]
    assign _T_5804 = _GEN_410 == 32'h1; // @[ISA_functions.scala 488:57:@4246.14]
    assign _T_5805 = _T_5802 & _T_5804; // @[ISA_functions.scala 488:49:@4247.14]
    assign _T_5813 = _T_5804 == 1'h0; // @[ISA_functions.scala 491:52:@4255.16]
    assign _T_5814 = _T_5802 & _T_5813; // @[ISA_functions.scala 491:49:@4256.16]
    assign _T_5816 = _GEN_410 == 32'h2; // @[ISA_functions.scala 491:81:@4257.16]
    assign _T_5817 = _T_5814 & _T_5816; // @[ISA_functions.scala 491:73:@4258.16]
    assign _T_5830 = _T_5816 == 1'h0; // @[ISA_functions.scala 494:76:@4269.18]
    assign _T_5831 = _T_5814 & _T_5830; // @[ISA_functions.scala 494:73:@4270.18]
    assign _T_5833 = _GEN_410 == 32'h3; // @[ISA_functions.scala 494:105:@4271.18]
    assign _T_5834 = _T_5831 & _T_5833; // @[ISA_functions.scala 494:97:@4272.18]
    assign _T_5852 = _T_5833 == 1'h0; // @[ISA_functions.scala 497:100:@4286.20]
    assign _T_5853 = _T_5831 & _T_5852; // @[ISA_functions.scala 497:97:@4287.20]
    assign _T_5855 = _GEN_410 == 32'h4; // @[ISA_functions.scala 497:129:@4288.20]
    assign _T_5856 = _T_5853 & _T_5855; // @[ISA_functions.scala 497:121:@4289.20]
    assign _T_5879 = _T_5855 == 1'h0; // @[ISA_functions.scala 500:124:@4306.22]
    assign _T_5880 = _T_5853 & _T_5879; // @[ISA_functions.scala 500:121:@4307.22]
    assign _T_5882 = _GEN_410 == 32'h5; // @[ISA_functions.scala 500:153:@4308.22]
    assign _T_5883 = _T_5880 & _T_5882; // @[ISA_functions.scala 500:145:@4309.22]
    assign _T_5911 = _T_5882 == 1'h0; // @[ISA_functions.scala 503:148:@4329.24]
    assign _T_5912 = _T_5880 & _T_5911; // @[ISA_functions.scala 503:145:@4330.24]
    assign _T_5914 = _GEN_410 == 32'h6; // @[ISA_functions.scala 503:177:@4331.24]
    assign _T_5915 = _T_5912 & _T_5914; // @[ISA_functions.scala 503:169:@4332.24]
    assign _T_5948 = _T_5914 == 1'h0; // @[ISA_functions.scala 506:172:@4355.26]
    assign _T_5949 = _T_5912 & _T_5948; // @[ISA_functions.scala 506:169:@4356.26]
    assign _T_5951 = _GEN_410 == 32'h7; // @[ISA_functions.scala 506:201:@4357.26]
    assign _T_5952 = _T_5949 & _T_5951; // @[ISA_functions.scala 506:193:@4358.26]
    assign _T_5990 = _T_5951 == 1'h0; // @[ISA_functions.scala 509:196:@4384.28]
    assign _T_5991 = _T_5949 & _T_5990; // @[ISA_functions.scala 509:193:@4385.28]
    assign _T_5993 = _GEN_410 == 32'h8; // @[ISA_functions.scala 509:225:@4386.28]
    assign _T_5994 = _T_5991 & _T_5993; // @[ISA_functions.scala 509:217:@4387.28]
    assign _T_6037 = _T_5993 == 1'h0; // @[ISA_functions.scala 512:220:@4416.30]
    assign _T_6038 = _T_5991 & _T_6037; // @[ISA_functions.scala 512:217:@4417.30]
    assign _T_6040 = _GEN_410 == 32'h9; // @[ISA_functions.scala 512:249:@4418.30]
    assign _T_6041 = _T_6038 & _T_6040; // @[ISA_functions.scala 512:241:@4419.30]
    assign _T_6089 = _T_6040 == 1'h0; // @[ISA_functions.scala 515:244:@4451.32]
    assign _T_6090 = _T_6038 & _T_6089; // @[ISA_functions.scala 515:241:@4452.32]
    assign _T_6092 = _GEN_410 == 32'ha; // @[ISA_functions.scala 515:273:@4453.32]
    assign _T_6093 = _T_6090 & _T_6092; // @[ISA_functions.scala 515:265:@4454.32]
    assign _T_6146 = _T_6092 == 1'h0; // @[ISA_functions.scala 518:268:@4489.34]
    assign _T_6147 = _T_6090 & _T_6146; // @[ISA_functions.scala 518:265:@4490.34]
    assign _T_6149 = _GEN_410 == 32'hb; // @[ISA_functions.scala 518:298:@4491.34]
    assign _T_6150 = _T_6147 & _T_6149; // @[ISA_functions.scala 518:290:@4492.34]
    assign _T_6208 = _T_6149 == 1'h0; // @[ISA_functions.scala 521:293:@4530.36]
    assign _T_6209 = _T_6147 & _T_6208; // @[ISA_functions.scala 521:290:@4531.36]
    assign _T_6211 = _GEN_410 == 32'hc; // @[ISA_functions.scala 521:323:@4532.36]
    assign _T_6212 = _T_6209 & _T_6211; // @[ISA_functions.scala 521:315:@4533.36]
    assign _T_6275 = _T_6211 == 1'h0; // @[ISA_functions.scala 524:318:@4574.38]
    assign _T_6276 = _T_6209 & _T_6275; // @[ISA_functions.scala 524:315:@4575.38]
    assign _T_6278 = _GEN_410 == 32'hd; // @[ISA_functions.scala 524:348:@4576.38]
    assign _T_6279 = _T_6276 & _T_6278; // @[ISA_functions.scala 524:340:@4577.38]
    assign _T_6347 = _T_6278 == 1'h0; // @[ISA_functions.scala 527:343:@4621.40]
    assign _T_6348 = _T_6276 & _T_6347; // @[ISA_functions.scala 527:340:@4622.40]
    assign _T_6350 = _GEN_410 == 32'he; // @[ISA_functions.scala 527:373:@4623.40]
    assign _T_6351 = _T_6348 & _T_6350; // @[ISA_functions.scala 527:365:@4624.40]
    assign _T_6424 = _T_6350 == 1'h0; // @[ISA_functions.scala 530:368:@4671.42]
    assign _T_6425 = _T_6348 & _T_6424; // @[ISA_functions.scala 530:365:@4672.42]
    assign _T_6427 = _GEN_410 == 32'hf; // @[ISA_functions.scala 530:398:@4673.42]
    assign _T_6428 = _T_6425 & _T_6427; // @[ISA_functions.scala 530:390:@4674.42]
    assign _T_6506 = _T_6427 == 1'h0; // @[ISA_functions.scala 533:393:@4724.44]
    assign _T_6507 = _T_6425 & _T_6506; // @[ISA_functions.scala 533:390:@4725.44]
    assign _T_6509 = _GEN_410 == 32'h10; // @[ISA_functions.scala 533:423:@4726.44]
    assign _T_6510 = _T_6507 & _T_6509; // @[ISA_functions.scala 533:415:@4727.44]
    assign _T_6593 = _T_6509 == 1'h0; // @[ISA_functions.scala 536:418:@4780.46]
    assign _T_6594 = _T_6507 & _T_6593; // @[ISA_functions.scala 536:415:@4781.46]
    assign _T_6596 = _GEN_410 == 32'h11; // @[ISA_functions.scala 536:448:@4782.46]
    assign _T_6597 = _T_6594 & _T_6596; // @[ISA_functions.scala 536:440:@4783.46]
    assign _T_6685 = _T_6596 == 1'h0; // @[ISA_functions.scala 539:443:@4839.48]
    assign _T_6686 = _T_6594 & _T_6685; // @[ISA_functions.scala 539:440:@4840.48]
    assign _T_6688 = _GEN_410 == 32'h12; // @[ISA_functions.scala 539:473:@4841.48]
    assign _T_6689 = _T_6686 & _T_6688; // @[ISA_functions.scala 539:465:@4842.48]
    assign _T_6782 = _T_6688 == 1'h0; // @[ISA_functions.scala 542:468:@4901.50]
    assign _T_6783 = _T_6686 & _T_6782; // @[ISA_functions.scala 542:465:@4902.50]
    assign _T_6785 = _GEN_410 == 32'h13; // @[ISA_functions.scala 542:498:@4903.50]
    assign _T_6786 = _T_6783 & _T_6785; // @[ISA_functions.scala 542:490:@4904.50]
    assign _T_6884 = _T_6785 == 1'h0; // @[ISA_functions.scala 545:493:@4966.52]
    assign _T_6885 = _T_6783 & _T_6884; // @[ISA_functions.scala 545:490:@4967.52]
    assign _T_6887 = _GEN_410 == 32'h14; // @[ISA_functions.scala 545:523:@4968.52]
    assign _T_6888 = _T_6885 & _T_6887; // @[ISA_functions.scala 545:515:@4969.52]
    assign _T_6991 = _T_6887 == 1'h0; // @[ISA_functions.scala 548:518:@5034.54]
    assign _T_6992 = _T_6885 & _T_6991; // @[ISA_functions.scala 548:515:@5035.54]
    assign _T_6994 = _GEN_410 == 32'h15; // @[ISA_functions.scala 548:548:@5036.54]
    assign _T_6995 = _T_6992 & _T_6994; // @[ISA_functions.scala 548:540:@5037.54]
    assign _T_7103 = _T_6994 == 1'h0; // @[ISA_functions.scala 551:543:@5105.56]
    assign _T_7104 = _T_6992 & _T_7103; // @[ISA_functions.scala 551:540:@5106.56]
    assign _T_7106 = _GEN_410 == 32'h16; // @[ISA_functions.scala 551:573:@5107.56]
    assign _T_7107 = _T_7104 & _T_7106; // @[ISA_functions.scala 551:565:@5108.56]
    assign _T_7220 = _T_7106 == 1'h0; // @[ISA_functions.scala 554:568:@5179.58]
    assign _T_7221 = _T_7104 & _T_7220; // @[ISA_functions.scala 554:565:@5180.58]
    assign _T_7223 = _GEN_410 == 32'h17; // @[ISA_functions.scala 554:598:@5181.58]
    assign _T_7224 = _T_7221 & _T_7223; // @[ISA_functions.scala 554:590:@5182.58]
    assign _T_7342 = _T_7223 == 1'h0; // @[ISA_functions.scala 557:593:@5256.60]
    assign _T_7343 = _T_7221 & _T_7342; // @[ISA_functions.scala 557:590:@5257.60]
    assign _T_7345 = _GEN_410 == 32'h18; // @[ISA_functions.scala 557:623:@5258.60]
    assign _T_7346 = _T_7343 & _T_7345; // @[ISA_functions.scala 557:615:@5259.60]
    assign _T_7469 = _T_7345 == 1'h0; // @[ISA_functions.scala 560:618:@5336.62]
    assign _T_7470 = _T_7343 & _T_7469; // @[ISA_functions.scala 560:615:@5337.62]
    assign _T_7472 = _GEN_410 == 32'h19; // @[ISA_functions.scala 560:648:@5338.62]
    assign _T_7473 = _T_7470 & _T_7472; // @[ISA_functions.scala 560:640:@5339.62]
    assign _T_7601 = _T_7472 == 1'h0; // @[ISA_functions.scala 563:643:@5419.64]
    assign _T_7602 = _T_7470 & _T_7601; // @[ISA_functions.scala 563:640:@5420.64]
    assign _T_7604 = _GEN_410 == 32'h1a; // @[ISA_functions.scala 563:673:@5421.64]
    assign _T_7605 = _T_7602 & _T_7604; // @[ISA_functions.scala 563:665:@5422.64]
    assign _T_7738 = _T_7604 == 1'h0; // @[ISA_functions.scala 566:668:@5505.66]
    assign _T_7739 = _T_7602 & _T_7738; // @[ISA_functions.scala 566:665:@5506.66]
    assign _T_7741 = _GEN_410 == 32'h1b; // @[ISA_functions.scala 566:698:@5507.66]
    assign _T_7742 = _T_7739 & _T_7741; // @[ISA_functions.scala 566:690:@5508.66]
    assign _T_7880 = _T_7741 == 1'h0; // @[ISA_functions.scala 569:693:@5594.68]
    assign _T_7881 = _T_7739 & _T_7880; // @[ISA_functions.scala 569:690:@5595.68]
    assign _T_7883 = _GEN_410 == 32'h1c; // @[ISA_functions.scala 569:723:@5596.68]
    assign _T_7884 = _T_7881 & _T_7883; // @[ISA_functions.scala 569:715:@5597.68]
    assign _T_8027 = _T_7883 == 1'h0; // @[ISA_functions.scala 572:718:@5686.70]
    assign _T_8028 = _T_7881 & _T_8027; // @[ISA_functions.scala 572:715:@5687.70]
    assign _T_8030 = _GEN_410 == 32'h1d; // @[ISA_functions.scala 572:748:@5688.70]
    assign _T_8031 = _T_8028 & _T_8030; // @[ISA_functions.scala 572:740:@5689.70]
    assign _T_8179 = _T_8030 == 1'h0; // @[ISA_functions.scala 575:743:@5781.72]
    assign _T_8180 = _T_8028 & _T_8179; // @[ISA_functions.scala 575:740:@5782.72]
    assign _T_8182 = _GEN_410 == 32'h1e; // @[ISA_functions.scala 575:773:@5783.72]
    assign _T_8183 = _T_8180 & _T_8182; // @[ISA_functions.scala 575:765:@5784.72]
    assign _GEN_411 = _T_8183 ? io_fromRegsPort_reg_file_30 : io_fromRegsPort_reg_file_31; // @[ISA_functions.scala 575:790:@5785.72]
    assign _GEN_412 = _T_8031 ? io_fromRegsPort_reg_file_29 : _GEN_411; // @[ISA_functions.scala 572:765:@5690.70]
    assign _GEN_413 = _T_7884 ? io_fromRegsPort_reg_file_28 : _GEN_412; // @[ISA_functions.scala 569:740:@5598.68]
    assign _GEN_414 = _T_7742 ? io_fromRegsPort_reg_file_27 : _GEN_413; // @[ISA_functions.scala 566:715:@5509.66]
    assign _GEN_415 = _T_7605 ? io_fromRegsPort_reg_file_26 : _GEN_414; // @[ISA_functions.scala 563:690:@5423.64]
    assign _GEN_416 = _T_7473 ? io_fromRegsPort_reg_file_25 : _GEN_415; // @[ISA_functions.scala 560:665:@5340.62]
    assign _GEN_417 = _T_7346 ? io_fromRegsPort_reg_file_24 : _GEN_416; // @[ISA_functions.scala 557:640:@5260.60]
    assign _GEN_418 = _T_7224 ? io_fromRegsPort_reg_file_23 : _GEN_417; // @[ISA_functions.scala 554:615:@5183.58]
    assign _GEN_419 = _T_7107 ? io_fromRegsPort_reg_file_22 : _GEN_418; // @[ISA_functions.scala 551:590:@5109.56]
    assign _GEN_420 = _T_6995 ? io_fromRegsPort_reg_file_21 : _GEN_419; // @[ISA_functions.scala 548:565:@5038.54]
    assign _GEN_421 = _T_6888 ? io_fromRegsPort_reg_file_20 : _GEN_420; // @[ISA_functions.scala 545:540:@4970.52]
    assign _GEN_422 = _T_6786 ? io_fromRegsPort_reg_file_19 : _GEN_421; // @[ISA_functions.scala 542:515:@4905.50]
    assign _GEN_423 = _T_6689 ? io_fromRegsPort_reg_file_18 : _GEN_422; // @[ISA_functions.scala 539:490:@4843.48]
    assign _GEN_424 = _T_6597 ? io_fromRegsPort_reg_file_17 : _GEN_423; // @[ISA_functions.scala 536:465:@4784.46]
    assign _GEN_425 = _T_6510 ? io_fromRegsPort_reg_file_16 : _GEN_424; // @[ISA_functions.scala 533:440:@4728.44]
    assign _GEN_426 = _T_6428 ? io_fromRegsPort_reg_file_15 : _GEN_425; // @[ISA_functions.scala 530:415:@4675.42]
    assign _GEN_427 = _T_6351 ? io_fromRegsPort_reg_file_14 : _GEN_426; // @[ISA_functions.scala 527:390:@4625.40]
    assign _GEN_428 = _T_6279 ? io_fromRegsPort_reg_file_13 : _GEN_427; // @[ISA_functions.scala 524:365:@4578.38]
    assign _GEN_429 = _T_6212 ? io_fromRegsPort_reg_file_12 : _GEN_428; // @[ISA_functions.scala 521:340:@4534.36]
    assign _GEN_430 = _T_6150 ? io_fromRegsPort_reg_file_11 : _GEN_429; // @[ISA_functions.scala 518:315:@4493.34]
    assign _GEN_431 = _T_6093 ? io_fromRegsPort_reg_file_10 : _GEN_430; // @[ISA_functions.scala 515:290:@4455.32]
    assign _GEN_432 = _T_6041 ? io_fromRegsPort_reg_file_09 : _GEN_431; // @[ISA_functions.scala 512:265:@4420.30]
    assign _GEN_433 = _T_5994 ? io_fromRegsPort_reg_file_08 : _GEN_432; // @[ISA_functions.scala 509:241:@4388.28]
    assign _GEN_434 = _T_5952 ? io_fromRegsPort_reg_file_07 : _GEN_433; // @[ISA_functions.scala 506:217:@4359.26]
    assign _GEN_435 = _T_5915 ? io_fromRegsPort_reg_file_06 : _GEN_434; // @[ISA_functions.scala 503:193:@4333.24]
    assign _GEN_436 = _T_5883 ? io_fromRegsPort_reg_file_05 : _GEN_435; // @[ISA_functions.scala 500:169:@4310.22]
    assign _GEN_437 = _T_5856 ? io_fromRegsPort_reg_file_04 : _GEN_436; // @[ISA_functions.scala 497:145:@4290.20]
    assign _GEN_438 = _T_5834 ? io_fromRegsPort_reg_file_03 : _GEN_437; // @[ISA_functions.scala 494:121:@4273.18]
    assign _GEN_439 = _T_5817 ? io_fromRegsPort_reg_file_02 : _GEN_438; // @[ISA_functions.scala 491:97:@4259.16]
    assign _GEN_440 = _T_5805 ? io_fromRegsPort_reg_file_01 : _GEN_439; // @[ISA_functions.scala 488:73:@4248.14]
    assign _GEN_441 = _T_5797 ? 32'h0 : _GEN_440; // @[ISA_functions.scala 485:44:@4240.12]
    assign _T_8194 = _T_91 | _T_185; // @[ISA_functions.scala 474:71:@5796.12]
    assign _T_8199 = _T_8194 | _T_224; // @[ISA_functions.scala 474:121:@5799.12]
    assign _T_8201 = io_fromMemoryPort_loadedData >> 32'h14; // @[ISA_functions.scala 475:48:@5801.14]
    assign _T_8204 = _T_8201 & 32'h1f; // @[ISA_functions.scala 475:70:@5803.14]
    assign _GEN_442 = _T_8199 ? _T_8204 : 32'h0; // @[ISA_functions.scala 474:172:@5800.12]
    assign _T_8209 = _GEN_442 == 32'h0; // @[ISA_functions.scala 485:28:@5810.12]
    assign _T_8214 = _T_8209 == 1'h0; // @[ISA_functions.scala 488:28:@5816.14]
    assign _T_8216 = _GEN_442 == 32'h1; // @[ISA_functions.scala 488:57:@5817.14]
    assign _T_8217 = _T_8214 & _T_8216; // @[ISA_functions.scala 488:49:@5818.14]
    assign _T_8225 = _T_8216 == 1'h0; // @[ISA_functions.scala 491:52:@5826.16]
    assign _T_8226 = _T_8214 & _T_8225; // @[ISA_functions.scala 491:49:@5827.16]
    assign _T_8228 = _GEN_442 == 32'h2; // @[ISA_functions.scala 491:81:@5828.16]
    assign _T_8229 = _T_8226 & _T_8228; // @[ISA_functions.scala 491:73:@5829.16]
    assign _T_8242 = _T_8228 == 1'h0; // @[ISA_functions.scala 494:76:@5840.18]
    assign _T_8243 = _T_8226 & _T_8242; // @[ISA_functions.scala 494:73:@5841.18]
    assign _T_8245 = _GEN_442 == 32'h3; // @[ISA_functions.scala 494:105:@5842.18]
    assign _T_8246 = _T_8243 & _T_8245; // @[ISA_functions.scala 494:97:@5843.18]
    assign _T_8264 = _T_8245 == 1'h0; // @[ISA_functions.scala 497:100:@5857.20]
    assign _T_8265 = _T_8243 & _T_8264; // @[ISA_functions.scala 497:97:@5858.20]
    assign _T_8267 = _GEN_442 == 32'h4; // @[ISA_functions.scala 497:129:@5859.20]
    assign _T_8268 = _T_8265 & _T_8267; // @[ISA_functions.scala 497:121:@5860.20]
    assign _T_8291 = _T_8267 == 1'h0; // @[ISA_functions.scala 500:124:@5877.22]
    assign _T_8292 = _T_8265 & _T_8291; // @[ISA_functions.scala 500:121:@5878.22]
    assign _T_8294 = _GEN_442 == 32'h5; // @[ISA_functions.scala 500:153:@5879.22]
    assign _T_8295 = _T_8292 & _T_8294; // @[ISA_functions.scala 500:145:@5880.22]
    assign _T_8323 = _T_8294 == 1'h0; // @[ISA_functions.scala 503:148:@5900.24]
    assign _T_8324 = _T_8292 & _T_8323; // @[ISA_functions.scala 503:145:@5901.24]
    assign _T_8326 = _GEN_442 == 32'h6; // @[ISA_functions.scala 503:177:@5902.24]
    assign _T_8327 = _T_8324 & _T_8326; // @[ISA_functions.scala 503:169:@5903.24]
    assign _T_8360 = _T_8326 == 1'h0; // @[ISA_functions.scala 506:172:@5926.26]
    assign _T_8361 = _T_8324 & _T_8360; // @[ISA_functions.scala 506:169:@5927.26]
    assign _T_8363 = _GEN_442 == 32'h7; // @[ISA_functions.scala 506:201:@5928.26]
    assign _T_8364 = _T_8361 & _T_8363; // @[ISA_functions.scala 506:193:@5929.26]
    assign _T_8402 = _T_8363 == 1'h0; // @[ISA_functions.scala 509:196:@5955.28]
    assign _T_8403 = _T_8361 & _T_8402; // @[ISA_functions.scala 509:193:@5956.28]
    assign _T_8405 = _GEN_442 == 32'h8; // @[ISA_functions.scala 509:225:@5957.28]
    assign _T_8406 = _T_8403 & _T_8405; // @[ISA_functions.scala 509:217:@5958.28]
    assign _T_8449 = _T_8405 == 1'h0; // @[ISA_functions.scala 512:220:@5987.30]
    assign _T_8450 = _T_8403 & _T_8449; // @[ISA_functions.scala 512:217:@5988.30]
    assign _T_8452 = _GEN_442 == 32'h9; // @[ISA_functions.scala 512:249:@5989.30]
    assign _T_8453 = _T_8450 & _T_8452; // @[ISA_functions.scala 512:241:@5990.30]
    assign _T_8501 = _T_8452 == 1'h0; // @[ISA_functions.scala 515:244:@6022.32]
    assign _T_8502 = _T_8450 & _T_8501; // @[ISA_functions.scala 515:241:@6023.32]
    assign _T_8504 = _GEN_442 == 32'ha; // @[ISA_functions.scala 515:273:@6024.32]
    assign _T_8505 = _T_8502 & _T_8504; // @[ISA_functions.scala 515:265:@6025.32]
    assign _T_8558 = _T_8504 == 1'h0; // @[ISA_functions.scala 518:268:@6060.34]
    assign _T_8559 = _T_8502 & _T_8558; // @[ISA_functions.scala 518:265:@6061.34]
    assign _T_8561 = _GEN_442 == 32'hb; // @[ISA_functions.scala 518:298:@6062.34]
    assign _T_8562 = _T_8559 & _T_8561; // @[ISA_functions.scala 518:290:@6063.34]
    assign _T_8620 = _T_8561 == 1'h0; // @[ISA_functions.scala 521:293:@6101.36]
    assign _T_8621 = _T_8559 & _T_8620; // @[ISA_functions.scala 521:290:@6102.36]
    assign _T_8623 = _GEN_442 == 32'hc; // @[ISA_functions.scala 521:323:@6103.36]
    assign _T_8624 = _T_8621 & _T_8623; // @[ISA_functions.scala 521:315:@6104.36]
    assign _T_8687 = _T_8623 == 1'h0; // @[ISA_functions.scala 524:318:@6145.38]
    assign _T_8688 = _T_8621 & _T_8687; // @[ISA_functions.scala 524:315:@6146.38]
    assign _T_8690 = _GEN_442 == 32'hd; // @[ISA_functions.scala 524:348:@6147.38]
    assign _T_8691 = _T_8688 & _T_8690; // @[ISA_functions.scala 524:340:@6148.38]
    assign _T_8759 = _T_8690 == 1'h0; // @[ISA_functions.scala 527:343:@6192.40]
    assign _T_8760 = _T_8688 & _T_8759; // @[ISA_functions.scala 527:340:@6193.40]
    assign _T_8762 = _GEN_442 == 32'he; // @[ISA_functions.scala 527:373:@6194.40]
    assign _T_8763 = _T_8760 & _T_8762; // @[ISA_functions.scala 527:365:@6195.40]
    assign _T_8836 = _T_8762 == 1'h0; // @[ISA_functions.scala 530:368:@6242.42]
    assign _T_8837 = _T_8760 & _T_8836; // @[ISA_functions.scala 530:365:@6243.42]
    assign _T_8839 = _GEN_442 == 32'hf; // @[ISA_functions.scala 530:398:@6244.42]
    assign _T_8840 = _T_8837 & _T_8839; // @[ISA_functions.scala 530:390:@6245.42]
    assign _T_8918 = _T_8839 == 1'h0; // @[ISA_functions.scala 533:393:@6295.44]
    assign _T_8919 = _T_8837 & _T_8918; // @[ISA_functions.scala 533:390:@6296.44]
    assign _T_8921 = _GEN_442 == 32'h10; // @[ISA_functions.scala 533:423:@6297.44]
    assign _T_8922 = _T_8919 & _T_8921; // @[ISA_functions.scala 533:415:@6298.44]
    assign _T_9005 = _T_8921 == 1'h0; // @[ISA_functions.scala 536:418:@6351.46]
    assign _T_9006 = _T_8919 & _T_9005; // @[ISA_functions.scala 536:415:@6352.46]
    assign _T_9008 = _GEN_442 == 32'h11; // @[ISA_functions.scala 536:448:@6353.46]
    assign _T_9009 = _T_9006 & _T_9008; // @[ISA_functions.scala 536:440:@6354.46]
    assign _T_9097 = _T_9008 == 1'h0; // @[ISA_functions.scala 539:443:@6410.48]
    assign _T_9098 = _T_9006 & _T_9097; // @[ISA_functions.scala 539:440:@6411.48]
    assign _T_9100 = _GEN_442 == 32'h12; // @[ISA_functions.scala 539:473:@6412.48]
    assign _T_9101 = _T_9098 & _T_9100; // @[ISA_functions.scala 539:465:@6413.48]
    assign _T_9194 = _T_9100 == 1'h0; // @[ISA_functions.scala 542:468:@6472.50]
    assign _T_9195 = _T_9098 & _T_9194; // @[ISA_functions.scala 542:465:@6473.50]
    assign _T_9197 = _GEN_442 == 32'h13; // @[ISA_functions.scala 542:498:@6474.50]
    assign _T_9198 = _T_9195 & _T_9197; // @[ISA_functions.scala 542:490:@6475.50]
    assign _T_9296 = _T_9197 == 1'h0; // @[ISA_functions.scala 545:493:@6537.52]
    assign _T_9297 = _T_9195 & _T_9296; // @[ISA_functions.scala 545:490:@6538.52]
    assign _T_9299 = _GEN_442 == 32'h14; // @[ISA_functions.scala 545:523:@6539.52]
    assign _T_9300 = _T_9297 & _T_9299; // @[ISA_functions.scala 545:515:@6540.52]
    assign _T_9403 = _T_9299 == 1'h0; // @[ISA_functions.scala 548:518:@6605.54]
    assign _T_9404 = _T_9297 & _T_9403; // @[ISA_functions.scala 548:515:@6606.54]
    assign _T_9406 = _GEN_442 == 32'h15; // @[ISA_functions.scala 548:548:@6607.54]
    assign _T_9407 = _T_9404 & _T_9406; // @[ISA_functions.scala 548:540:@6608.54]
    assign _T_9515 = _T_9406 == 1'h0; // @[ISA_functions.scala 551:543:@6676.56]
    assign _T_9516 = _T_9404 & _T_9515; // @[ISA_functions.scala 551:540:@6677.56]
    assign _T_9518 = _GEN_442 == 32'h16; // @[ISA_functions.scala 551:573:@6678.56]
    assign _T_9519 = _T_9516 & _T_9518; // @[ISA_functions.scala 551:565:@6679.56]
    assign _T_9632 = _T_9518 == 1'h0; // @[ISA_functions.scala 554:568:@6750.58]
    assign _T_9633 = _T_9516 & _T_9632; // @[ISA_functions.scala 554:565:@6751.58]
    assign _T_9635 = _GEN_442 == 32'h17; // @[ISA_functions.scala 554:598:@6752.58]
    assign _T_9636 = _T_9633 & _T_9635; // @[ISA_functions.scala 554:590:@6753.58]
    assign _T_9754 = _T_9635 == 1'h0; // @[ISA_functions.scala 557:593:@6827.60]
    assign _T_9755 = _T_9633 & _T_9754; // @[ISA_functions.scala 557:590:@6828.60]
    assign _T_9757 = _GEN_442 == 32'h18; // @[ISA_functions.scala 557:623:@6829.60]
    assign _T_9758 = _T_9755 & _T_9757; // @[ISA_functions.scala 557:615:@6830.60]
    assign _T_9881 = _T_9757 == 1'h0; // @[ISA_functions.scala 560:618:@6907.62]
    assign _T_9882 = _T_9755 & _T_9881; // @[ISA_functions.scala 560:615:@6908.62]
    assign _T_9884 = _GEN_442 == 32'h19; // @[ISA_functions.scala 560:648:@6909.62]
    assign _T_9885 = _T_9882 & _T_9884; // @[ISA_functions.scala 560:640:@6910.62]
    assign _T_10013 = _T_9884 == 1'h0; // @[ISA_functions.scala 563:643:@6990.64]
    assign _T_10014 = _T_9882 & _T_10013; // @[ISA_functions.scala 563:640:@6991.64]
    assign _T_10016 = _GEN_442 == 32'h1a; // @[ISA_functions.scala 563:673:@6992.64]
    assign _T_10017 = _T_10014 & _T_10016; // @[ISA_functions.scala 563:665:@6993.64]
    assign _T_10150 = _T_10016 == 1'h0; // @[ISA_functions.scala 566:668:@7076.66]
    assign _T_10151 = _T_10014 & _T_10150; // @[ISA_functions.scala 566:665:@7077.66]
    assign _T_10153 = _GEN_442 == 32'h1b; // @[ISA_functions.scala 566:698:@7078.66]
    assign _T_10154 = _T_10151 & _T_10153; // @[ISA_functions.scala 566:690:@7079.66]
    assign _T_10292 = _T_10153 == 1'h0; // @[ISA_functions.scala 569:693:@7165.68]
    assign _T_10293 = _T_10151 & _T_10292; // @[ISA_functions.scala 569:690:@7166.68]
    assign _T_10295 = _GEN_442 == 32'h1c; // @[ISA_functions.scala 569:723:@7167.68]
    assign _T_10296 = _T_10293 & _T_10295; // @[ISA_functions.scala 569:715:@7168.68]
    assign _T_10439 = _T_10295 == 1'h0; // @[ISA_functions.scala 572:718:@7257.70]
    assign _T_10440 = _T_10293 & _T_10439; // @[ISA_functions.scala 572:715:@7258.70]
    assign _T_10442 = _GEN_442 == 32'h1d; // @[ISA_functions.scala 572:748:@7259.70]
    assign _T_10443 = _T_10440 & _T_10442; // @[ISA_functions.scala 572:740:@7260.70]
    assign _T_10591 = _T_10442 == 1'h0; // @[ISA_functions.scala 575:743:@7352.72]
    assign _T_10592 = _T_10440 & _T_10591; // @[ISA_functions.scala 575:740:@7353.72]
    assign _T_10594 = _GEN_442 == 32'h1e; // @[ISA_functions.scala 575:773:@7354.72]
    assign _T_10595 = _T_10592 & _T_10594; // @[ISA_functions.scala 575:765:@7355.72]
    assign _GEN_443 = _T_10595 ? io_fromRegsPort_reg_file_30 : io_fromRegsPort_reg_file_31; // @[ISA_functions.scala 575:790:@7356.72]
    assign _GEN_444 = _T_10443 ? io_fromRegsPort_reg_file_29 : _GEN_443; // @[ISA_functions.scala 572:765:@7261.70]
    assign _GEN_445 = _T_10296 ? io_fromRegsPort_reg_file_28 : _GEN_444; // @[ISA_functions.scala 569:740:@7169.68]
    assign _GEN_446 = _T_10154 ? io_fromRegsPort_reg_file_27 : _GEN_445; // @[ISA_functions.scala 566:715:@7080.66]
    assign _GEN_447 = _T_10017 ? io_fromRegsPort_reg_file_26 : _GEN_446; // @[ISA_functions.scala 563:690:@6994.64]
    assign _GEN_448 = _T_9885 ? io_fromRegsPort_reg_file_25 : _GEN_447; // @[ISA_functions.scala 560:665:@6911.62]
    assign _GEN_449 = _T_9758 ? io_fromRegsPort_reg_file_24 : _GEN_448; // @[ISA_functions.scala 557:640:@6831.60]
    assign _GEN_450 = _T_9636 ? io_fromRegsPort_reg_file_23 : _GEN_449; // @[ISA_functions.scala 554:615:@6754.58]
    assign _GEN_451 = _T_9519 ? io_fromRegsPort_reg_file_22 : _GEN_450; // @[ISA_functions.scala 551:590:@6680.56]
    assign _GEN_452 = _T_9407 ? io_fromRegsPort_reg_file_21 : _GEN_451; // @[ISA_functions.scala 548:565:@6609.54]
    assign _GEN_453 = _T_9300 ? io_fromRegsPort_reg_file_20 : _GEN_452; // @[ISA_functions.scala 545:540:@6541.52]
    assign _GEN_454 = _T_9198 ? io_fromRegsPort_reg_file_19 : _GEN_453; // @[ISA_functions.scala 542:515:@6476.50]
    assign _GEN_455 = _T_9101 ? io_fromRegsPort_reg_file_18 : _GEN_454; // @[ISA_functions.scala 539:490:@6414.48]
    assign _GEN_456 = _T_9009 ? io_fromRegsPort_reg_file_17 : _GEN_455; // @[ISA_functions.scala 536:465:@6355.46]
    assign _GEN_457 = _T_8922 ? io_fromRegsPort_reg_file_16 : _GEN_456; // @[ISA_functions.scala 533:440:@6299.44]
    assign _GEN_458 = _T_8840 ? io_fromRegsPort_reg_file_15 : _GEN_457; // @[ISA_functions.scala 530:415:@6246.42]
    assign _GEN_459 = _T_8763 ? io_fromRegsPort_reg_file_14 : _GEN_458; // @[ISA_functions.scala 527:390:@6196.40]
    assign _GEN_460 = _T_8691 ? io_fromRegsPort_reg_file_13 : _GEN_459; // @[ISA_functions.scala 524:365:@6149.38]
    assign _GEN_461 = _T_8624 ? io_fromRegsPort_reg_file_12 : _GEN_460; // @[ISA_functions.scala 521:340:@6105.36]
    assign _GEN_462 = _T_8562 ? io_fromRegsPort_reg_file_11 : _GEN_461; // @[ISA_functions.scala 518:315:@6064.34]
    assign _GEN_463 = _T_8505 ? io_fromRegsPort_reg_file_10 : _GEN_462; // @[ISA_functions.scala 515:290:@6026.32]
    assign _GEN_464 = _T_8453 ? io_fromRegsPort_reg_file_09 : _GEN_463; // @[ISA_functions.scala 512:265:@5991.30]
    assign _GEN_465 = _T_8406 ? io_fromRegsPort_reg_file_08 : _GEN_464; // @[ISA_functions.scala 509:241:@5959.28]
    assign _GEN_466 = _T_8364 ? io_fromRegsPort_reg_file_07 : _GEN_465; // @[ISA_functions.scala 506:217:@5930.26]
    assign _GEN_467 = _T_8327 ? io_fromRegsPort_reg_file_06 : _GEN_466; // @[ISA_functions.scala 503:193:@5904.24]
    assign _GEN_468 = _T_8295 ? io_fromRegsPort_reg_file_05 : _GEN_467; // @[ISA_functions.scala 500:169:@5881.22]
    assign _GEN_469 = _T_8268 ? io_fromRegsPort_reg_file_04 : _GEN_468; // @[ISA_functions.scala 497:145:@5861.20]
    assign _GEN_470 = _T_8246 ? io_fromRegsPort_reg_file_03 : _GEN_469; // @[ISA_functions.scala 494:121:@5844.18]
    assign _GEN_471 = _T_8229 ? io_fromRegsPort_reg_file_02 : _GEN_470; // @[ISA_functions.scala 491:97:@5830.16]
    assign _GEN_472 = _T_8217 ? io_fromRegsPort_reg_file_01 : _GEN_471; // @[ISA_functions.scala 488:73:@5819.14]
    assign _GEN_473 = _T_8209 ? 32'h0 : _GEN_472; // @[ISA_functions.scala 485:44:@5811.12]
    assign _T_10598 = _GEN_409 == 32'h1; // @[ISA_functions.scala 161:36:@7363.12]
    assign _T_10599 = _GEN_441 + _GEN_473; // @[ISA_functions.scala 162:43:@7365.14]
    assign _T_10600 = _GEN_441 + _GEN_473; // @[ISA_functions.scala 162:43:@7366.14]
    assign _T_10603 = _T_10598 == 1'h0; // @[ISA_functions.scala 164:28:@7371.14]
    assign _T_10604 = _GEN_409 == 32'h2; // @[ISA_functions.scala 164:71:@7372.14]
    assign _T_10605 = _T_10603 & _T_10604; // @[ISA_functions.scala 164:55:@7373.14]
    assign _T_10607 = _GEN_473 * 32'hffffffff; // @[ISA_functions.scala 165:55:@7375.16]
    assign _GEN_6225 = {{32'd0}, _GEN_441}; // @[ISA_functions.scala 165:43:@7376.16]
    assign _T_10608 = _GEN_6225 + _T_10607; // @[ISA_functions.scala 165:43:@7376.16]
    assign _T_10609 = _GEN_6225 + _T_10607; // @[ISA_functions.scala 165:43:@7377.16]
    assign _T_10615 = _T_10604 == 1'h0; // @[ISA_functions.scala 167:58:@7384.16]
    assign _T_10616 = _T_10603 & _T_10615; // @[ISA_functions.scala 167:55:@7385.16]
    assign _T_10617 = _GEN_409 == 32'h6; // @[ISA_functions.scala 167:101:@7386.16]
    assign _T_10618 = _T_10616 & _T_10617; // @[ISA_functions.scala 167:85:@7387.16]
    assign _T_10619 = _GEN_441 & _GEN_473; // @[ISA_functions.scala 168:43:@7389.18]
    assign _T_10629 = _T_10617 == 1'h0; // @[ISA_functions.scala 170:88:@7399.18]
    assign _T_10630 = _T_10616 & _T_10629; // @[ISA_functions.scala 170:85:@7400.18]
    assign _T_10631 = _GEN_409 == 32'h7; // @[ISA_functions.scala 170:131:@7401.18]
    assign _T_10632 = _T_10630 & _T_10631; // @[ISA_functions.scala 170:115:@7402.18]
    assign _T_10633 = _GEN_441 | _GEN_473; // @[ISA_functions.scala 171:43:@7404.20]
    assign _T_10647 = _T_10631 == 1'h0; // @[ISA_functions.scala 173:118:@7417.20]
    assign _T_10648 = _T_10630 & _T_10647; // @[ISA_functions.scala 173:115:@7418.20]
    assign _T_10649 = _GEN_409 == 32'h8; // @[ISA_functions.scala 173:160:@7419.20]
    assign _T_10650 = _T_10648 & _T_10649; // @[ISA_functions.scala 173:144:@7420.20]
    assign _T_10651 = _GEN_441 ^ _GEN_473; // @[ISA_functions.scala 174:43:@7422.22]
    assign _T_10669 = _T_10649 == 1'h0; // @[ISA_functions.scala 176:147:@7438.22]
    assign _T_10670 = _T_10648 & _T_10669; // @[ISA_functions.scala 176:144:@7439.22]
    assign _T_10671 = _GEN_409 == 32'h9; // @[ISA_functions.scala 176:190:@7440.22]
    assign _T_10672 = _T_10670 & _T_10671; // @[ISA_functions.scala 176:174:@7441.22]
    assign _T_10673 = $signed(_GEN_441); // @[ISA_functions.scala 176:217:@7442.22]
    assign _T_10674 = $signed(_GEN_473); // @[ISA_functions.scala 176:237:@7443.22]
    assign _T_10675 = $signed(_T_10673) < $signed(_T_10674); // @[ISA_functions.scala 176:225:@7444.22]
    assign _T_10676 = _T_10672 & _T_10675; // @[ISA_functions.scala 176:203:@7445.22]
    assign _T_10703 = _T_10675 == 1'h0; // @[ISA_functions.scala 179:206:@7469.24]
    assign _T_10704 = _T_10672 & _T_10703; // @[ISA_functions.scala 179:203:@7470.24]
    assign _T_10727 = _T_10671 == 1'h0; // @[ISA_functions.scala 182:177:@7490.26]
    assign _T_10728 = _T_10670 & _T_10727; // @[ISA_functions.scala 182:174:@7491.26]
    assign _T_10729 = _GEN_409 == 32'ha; // @[ISA_functions.scala 182:220:@7492.26]
    assign _T_10730 = _T_10728 & _T_10729; // @[ISA_functions.scala 182:204:@7493.26]
    assign _T_10731 = _GEN_441 < _GEN_473; // @[ISA_functions.scala 182:247:@7494.26]
    assign _T_10732 = _T_10730 & _T_10731; // @[ISA_functions.scala 182:234:@7495.26]
    assign _T_10761 = _T_10731 == 1'h0; // @[ISA_functions.scala 185:237:@7520.28]
    assign _T_10762 = _T_10730 & _T_10761; // @[ISA_functions.scala 185:234:@7521.28]
    assign _T_10789 = _T_10729 == 1'h0; // @[ISA_functions.scala 188:207:@7544.30]
    assign _T_10790 = _T_10728 & _T_10789; // @[ISA_functions.scala 188:204:@7545.30]
    assign _T_10791 = _GEN_409 == 32'h3; // @[ISA_functions.scala 188:251:@7546.30]
    assign _T_10792 = _T_10790 & _T_10791; // @[ISA_functions.scala 188:235:@7547.30]
    assign _T_10793 = _GEN_473[18:0]; // @[ISA_functions.scala 189:55:@7549.32]
    assign _T_10795 = _T_10793 & 19'h1f; // @[ISA_functions.scala 189:62:@7550.32]
    assign _GEN_6226 = {{524287'd0}, _GEN_441}; // @[ISA_functions.scala 189:43:@7551.32]
    assign _T_10796 = _GEN_6226 << _T_10795; // @[ISA_functions.scala 189:43:@7551.32]
    assign _T_10797 = _T_10796[31:0]; // @[ISA_functions.scala 189:76:@7552.32]
    assign _T_10827 = _T_10791 == 1'h0; // @[ISA_functions.scala 191:238:@7577.32]
    assign _T_10828 = _T_10790 & _T_10827; // @[ISA_functions.scala 191:235:@7578.32]
    assign _T_10829 = _GEN_409 == 32'h5; // @[ISA_functions.scala 191:281:@7579.32]
    assign _T_10830 = _T_10828 & _T_10829; // @[ISA_functions.scala 191:265:@7580.32]
    assign _T_10833 = _GEN_473 & 32'h1f; // @[ISA_functions.scala 192:67:@7583.34]
    assign _T_10834 = $signed(_T_10673) >>> _T_10833; // @[ISA_functions.scala 192:53:@7584.34]
    assign _T_10835 = $unsigned(_T_10834); // @[ISA_functions.scala 192:82:@7585.34]
    assign _T_10869 = _T_10829 == 1'h0; // @[ISA_functions.scala 194:268:@7613.34]
    assign _T_10870 = _T_10828 & _T_10869; // @[ISA_functions.scala 194:265:@7614.34]
    assign _T_10871 = _GEN_409 == 32'h4; // @[ISA_functions.scala 194:311:@7615.34]
    assign _T_10872 = _T_10870 & _T_10871; // @[ISA_functions.scala 194:295:@7616.34]
    assign _T_10875 = _GEN_441 >> _T_10833; // @[ISA_functions.scala 195:43:@7619.36]
    assign _T_10914 = _T_10871 == 1'h0; // @[ISA_functions.scala 197:298:@7651.36]
    assign _T_10915 = _T_10870 & _T_10914; // @[ISA_functions.scala 197:295:@7652.36]
    assign _T_10916 = _GEN_409 == 32'hb; // @[ISA_functions.scala 197:341:@7653.36]
    assign _T_10917 = _T_10915 & _T_10916; // @[ISA_functions.scala 197:325:@7654.36]
    assign _GEN_474 = _T_10917 ? _GEN_441 : 32'h0; // @[ISA_functions.scala 197:357:@7655.36]
    assign _GEN_475 = _T_10872 ? _T_10875 : _GEN_474; // @[ISA_functions.scala 194:325:@7617.34]
    assign _GEN_476 = _T_10830 ? _T_10835 : _GEN_475; // @[ISA_functions.scala 191:295:@7581.32]
    assign _GEN_477 = _T_10792 ? _T_10797 : _GEN_476; // @[ISA_functions.scala 188:265:@7548.30]
    assign _GEN_478 = _T_10762 ? 32'h0 : _GEN_477; // @[ISA_functions.scala 185:261:@7522.28]
    assign _GEN_479 = _T_10732 ? 32'h1 : _GEN_478; // @[ISA_functions.scala 182:260:@7496.26]
    assign _GEN_480 = _T_10704 ? 32'h0 : _GEN_479; // @[ISA_functions.scala 179:248:@7471.24]
    assign _GEN_481 = _T_10676 ? 32'h1 : _GEN_480; // @[ISA_functions.scala 176:247:@7446.22]
    assign _GEN_482 = _T_10650 ? _T_10651 : _GEN_481; // @[ISA_functions.scala 173:174:@7421.20]
    assign _GEN_483 = _T_10632 ? _T_10633 : _GEN_482; // @[ISA_functions.scala 170:144:@7403.18]
    assign _GEN_484 = _T_10618 ? _T_10619 : _GEN_483; // @[ISA_functions.scala 167:115:@7388.16]
    assign _GEN_485 = _T_10605 ? _T_10609 : {{32'd0}, _GEN_484}; // @[ISA_functions.scala 164:85:@7374.14]
    assign _GEN_486 = _T_10598 ? {{32'd0}, _T_10600} : _GEN_485; // @[ISA_functions.scala 161:50:@7364.12]
    assign _GEN_622 = io_fromMemoryPort_sync ? 3'h4 : _GEN_329; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_623 = io_fromMemoryPort_sync ? _T_50 : _GEN_330; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_624 = io_fromMemoryPort_sync ? 32'h0 : _GEN_331; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_625 = io_fromMemoryPort_sync ? 32'h1 : _GEN_332; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_626 = io_fromMemoryPort_sync ? 32'h1 : _GEN_333; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_627 = io_fromMemoryPort_sync ? _T_50 : _GEN_334; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_628 = io_fromMemoryPort_sync ? _GEN_352 : regfileWrite_signal_r_dst; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_629 = io_fromMemoryPort_sync ? _GEN_486 : {{32'd0}, _GEN_336}; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_630 = io_fromMemoryPort_sync ? _T_50 : _GEN_337; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_631 = io_fromMemoryPort_sync ? 32'h0 : _GEN_338; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_632 = io_fromMemoryPort_sync ? 32'h1 : _GEN_339; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_633 = io_fromMemoryPort_sync ? 32'h1 : _GEN_340; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_634 = io_fromMemoryPort_sync ? _GEN_352 : _GEN_103; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_635 = io_fromMemoryPort_sync ? _GEN_486 : {{32'd0}, _GEN_104}; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_636 = io_fromMemoryPort_sync ? 1'h0 : _GEN_341; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_637 = io_fromMemoryPort_sync ? 1'h1 : _GEN_342; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_638 = io_fromMemoryPort_sync ? 1'h1 : _GEN_343; // @[ISA.scala 227:62:@1715.10]
    assign _GEN_639 = _T_335 ? _GEN_622 : _GEN_329; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_640 = _T_335 ? _GEN_623 : _GEN_330; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_641 = _T_335 ? _GEN_624 : _GEN_331; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_642 = _T_335 ? _GEN_625 : _GEN_332; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_643 = _T_335 ? _GEN_626 : _GEN_333; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_644 = _T_335 ? _GEN_627 : _GEN_334; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_645 = _T_335 ? _GEN_628 : regfileWrite_signal_r_dst; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_646 = _T_335 ? _GEN_629 : {{32'd0}, _GEN_336}; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_647 = _T_335 ? _GEN_630 : _GEN_337; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_648 = _T_335 ? _GEN_631 : _GEN_338; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_649 = _T_335 ? _GEN_632 : _GEN_339; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_650 = _T_335 ? _GEN_633 : _GEN_340; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_651 = _T_335 ? _GEN_634 : _GEN_103; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_652 = _T_335 ? _GEN_635 : {{32'd0}, _GEN_104}; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_653 = _T_335 ? _GEN_636 : _GEN_341; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_654 = _T_335 ? _GEN_637 : _GEN_342; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_655 = _T_335 ? _GEN_638 : _GEN_343; // @[ISA.scala 226:84:@1714.8]
    assign _GEN_656 = _T_85 ? _GEN_639 : _GEN_329; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_657 = _T_85 ? _GEN_640 : _GEN_330; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_658 = _T_85 ? _GEN_641 : _GEN_331; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_659 = _T_85 ? _GEN_642 : _GEN_332; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_660 = _T_85 ? _GEN_643 : _GEN_333; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_661 = _T_85 ? _GEN_644 : _GEN_334; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_662 = _T_85 ? _GEN_645 : regfileWrite_signal_r_dst; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_663 = _T_85 ? _GEN_646 : {{32'd0}, _GEN_336}; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_664 = _T_85 ? _GEN_647 : _GEN_337; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_665 = _T_85 ? _GEN_648 : _GEN_338; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_666 = _T_85 ? _GEN_649 : _GEN_339; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_667 = _T_85 ? _GEN_650 : _GEN_340; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_668 = _T_85 ? _GEN_651 : _GEN_103; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_669 = _T_85 ? _GEN_652 : {{32'd0}, _GEN_104}; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_670 = _T_85 ? _GEN_653 : _GEN_341; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_671 = _T_85 ? _GEN_654 : _GEN_342; // @[ISA.scala 225:44:@1543.6]
    assign _GEN_672 = _T_85 ? _GEN_655 : _GEN_343; // @[ISA.scala 225:44:@1543.6]
    assign _T_31159 = _GEN_486 == 64'h0; // @[ISA_functions.scala 91:81:@21596.14]
    assign _T_31160 = _T_5066 & _T_31159; // @[ISA_functions.scala 91:67:@21597.14]
    assign _T_31171 = _T_110 | _T_128; // @[ISA_functions.scala 251:71:@21604.16]
    assign _T_31176 = _T_31171 | _T_153; // @[ISA_functions.scala 251:120:@21607.16]
    assign _T_31178 = io_fromMemoryPort_loadedData >> 32'h1f; // @[ISA_functions.scala 251:190:@21608.16]
    assign _T_31181 = _T_31178 & 32'h1; // @[ISA_functions.scala 251:212:@21610.16]
    assign _T_31183 = _T_31181 == 32'h0; // @[ISA_functions.scala 251:225:@21611.16]
    assign _T_31184 = _T_31176 & _T_31183; // @[ISA_functions.scala 251:171:@21612.16]
    assign _T_31210 = _T_31183 == 1'h0; // @[ISA_functions.scala 254:179:@21631.18]
    assign _T_31211 = _T_31176 & _T_31210; // @[ISA_functions.scala 254:176:@21632.18]
    assign _T_31217 = 32'hfffff000 | _T_8201; // @[ISA_functions.scala 255:57:@21637.20]
    assign _T_31233 = _T_31176 == 1'h0; // @[ISA_functions.scala 257:28:@21649.20]
    assign _T_31238 = _T_31233 & _T_185; // @[ISA_functions.scala 257:177:@21652.20]
    assign _T_31246 = _T_31238 & _T_31183; // @[ISA_functions.scala 257:226:@21657.20]
    assign _T_31251 = _T_8201 & 32'hfe0; // @[ISA_functions.scala 258:71:@21661.22]
    assign _T_31257 = _T_31251 | _T_2333; // @[ISA_functions.scala 258:87:@21665.22]
    assign _T_31288 = _T_31238 & _T_31210; // @[ISA_functions.scala 260:226:@21686.22]
    assign _T_31302 = 32'hfffff000 | _T_31257; // @[ISA_functions.scala 261:57:@21696.24]
    assign _T_31325 = _T_31233 & _T_219; // @[ISA_functions.scala 263:177:@21712.24]
    assign _T_31330 = _T_31325 & _T_224; // @[ISA_functions.scala 263:227:@21715.24]
    assign _T_31338 = _T_31330 & _T_31183; // @[ISA_functions.scala 263:276:@21720.24]
    assign _GEN_6231 = {{524287'd0}, io_fromMemoryPort_loadedData}; // @[ISA_functions.scala 264:50:@21722.26]
    assign _T_31340 = _GEN_6231 << 19'h4; // @[ISA_functions.scala 264:50:@21722.26]
    assign _T_31341 = _T_31340[31:0]; // @[ISA_functions.scala 264:63:@21723.26]
    assign _T_31343 = _T_31341 & 32'h800; // @[ISA_functions.scala 264:71:@21724.26]
    assign _T_31348 = _T_8201 & 32'h7e0; // @[ISA_functions.scala 264:126:@21727.26]
    assign _T_31349 = _T_31343 | _T_31348; // @[ISA_functions.scala 264:87:@21728.26]
    assign _T_31354 = _T_2330 & 32'h1e; // @[ISA_functions.scala 264:181:@21731.26]
    assign _T_31355 = _T_31349 | _T_31354; // @[ISA_functions.scala 264:143:@21732.26]
    assign _T_31393 = _T_31330 & _T_31210; // @[ISA_functions.scala 266:276:@21757.26]
    assign _T_31413 = 32'hfffff000 | _T_31355; // @[ISA_functions.scala 267:57:@21771.28]
    assign _T_31443 = _T_31325 & _T_265; // @[ISA_functions.scala 269:227:@21791.28]
    assign _T_31453 = _T_31443 & _T_275; // @[ISA_functions.scala 269:277:@21797.28]
    assign _T_31456 = io_fromMemoryPort_loadedData & 32'hfffff000; // @[ISA_functions.scala 270:47:@21800.30]
    assign _T_31498 = _T_31443 & _T_328; // @[ISA_functions.scala 272:277:@21827.30]
    assign _T_31503 = _T_31498 & _T_333; // @[ISA_functions.scala 272:378:@21830.30]
    assign _T_31511 = _T_31503 & _T_31183; // @[ISA_functions.scala 272:428:@21835.30]
    assign _T_31513 = io_fromMemoryPort_loadedData & 32'hff000; // @[ISA_functions.scala 273:49:@21837.32]
    assign _T_31515 = io_fromMemoryPort_loadedData >> 32'h9; // @[ISA_functions.scala 273:85:@21838.32]
    assign _T_31518 = _T_31515 & 32'h800; // @[ISA_functions.scala 273:106:@21840.32]
    assign _T_31519 = _T_31513 | _T_31518; // @[ISA_functions.scala 273:68:@21841.32]
    assign _T_31524 = _T_8201 & 32'h7fe; // @[ISA_functions.scala 273:162:@21844.32]
    assign _T_31525 = _T_31519 | _T_31524; // @[ISA_functions.scala 273:123:@21845.32]
    assign _T_31582 = _T_31503 & _T_31210; // @[ISA_functions.scala 275:428:@21881.32]
    assign _T_31599 = 32'hfff00000 | _T_31525; // @[ISA_functions.scala 276:60:@21893.34]
    assign _GEN_868 = _T_31582 ? _T_31599 : 32'h0; // @[ISA_functions.scala 275:499:@21882.32]
    assign _GEN_869 = _T_31511 ? _T_31525 : _GEN_868; // @[ISA_functions.scala 272:498:@21836.30]
    assign _GEN_870 = _T_31453 ? _T_31456 : _GEN_869; // @[ISA_functions.scala 269:378:@21798.28]
    assign _GEN_871 = _T_31393 ? _T_31413 : _GEN_870; // @[ISA_functions.scala 266:347:@21758.26]
    assign _GEN_872 = _T_31338 ? _T_31355 : _GEN_871; // @[ISA_functions.scala 263:346:@21721.24]
    assign _GEN_873 = _T_31288 ? _T_31302 : _GEN_872; // @[ISA_functions.scala 260:297:@21687.22]
    assign _GEN_874 = _T_31246 ? _T_31257 : _GEN_873; // @[ISA_functions.scala 257:296:@21658.20]
    assign _GEN_875 = _T_31211 ? _T_31217 : _GEN_874; // @[ISA_functions.scala 254:247:@21633.18]
    assign _GEN_876 = _T_31184 ? _T_8201 : _GEN_875; // @[ISA_functions.scala 251:241:@21613.16]
    assign _T_31601 = pcReg_signal_r + _GEN_876; // @[ISA_functions.scala 92:40:@21899.16]
    assign _T_31602 = pcReg_signal_r + _GEN_876; // @[ISA_functions.scala 92:40:@21900.16]
    assign _T_34242 = _T_31160 == 1'h0; // @[ISA_functions.scala 94:28:@23640.16]
    assign _T_36879 = _GEN_486 != 64'h0; // @[ISA_functions.scala 94:164:@25375.16]
    assign _T_36880 = _T_5068 & _T_36879; // @[ISA_functions.scala 94:150:@25376.16]
    assign _T_36881 = _T_34242 & _T_36880; // @[ISA_functions.scala 94:103:@25377.16]
    assign _T_42603 = _T_36880 == 1'h0; // @[ISA_functions.scala 97:106:@29157.18]
    assign _T_42604 = _T_34242 & _T_42603; // @[ISA_functions.scala 97:103:@29158.18]
    assign _T_45241 = _GEN_486 == 64'h1; // @[ISA_functions.scala 97:242:@30893.18]
    assign _T_45242 = _T_5146 & _T_45241; // @[ISA_functions.scala 97:228:@30894.18]
    assign _T_45243 = _T_42604 & _T_45242; // @[ISA_functions.scala 97:181:@30895.18]
    assign _T_53606 = _T_45242 == 1'h0; // @[ISA_functions.scala 100:184:@36413.20]
    assign _T_53607 = _T_42604 & _T_53606; // @[ISA_functions.scala 100:181:@36414.20]
    assign _T_56245 = _T_5148 & _T_31159; // @[ISA_functions.scala 100:306:@38150.20]
    assign _T_56246 = _T_53607 & _T_56245; // @[ISA_functions.scala 100:259:@38151.20]
    assign _T_67250 = _T_56245 == 1'h0; // @[ISA_functions.scala 103:262:@45407.22]
    assign _T_67251 = _T_53607 & _T_67250; // @[ISA_functions.scala 103:259:@45408.22]
    assign _T_69889 = _T_5201 & _T_45241; // @[ISA_functions.scala 103:385:@47144.22]
    assign _T_69890 = _T_67251 & _T_69889; // @[ISA_functions.scala 103:337:@47145.22]
    assign _T_83535 = _T_69889 == 1'h0; // @[ISA_functions.scala 106:340:@56139.24]
    assign _T_83536 = _T_67251 & _T_83535; // @[ISA_functions.scala 106:337:@56140.24]
    assign _T_86174 = _T_5203 & _T_31159; // @[ISA_functions.scala 106:464:@57876.24]
    assign _T_86175 = _T_83536 & _T_86174; // @[ISA_functions.scala 106:416:@57877.24]
    assign _T_86619 = pcReg_signal_r + 32'h4; // @[ISA_functions.scala 110:40:@58184.26]
    assign _T_86620 = pcReg_signal_r + 32'h4; // @[ISA_functions.scala 110:40:@58185.26]
    assign _GEN_1822 = _T_86175 ? _T_31602 : _T_86620; // @[ISA_functions.scala 106:495:@57878.24]
    assign _GEN_1823 = _T_69890 ? _T_31602 : _GEN_1822; // @[ISA_functions.scala 103:416:@47146.22]
    assign _GEN_1824 = _T_56246 ? _T_31602 : _GEN_1823; // @[ISA_functions.scala 100:337:@38152.20]
    assign _GEN_1825 = _T_45243 ? _T_31602 : _GEN_1824; // @[ISA_functions.scala 97:259:@30896.18]
    assign _GEN_1826 = _T_36881 ? _T_31602 : _GEN_1825; // @[ISA_functions.scala 94:181:@25378.16]
    assign _GEN_1827 = _T_31160 ? _T_31602 : _GEN_1826; // @[ISA_functions.scala 91:98:@21598.14]
    assign _GEN_4106 = io_fromMemoryPort_sync ? 3'h4 : _GEN_656; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4107 = io_fromMemoryPort_sync ? _GEN_1827 : _GEN_657; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4108 = io_fromMemoryPort_sync ? 32'h0 : _GEN_658; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4109 = io_fromMemoryPort_sync ? 32'h1 : _GEN_659; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4110 = io_fromMemoryPort_sync ? 32'h1 : _GEN_660; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4111 = io_fromMemoryPort_sync ? _GEN_1827 : _GEN_661; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4112 = io_fromMemoryPort_sync ? regfileWrite_signal_r_dst : _GEN_662; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4113 = io_fromMemoryPort_sync ? {{32'd0}, regfileWrite_signal_r_dstData} : _GEN_663; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4114 = io_fromMemoryPort_sync ? _GEN_1827 : _GEN_664; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4115 = io_fromMemoryPort_sync ? 32'h0 : _GEN_665; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4116 = io_fromMemoryPort_sync ? 32'h1 : _GEN_666; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4117 = io_fromMemoryPort_sync ? 32'h1 : _GEN_667; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4118 = io_fromMemoryPort_sync ? 1'h0 : _GEN_670; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4119 = io_fromMemoryPort_sync ? 1'h1 : _GEN_671; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4120 = io_fromMemoryPort_sync ? 1'h0 : _GEN_672; // @[ISA.scala 251:70:@13955.12]
    assign _GEN_4121 = _T_578 ? _GEN_4106 : _GEN_656; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4122 = _T_578 ? _GEN_4107 : _GEN_657; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4123 = _T_578 ? _GEN_4108 : _GEN_658; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4124 = _T_578 ? _GEN_4109 : _GEN_659; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4125 = _T_578 ? _GEN_4110 : _GEN_660; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4126 = _T_578 ? _GEN_4111 : _GEN_661; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4127 = _T_578 ? _GEN_4112 : _GEN_662; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4128 = _T_578 ? _GEN_4113 : _GEN_663; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4129 = _T_578 ? _GEN_4114 : _GEN_664; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4130 = _T_578 ? _GEN_4115 : _GEN_665; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4131 = _T_578 ? _GEN_4116 : _GEN_666; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4132 = _T_578 ? _GEN_4117 : _GEN_667; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4133 = _T_578 ? _GEN_4118 : _GEN_670; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4134 = _T_578 ? _GEN_4119 : _GEN_671; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4135 = _T_578 ? _GEN_4120 : _GEN_672; // @[ISA.scala 250:92:@13954.10]
    assign _GEN_4136 = _T_337 ? _GEN_4121 : _GEN_656; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4137 = _T_337 ? _GEN_4122 : _GEN_657; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4138 = _T_337 ? _GEN_4123 : _GEN_658; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4139 = _T_337 ? _GEN_4124 : _GEN_659; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4140 = _T_337 ? _GEN_4125 : _GEN_660; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4141 = _T_337 ? _GEN_4126 : _GEN_661; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4142 = _T_337 ? _GEN_4127 : _GEN_662; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4143 = _T_337 ? _GEN_4128 : _GEN_663; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4144 = _T_337 ? _GEN_4129 : _GEN_664; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4145 = _T_337 ? _GEN_4130 : _GEN_665; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4146 = _T_337 ? _GEN_4131 : _GEN_666; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4147 = _T_337 ? _GEN_4132 : _GEN_667; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4148 = _T_337 ? _GEN_4133 : _GEN_670; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4149 = _T_337 ? _GEN_4134 : _GEN_671; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4150 = _T_337 ? _GEN_4135 : _GEN_672; // @[ISA.scala 249:85:@13783.8]
    assign _GEN_4151 = _T_85 ? _GEN_4136 : _GEN_656; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4152 = _T_85 ? _GEN_4137 : _GEN_657; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4153 = _T_85 ? _GEN_4138 : _GEN_658; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4154 = _T_85 ? _GEN_4139 : _GEN_659; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4155 = _T_85 ? _GEN_4140 : _GEN_660; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4156 = _T_85 ? _GEN_4141 : _GEN_661; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4157 = _T_85 ? _GEN_4142 : _GEN_662; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4158 = _T_85 ? _GEN_4143 : _GEN_663; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4159 = _T_85 ? _GEN_4144 : _GEN_664; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4160 = _T_85 ? _GEN_4145 : _GEN_665; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4161 = _T_85 ? _GEN_4146 : _GEN_666; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4162 = _T_85 ? _GEN_4147 : _GEN_667; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4163 = _T_85 ? _GEN_4148 : _GEN_670; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4164 = _T_85 ? _GEN_4149 : _GEN_671; // @[ISA.scala 248:44:@13611.6]
    assign _GEN_4165 = _T_85 ? _GEN_4150 : _GEN_672; // @[ISA.scala 248:44:@13611.6]
    assign _T_223492 = _GEN_441 + _GEN_876; // @[ISA_functions.scala 162:43:@149070.18]
    assign _T_223493 = _GEN_441 + _GEN_876; // @[ISA_functions.scala 162:43:@149071.18]
    assign _T_223500 = _GEN_876 * 32'hffffffff; // @[ISA_functions.scala 165:55:@149080.20]
    assign _T_223501 = _GEN_6225 + _T_223500; // @[ISA_functions.scala 165:43:@149081.20]
    assign _T_223502 = _GEN_6225 + _T_223500; // @[ISA_functions.scala 165:43:@149082.20]
    assign _T_223512 = _GEN_441 & _GEN_876; // @[ISA_functions.scala 168:43:@149094.22]
    assign _T_223526 = _GEN_441 | _GEN_876; // @[ISA_functions.scala 171:43:@149109.24]
    assign _T_223544 = _GEN_441 ^ _GEN_876; // @[ISA_functions.scala 174:43:@149127.26]
    assign _T_223567 = $signed(_GEN_876); // @[ISA_functions.scala 176:237:@149148.26]
    assign _T_223568 = $signed(_T_10673) < $signed(_T_223567); // @[ISA_functions.scala 176:225:@149149.26]
    assign _T_223596 = _T_223568 == 1'h0; // @[ISA_functions.scala 179:206:@149174.28]
    assign _T_223624 = _GEN_441 < _GEN_876; // @[ISA_functions.scala 182:247:@149199.30]
    assign _T_223654 = _T_223624 == 1'h0; // @[ISA_functions.scala 185:237:@149225.32]
    assign _T_223686 = _GEN_876[18:0]; // @[ISA_functions.scala 189:55:@149254.36]
    assign _T_223688 = _T_223686 & 19'h1f; // @[ISA_functions.scala 189:62:@149255.36]
    assign _T_223689 = _GEN_6226 << _T_223688; // @[ISA_functions.scala 189:43:@149256.36]
    assign _T_223690 = _T_223689[31:0]; // @[ISA_functions.scala 189:76:@149257.36]
    assign _T_223726 = _GEN_876 & 32'h1f; // @[ISA_functions.scala 192:67:@149288.38]
    assign _T_223727 = $signed(_T_10673) >>> _T_223726; // @[ISA_functions.scala 192:53:@149289.38]
    assign _T_223728 = $unsigned(_T_223727); // @[ISA_functions.scala 192:82:@149290.38]
    assign _T_223768 = _GEN_441 >> _T_223726; // @[ISA_functions.scala 195:43:@149324.40]
    assign _GEN_4243 = {{32'd0}, _T_223493}; // @[ISA_functions.scala 161:50:@149069.16]
    assign _T_228862 = _T_5012 | _T_5022; // @[ISA_functions.scala 429:45:@152675.16]
    assign _T_228873 = _T_228862 == 1'h0; // @[ISA_functions.scala 432:28:@152683.18]
    assign _T_228876 = _T_5014 | _T_5024; // @[ISA_functions.scala 432:101:@152686.18]
    assign _T_228877 = _T_228873 & _T_228876; // @[ISA_functions.scala 432:76:@152687.18]
    assign _T_228887 = _T_228876 == 1'h0; // @[ISA_functions.scala 435:79:@152699.20]
    assign _T_228888 = _T_228873 & _T_228887; // @[ISA_functions.scala 435:76:@152700.20]
    assign _T_228891 = _T_5016 | _T_5026; // @[ISA_functions.scala 435:152:@152703.20]
    assign _T_228892 = _T_228888 & _T_228891; // @[ISA_functions.scala 435:127:@152704.20]
    assign _T_228908 = _T_228891 == 1'h0; // @[ISA_functions.scala 438:130:@152721.22]
    assign _T_228909 = _T_228888 & _T_228908; // @[ISA_functions.scala 438:127:@152722.22]
    assign _T_228911 = _T_228909 & _T_5018; // @[ISA_functions.scala 438:178:@152724.22]
    assign _T_228931 = _T_5018 == 1'h0; // @[ISA_functions.scala 441:181:@152744.24]
    assign _T_228932 = _T_228909 & _T_228931; // @[ISA_functions.scala 441:178:@152745.24]
    assign _T_228934 = _T_228932 & _T_5020; // @[ISA_functions.scala 441:204:@152747.24]
    assign _GEN_4321 = _T_228934 ? 32'h4 : 32'h0; // @[ISA_functions.scala 441:230:@152748.24]
    assign _GEN_4322 = _T_228911 ? 32'h5 : _GEN_4321; // @[ISA_functions.scala 438:204:@152725.22]
    assign _GEN_4323 = _T_228892 ? 32'h1 : _GEN_4322; // @[ISA_functions.scala 435:178:@152705.20]
    assign _GEN_4324 = _T_228877 ? 32'h2 : _GEN_4323; // @[ISA_functions.scala 432:127:@152688.18]
    assign _GEN_4325 = _T_228862 ? 32'h3 : _GEN_4324; // @[ISA_functions.scala 429:71:@152676.16]
    assign _GEN_4462 = io_fromMemoryPort_sync ? 3'h0 : _GEN_4151; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4463 = io_fromMemoryPort_sync ? _GEN_4243 : {{32'd0}, _GEN_4152}; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4464 = io_fromMemoryPort_sync ? _GEN_473 : _GEN_4153; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4465 = io_fromMemoryPort_sync ? _GEN_4325 : _GEN_4154; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4466 = io_fromMemoryPort_sync ? 32'h2 : _GEN_4155; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4467 = io_fromMemoryPort_sync ? pcReg_signal_r : _GEN_4156; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4468 = io_fromMemoryPort_sync ? regfileWrite_signal_r_dst : _GEN_4157; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4469 = io_fromMemoryPort_sync ? {{32'd0}, regfileWrite_signal_r_dstData} : _GEN_4158; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4470 = io_fromMemoryPort_sync ? _GEN_4243 : {{32'd0}, _GEN_4159}; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4471 = io_fromMemoryPort_sync ? _GEN_473 : _GEN_4160; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4472 = io_fromMemoryPort_sync ? _GEN_4325 : _GEN_4161; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4473 = io_fromMemoryPort_sync ? 32'h2 : _GEN_4162; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4474 = io_fromMemoryPort_sync ? 1'h0 : _GEN_4163; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4475 = io_fromMemoryPort_sync ? 1'h1 : _GEN_4164; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4476 = io_fromMemoryPort_sync ? 1'h0 : _GEN_4165; // @[ISA.scala 275:78:@147185.14]
    assign _GEN_4477 = _T_821 ? _GEN_4462 : _GEN_4151; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4478 = _T_821 ? _GEN_4463 : {{32'd0}, _GEN_4152}; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4479 = _T_821 ? _GEN_4464 : _GEN_4153; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4480 = _T_821 ? _GEN_4465 : _GEN_4154; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4481 = _T_821 ? _GEN_4466 : _GEN_4155; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4482 = _T_821 ? _GEN_4467 : _GEN_4156; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4483 = _T_821 ? _GEN_4468 : _GEN_4157; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4484 = _T_821 ? _GEN_4469 : _GEN_4158; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4485 = _T_821 ? _GEN_4470 : {{32'd0}, _GEN_4159}; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4486 = _T_821 ? _GEN_4471 : _GEN_4160; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4487 = _T_821 ? _GEN_4472 : _GEN_4161; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4488 = _T_821 ? _GEN_4473 : _GEN_4162; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4489 = _T_821 ? _GEN_4474 : _GEN_4163; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4490 = _T_821 ? _GEN_4475 : _GEN_4164; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4491 = _T_821 ? _GEN_4476 : _GEN_4165; // @[ISA.scala 274:100:@147184.12]
    assign _GEN_4492 = _T_580 ? _GEN_4477 : _GEN_4151; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4493 = _T_580 ? _GEN_4478 : {{32'd0}, _GEN_4152}; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4494 = _T_580 ? _GEN_4479 : _GEN_4153; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4495 = _T_580 ? _GEN_4480 : _GEN_4154; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4496 = _T_580 ? _GEN_4481 : _GEN_4155; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4497 = _T_580 ? _GEN_4482 : _GEN_4156; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4498 = _T_580 ? _GEN_4483 : _GEN_4157; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4499 = _T_580 ? _GEN_4484 : _GEN_4158; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4500 = _T_580 ? _GEN_4485 : {{32'd0}, _GEN_4159}; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4501 = _T_580 ? _GEN_4486 : _GEN_4160; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4502 = _T_580 ? _GEN_4487 : _GEN_4161; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4503 = _T_580 ? _GEN_4488 : _GEN_4162; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4504 = _T_580 ? _GEN_4489 : _GEN_4163; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4505 = _T_580 ? _GEN_4490 : _GEN_4164; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4506 = _T_580 ? _GEN_4491 : _GEN_4165; // @[ISA.scala 273:93:@147013.10]
    assign _GEN_4507 = _T_337 ? _GEN_4492 : _GEN_4151; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4508 = _T_337 ? _GEN_4493 : {{32'd0}, _GEN_4152}; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4509 = _T_337 ? _GEN_4494 : _GEN_4153; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4510 = _T_337 ? _GEN_4495 : _GEN_4154; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4511 = _T_337 ? _GEN_4496 : _GEN_4155; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4512 = _T_337 ? _GEN_4497 : _GEN_4156; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4513 = _T_337 ? _GEN_4498 : _GEN_4157; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4514 = _T_337 ? _GEN_4499 : _GEN_4158; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4515 = _T_337 ? _GEN_4500 : {{32'd0}, _GEN_4159}; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4516 = _T_337 ? _GEN_4501 : _GEN_4160; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4517 = _T_337 ? _GEN_4502 : _GEN_4161; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4518 = _T_337 ? _GEN_4503 : _GEN_4162; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4519 = _T_337 ? _GEN_4504 : _GEN_4163; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4520 = _T_337 ? _GEN_4505 : _GEN_4164; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4521 = _T_337 ? _GEN_4506 : _GEN_4165; // @[ISA.scala 272:85:@146841.8]
    assign _GEN_4522 = _T_85 ? _GEN_4507 : _GEN_4151; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4523 = _T_85 ? _GEN_4508 : {{32'd0}, _GEN_4152}; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4524 = _T_85 ? _GEN_4509 : _GEN_4153; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4525 = _T_85 ? _GEN_4510 : _GEN_4154; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4526 = _T_85 ? _GEN_4511 : _GEN_4155; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4527 = _T_85 ? _GEN_4512 : _GEN_4156; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4528 = _T_85 ? _GEN_4513 : _GEN_4157; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4529 = _T_85 ? _GEN_4514 : _GEN_4158; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4530 = _T_85 ? _GEN_4515 : {{32'd0}, _GEN_4159}; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4531 = _T_85 ? _GEN_4516 : _GEN_4160; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4532 = _T_85 ? _GEN_4517 : _GEN_4161; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4533 = _T_85 ? _GEN_4518 : _GEN_4162; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4534 = _T_85 ? _GEN_4519 : _GEN_4163; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4535 = _T_85 ? _GEN_4520 : _GEN_4164; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_4536 = _T_85 ? _GEN_4521 : _GEN_4165; // @[ISA.scala 271:44:@146669.6]
    assign _GEN_6281 = {{32'd0}, _GEN_876}; // @[ISA_functions.scala 165:43:@161117.24]
    assign _GEN_4658 = {{32'd0}, _T_31602}; // @[ISA_functions.scala 161:50:@161706.20]
    assign _GEN_4659 = _T_5755 ? _GEN_6281 : _GEN_4658; // @[ISA_functions.scala 240:67:@160802.18]
    assign _GEN_4751 = io_fromMemoryPort_sync ? 3'h4 : _GEN_4522; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4752 = io_fromMemoryPort_sync ? {{32'd0}, _T_50} : _GEN_4523; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4753 = io_fromMemoryPort_sync ? 32'h0 : _GEN_4524; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4754 = io_fromMemoryPort_sync ? 32'h1 : _GEN_4525; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4755 = io_fromMemoryPort_sync ? 32'h1 : _GEN_4526; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4756 = io_fromMemoryPort_sync ? _T_50 : _GEN_4527; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4757 = io_fromMemoryPort_sync ? _GEN_352 : _GEN_4528; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4758 = io_fromMemoryPort_sync ? _GEN_4659 : _GEN_4529; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4759 = io_fromMemoryPort_sync ? {{32'd0}, _T_50} : _GEN_4530; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4760 = io_fromMemoryPort_sync ? 32'h0 : _GEN_4531; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4761 = io_fromMemoryPort_sync ? 32'h1 : _GEN_4532; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4762 = io_fromMemoryPort_sync ? 32'h1 : _GEN_4533; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4763 = io_fromMemoryPort_sync ? _GEN_352 : _GEN_668; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4764 = io_fromMemoryPort_sync ? _GEN_4659 : _GEN_669; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4765 = io_fromMemoryPort_sync ? 1'h0 : _GEN_4534; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4766 = io_fromMemoryPort_sync ? 1'h1 : _GEN_4535; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4767 = io_fromMemoryPort_sync ? 1'h1 : _GEN_4536; // @[ISA.scala 301:86:@159025.16]
    assign _GEN_4768 = _T_1064 ? _GEN_4751 : _GEN_4522; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4769 = _T_1064 ? _GEN_4752 : _GEN_4523; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4770 = _T_1064 ? _GEN_4753 : _GEN_4524; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4771 = _T_1064 ? _GEN_4754 : _GEN_4525; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4772 = _T_1064 ? _GEN_4755 : _GEN_4526; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4773 = _T_1064 ? _GEN_4756 : _GEN_4527; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4774 = _T_1064 ? _GEN_4757 : _GEN_4528; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4775 = _T_1064 ? _GEN_4758 : _GEN_4529; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4776 = _T_1064 ? _GEN_4759 : _GEN_4530; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4777 = _T_1064 ? _GEN_4760 : _GEN_4531; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4778 = _T_1064 ? _GEN_4761 : _GEN_4532; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4779 = _T_1064 ? _GEN_4762 : _GEN_4533; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4780 = _T_1064 ? _GEN_4763 : _GEN_668; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4781 = _T_1064 ? _GEN_4764 : _GEN_669; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4782 = _T_1064 ? _GEN_4765 : _GEN_4534; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4783 = _T_1064 ? _GEN_4766 : _GEN_4535; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4784 = _T_1064 ? _GEN_4767 : _GEN_4536; // @[ISA.scala 300:108:@159024.14]
    assign _GEN_4785 = _T_823 ? _GEN_4768 : _GEN_4522; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4786 = _T_823 ? _GEN_4769 : _GEN_4523; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4787 = _T_823 ? _GEN_4770 : _GEN_4524; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4788 = _T_823 ? _GEN_4771 : _GEN_4525; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4789 = _T_823 ? _GEN_4772 : _GEN_4526; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4790 = _T_823 ? _GEN_4773 : _GEN_4527; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4791 = _T_823 ? _GEN_4774 : _GEN_4528; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4792 = _T_823 ? _GEN_4775 : _GEN_4529; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4793 = _T_823 ? _GEN_4776 : _GEN_4530; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4794 = _T_823 ? _GEN_4777 : _GEN_4531; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4795 = _T_823 ? _GEN_4778 : _GEN_4532; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4796 = _T_823 ? _GEN_4779 : _GEN_4533; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4797 = _T_823 ? _GEN_4780 : _GEN_668; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4798 = _T_823 ? _GEN_4781 : _GEN_669; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4799 = _T_823 ? _GEN_4782 : _GEN_4534; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4800 = _T_823 ? _GEN_4783 : _GEN_4535; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4801 = _T_823 ? _GEN_4784 : _GEN_4536; // @[ISA.scala 299:101:@158853.12]
    assign _GEN_4802 = _T_580 ? _GEN_4785 : _GEN_4522; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4803 = _T_580 ? _GEN_4786 : _GEN_4523; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4804 = _T_580 ? _GEN_4787 : _GEN_4524; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4805 = _T_580 ? _GEN_4788 : _GEN_4525; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4806 = _T_580 ? _GEN_4789 : _GEN_4526; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4807 = _T_580 ? _GEN_4790 : _GEN_4527; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4808 = _T_580 ? _GEN_4791 : _GEN_4528; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4809 = _T_580 ? _GEN_4792 : _GEN_4529; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4810 = _T_580 ? _GEN_4793 : _GEN_4530; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4811 = _T_580 ? _GEN_4794 : _GEN_4531; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4812 = _T_580 ? _GEN_4795 : _GEN_4532; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4813 = _T_580 ? _GEN_4796 : _GEN_4533; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4814 = _T_580 ? _GEN_4797 : _GEN_668; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4815 = _T_580 ? _GEN_4798 : _GEN_669; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4816 = _T_580 ? _GEN_4799 : _GEN_4534; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4817 = _T_580 ? _GEN_4800 : _GEN_4535; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4818 = _T_580 ? _GEN_4801 : _GEN_4536; // @[ISA.scala 298:93:@158681.10]
    assign _GEN_4819 = _T_337 ? _GEN_4802 : _GEN_4522; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4820 = _T_337 ? _GEN_4803 : _GEN_4523; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4821 = _T_337 ? _GEN_4804 : _GEN_4524; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4822 = _T_337 ? _GEN_4805 : _GEN_4525; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4823 = _T_337 ? _GEN_4806 : _GEN_4526; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4824 = _T_337 ? _GEN_4807 : _GEN_4527; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4825 = _T_337 ? _GEN_4808 : _GEN_4528; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4826 = _T_337 ? _GEN_4809 : _GEN_4529; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4827 = _T_337 ? _GEN_4810 : _GEN_4530; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4828 = _T_337 ? _GEN_4811 : _GEN_4531; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4829 = _T_337 ? _GEN_4812 : _GEN_4532; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4830 = _T_337 ? _GEN_4813 : _GEN_4533; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4831 = _T_337 ? _GEN_4814 : _GEN_668; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4832 = _T_337 ? _GEN_4815 : _GEN_669; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4833 = _T_337 ? _GEN_4816 : _GEN_4534; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4834 = _T_337 ? _GEN_4817 : _GEN_4535; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4835 = _T_337 ? _GEN_4818 : _GEN_4536; // @[ISA.scala 297:85:@158509.8]
    assign _GEN_4836 = _T_85 ? _GEN_4819 : _GEN_4522; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4837 = _T_85 ? _GEN_4820 : _GEN_4523; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4838 = _T_85 ? _GEN_4821 : _GEN_4524; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4839 = _T_85 ? _GEN_4822 : _GEN_4525; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4840 = _T_85 ? _GEN_4823 : _GEN_4526; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4841 = _T_85 ? _GEN_4824 : _GEN_4527; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4842 = _T_85 ? _GEN_4825 : _GEN_4528; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4843 = _T_85 ? _GEN_4826 : _GEN_4529; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4844 = _T_85 ? _GEN_4827 : _GEN_4530; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4845 = _T_85 ? _GEN_4828 : _GEN_4531; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4846 = _T_85 ? _GEN_4829 : _GEN_4532; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4847 = _T_85 ? _GEN_4830 : _GEN_4533; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4848 = _T_85 ? _GEN_4831 : _GEN_668; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4849 = _T_85 ? _GEN_4832 : _GEN_669; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4850 = _T_85 ? _GEN_4833 : _GEN_4534; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4851 = _T_85 ? _GEN_4834 : _GEN_4535; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4852 = _T_85 ? _GEN_4835 : _GEN_4536; // @[ISA.scala 296:44:@158337.6]
    assign _GEN_4922 = io_fromMemoryPort_sync ? 3'h4 : _GEN_4836; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4923 = io_fromMemoryPort_sync ? {{32'd0}, _T_31602} : _GEN_4837; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4924 = io_fromMemoryPort_sync ? 32'h0 : _GEN_4838; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4925 = io_fromMemoryPort_sync ? 32'h1 : _GEN_4839; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4926 = io_fromMemoryPort_sync ? 32'h1 : _GEN_4840; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4927 = io_fromMemoryPort_sync ? _T_31602 : _GEN_4841; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4928 = io_fromMemoryPort_sync ? _GEN_352 : _GEN_4842; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4929 = io_fromMemoryPort_sync ? {{32'd0}, _T_50} : _GEN_4843; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4930 = io_fromMemoryPort_sync ? {{32'd0}, _T_31602} : _GEN_4844; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4931 = io_fromMemoryPort_sync ? 32'h0 : _GEN_4845; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4932 = io_fromMemoryPort_sync ? 32'h1 : _GEN_4846; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4933 = io_fromMemoryPort_sync ? 32'h1 : _GEN_4847; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4934 = io_fromMemoryPort_sync ? _GEN_352 : _GEN_4848; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4935 = io_fromMemoryPort_sync ? {{32'd0}, _T_50} : _GEN_4849; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4936 = io_fromMemoryPort_sync ? 1'h0 : _GEN_4850; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4937 = io_fromMemoryPort_sync ? 1'h1 : _GEN_4851; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4938 = io_fromMemoryPort_sync ? 1'h1 : _GEN_4852; // @[ISA.scala 331:94:@165852.18]
    assign _GEN_4939 = _T_1307 ? _GEN_4922 : _GEN_4836; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4940 = _T_1307 ? _GEN_4923 : _GEN_4837; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4941 = _T_1307 ? _GEN_4924 : _GEN_4838; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4942 = _T_1307 ? _GEN_4925 : _GEN_4839; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4943 = _T_1307 ? _GEN_4926 : _GEN_4840; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4944 = _T_1307 ? _GEN_4927 : _GEN_4841; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4945 = _T_1307 ? _GEN_4928 : _GEN_4842; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4946 = _T_1307 ? _GEN_4929 : _GEN_4843; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4947 = _T_1307 ? _GEN_4930 : _GEN_4844; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4948 = _T_1307 ? _GEN_4931 : _GEN_4845; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4949 = _T_1307 ? _GEN_4932 : _GEN_4846; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4950 = _T_1307 ? _GEN_4933 : _GEN_4847; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4951 = _T_1307 ? _GEN_4934 : _GEN_4848; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4952 = _T_1307 ? _GEN_4935 : _GEN_4849; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4953 = _T_1307 ? _GEN_4936 : _GEN_4850; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4954 = _T_1307 ? _GEN_4937 : _GEN_4851; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4955 = _T_1307 ? _GEN_4938 : _GEN_4852; // @[ISA.scala 330:116:@165851.16]
    assign _GEN_4956 = _T_1066 ? _GEN_4939 : _GEN_4836; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4957 = _T_1066 ? _GEN_4940 : _GEN_4837; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4958 = _T_1066 ? _GEN_4941 : _GEN_4838; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4959 = _T_1066 ? _GEN_4942 : _GEN_4839; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4960 = _T_1066 ? _GEN_4943 : _GEN_4840; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4961 = _T_1066 ? _GEN_4944 : _GEN_4841; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4962 = _T_1066 ? _GEN_4945 : _GEN_4842; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4963 = _T_1066 ? _GEN_4946 : _GEN_4843; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4964 = _T_1066 ? _GEN_4947 : _GEN_4844; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4965 = _T_1066 ? _GEN_4948 : _GEN_4845; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4966 = _T_1066 ? _GEN_4949 : _GEN_4846; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4967 = _T_1066 ? _GEN_4950 : _GEN_4847; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4968 = _T_1066 ? _GEN_4951 : _GEN_4848; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4969 = _T_1066 ? _GEN_4952 : _GEN_4849; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4970 = _T_1066 ? _GEN_4953 : _GEN_4850; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4971 = _T_1066 ? _GEN_4954 : _GEN_4851; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4972 = _T_1066 ? _GEN_4955 : _GEN_4852; // @[ISA.scala 329:109:@165680.14]
    assign _GEN_4973 = _T_823 ? _GEN_4956 : _GEN_4836; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4974 = _T_823 ? _GEN_4957 : _GEN_4837; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4975 = _T_823 ? _GEN_4958 : _GEN_4838; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4976 = _T_823 ? _GEN_4959 : _GEN_4839; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4977 = _T_823 ? _GEN_4960 : _GEN_4840; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4978 = _T_823 ? _GEN_4961 : _GEN_4841; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4979 = _T_823 ? _GEN_4962 : _GEN_4842; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4980 = _T_823 ? _GEN_4963 : _GEN_4843; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4981 = _T_823 ? _GEN_4964 : _GEN_4844; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4982 = _T_823 ? _GEN_4965 : _GEN_4845; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4983 = _T_823 ? _GEN_4966 : _GEN_4846; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4984 = _T_823 ? _GEN_4967 : _GEN_4847; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4985 = _T_823 ? _GEN_4968 : _GEN_4848; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4986 = _T_823 ? _GEN_4969 : _GEN_4849; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4987 = _T_823 ? _GEN_4970 : _GEN_4850; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4988 = _T_823 ? _GEN_4971 : _GEN_4851; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4989 = _T_823 ? _GEN_4972 : _GEN_4852; // @[ISA.scala 328:101:@165508.12]
    assign _GEN_4990 = _T_580 ? _GEN_4973 : _GEN_4836; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_4991 = _T_580 ? _GEN_4974 : _GEN_4837; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_4992 = _T_580 ? _GEN_4975 : _GEN_4838; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_4993 = _T_580 ? _GEN_4976 : _GEN_4839; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_4994 = _T_580 ? _GEN_4977 : _GEN_4840; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_4995 = _T_580 ? _GEN_4978 : _GEN_4841; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_4996 = _T_580 ? _GEN_4979 : _GEN_4842; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_4997 = _T_580 ? _GEN_4980 : _GEN_4843; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_4998 = _T_580 ? _GEN_4981 : _GEN_4844; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_4999 = _T_580 ? _GEN_4982 : _GEN_4845; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_5000 = _T_580 ? _GEN_4983 : _GEN_4846; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_5001 = _T_580 ? _GEN_4984 : _GEN_4847; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_5002 = _T_580 ? _GEN_4985 : _GEN_4848; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_5003 = _T_580 ? _GEN_4986 : _GEN_4849; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_5004 = _T_580 ? _GEN_4987 : _GEN_4850; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_5005 = _T_580 ? _GEN_4988 : _GEN_4851; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_5006 = _T_580 ? _GEN_4989 : _GEN_4852; // @[ISA.scala 327:93:@165336.10]
    assign _GEN_5007 = _T_337 ? _GEN_4990 : _GEN_4836; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5008 = _T_337 ? _GEN_4991 : _GEN_4837; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5009 = _T_337 ? _GEN_4992 : _GEN_4838; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5010 = _T_337 ? _GEN_4993 : _GEN_4839; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5011 = _T_337 ? _GEN_4994 : _GEN_4840; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5012 = _T_337 ? _GEN_4995 : _GEN_4841; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5013 = _T_337 ? _GEN_4996 : _GEN_4842; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5014 = _T_337 ? _GEN_4997 : _GEN_4843; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5015 = _T_337 ? _GEN_4998 : _GEN_4844; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5016 = _T_337 ? _GEN_4999 : _GEN_4845; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5017 = _T_337 ? _GEN_5000 : _GEN_4846; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5018 = _T_337 ? _GEN_5001 : _GEN_4847; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5019 = _T_337 ? _GEN_5002 : _GEN_4848; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5020 = _T_337 ? _GEN_5003 : _GEN_4849; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5021 = _T_337 ? _GEN_5004 : _GEN_4850; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5022 = _T_337 ? _GEN_5005 : _GEN_4851; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5023 = _T_337 ? _GEN_5006 : _GEN_4852; // @[ISA.scala 326:85:@165164.8]
    assign _GEN_5024 = _T_85 ? _GEN_5007 : _GEN_4836; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5025 = _T_85 ? _GEN_5008 : _GEN_4837; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5026 = _T_85 ? _GEN_5009 : _GEN_4838; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5027 = _T_85 ? _GEN_5010 : _GEN_4839; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5028 = _T_85 ? _GEN_5011 : _GEN_4840; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5029 = _T_85 ? _GEN_5012 : _GEN_4841; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5030 = _T_85 ? _GEN_5013 : _GEN_4842; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5031 = _T_85 ? _GEN_5014 : _GEN_4843; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5032 = _T_85 ? _GEN_5015 : _GEN_4844; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5033 = _T_85 ? _GEN_5016 : _GEN_4845; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5034 = _T_85 ? _GEN_5017 : _GEN_4846; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5035 = _T_85 ? _GEN_5018 : _GEN_4847; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5036 = _T_85 ? _GEN_5019 : _GEN_4848; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5037 = _T_85 ? _GEN_5020 : _GEN_4849; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5038 = _T_85 ? _GEN_5021 : _GEN_4850; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5039 = _T_85 ? _GEN_5022 : _GEN_4851; // @[ISA.scala 325:44:@164992.6]
    assign _GEN_5040 = _T_85 ? _GEN_5023 : _GEN_4852; // @[ISA.scala 325:44:@164992.6]
    assign _T_257102 = _T_10672 & _T_223568; // @[ISA_functions.scala 176:203:@172339.32]
    assign _T_257130 = _T_10672 & _T_223596; // @[ISA_functions.scala 179:203:@172364.34]
    assign _T_257158 = _T_10730 & _T_223624; // @[ISA_functions.scala 182:234:@172389.36]
    assign _T_257188 = _T_10730 & _T_223654; // @[ISA_functions.scala 185:234:@172415.38]
    assign _GEN_5189 = _T_10872 ? _T_223768 : _GEN_474; // @[ISA_functions.scala 194:325:@172511.44]
    assign _GEN_5190 = _T_10830 ? _T_223728 : _GEN_5189; // @[ISA_functions.scala 191:295:@172475.42]
    assign _GEN_5191 = _T_10792 ? _T_223690 : _GEN_5190; // @[ISA_functions.scala 188:265:@172442.40]
    assign _GEN_5192 = _T_257188 ? 32'h0 : _GEN_5191; // @[ISA_functions.scala 185:261:@172416.38]
    assign _GEN_5193 = _T_257158 ? 32'h1 : _GEN_5192; // @[ISA_functions.scala 182:260:@172390.36]
    assign _GEN_5194 = _T_257130 ? 32'h0 : _GEN_5193; // @[ISA_functions.scala 179:248:@172365.34]
    assign _GEN_5195 = _T_257102 ? 32'h1 : _GEN_5194; // @[ISA_functions.scala 176:247:@172340.32]
    assign _GEN_5196 = _T_10650 ? _T_223544 : _GEN_5195; // @[ISA_functions.scala 173:174:@172315.30]
    assign _GEN_5197 = _T_10632 ? _T_223526 : _GEN_5196; // @[ISA_functions.scala 170:144:@172297.28]
    assign _GEN_5198 = _T_10618 ? _T_223512 : _GEN_5197; // @[ISA_functions.scala 167:115:@172282.26]
    assign _GEN_5199 = _T_10605 ? _T_223502 : {{32'd0}, _GEN_5198}; // @[ISA_functions.scala 164:85:@172268.24]
    assign _GEN_5200 = _T_10598 ? {{32'd0}, _T_223493} : _GEN_5199; // @[ISA_functions.scala 161:50:@172258.22]
    assign _GEN_5313 = io_fromMemoryPort_sync ? 3'h4 : _GEN_5024; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5314 = io_fromMemoryPort_sync ? {{32'd0}, _T_50} : _GEN_5025; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5315 = io_fromMemoryPort_sync ? 32'h0 : _GEN_5026; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5316 = io_fromMemoryPort_sync ? 32'h1 : _GEN_5027; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5317 = io_fromMemoryPort_sync ? 32'h1 : _GEN_5028; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5318 = io_fromMemoryPort_sync ? _T_50 : _GEN_5029; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5319 = io_fromMemoryPort_sync ? _GEN_352 : _GEN_5030; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5320 = io_fromMemoryPort_sync ? _GEN_5200 : _GEN_5031; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5321 = io_fromMemoryPort_sync ? {{32'd0}, _T_50} : _GEN_5032; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5322 = io_fromMemoryPort_sync ? 32'h0 : _GEN_5033; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5323 = io_fromMemoryPort_sync ? 32'h1 : _GEN_5034; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5324 = io_fromMemoryPort_sync ? 32'h1 : _GEN_5035; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5325 = io_fromMemoryPort_sync ? _GEN_352 : _GEN_5036; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5326 = io_fromMemoryPort_sync ? _GEN_5200 : _GEN_5037; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5327 = io_fromMemoryPort_sync ? 1'h0 : _GEN_5038; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5328 = io_fromMemoryPort_sync ? 1'h1 : _GEN_5039; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5329 = io_fromMemoryPort_sync ? 1'h1 : _GEN_5040; // @[ISA.scala 363:102:@167880.20]
    assign _GEN_5330 = _T_1550 ? _GEN_5313 : _GEN_5024; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5331 = _T_1550 ? _GEN_5314 : _GEN_5025; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5332 = _T_1550 ? _GEN_5315 : _GEN_5026; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5333 = _T_1550 ? _GEN_5316 : _GEN_5027; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5334 = _T_1550 ? _GEN_5317 : _GEN_5028; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5335 = _T_1550 ? _GEN_5318 : _GEN_5029; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5336 = _T_1550 ? _GEN_5319 : _GEN_5030; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5337 = _T_1550 ? _GEN_5320 : _GEN_5031; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5338 = _T_1550 ? _GEN_5321 : _GEN_5032; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5339 = _T_1550 ? _GEN_5322 : _GEN_5033; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5340 = _T_1550 ? _GEN_5323 : _GEN_5034; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5341 = _T_1550 ? _GEN_5324 : _GEN_5035; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5342 = _T_1550 ? _GEN_5325 : _GEN_5036; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5343 = _T_1550 ? _GEN_5326 : _GEN_5037; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5344 = _T_1550 ? _GEN_5327 : _GEN_5038; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5345 = _T_1550 ? _GEN_5328 : _GEN_5039; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5346 = _T_1550 ? _GEN_5329 : _GEN_5040; // @[ISA.scala 362:126:@167879.18]
    assign _GEN_5347 = _T_1309 ? _GEN_5330 : _GEN_5024; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5348 = _T_1309 ? _GEN_5331 : _GEN_5025; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5349 = _T_1309 ? _GEN_5332 : _GEN_5026; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5350 = _T_1309 ? _GEN_5333 : _GEN_5027; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5351 = _T_1309 ? _GEN_5334 : _GEN_5028; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5352 = _T_1309 ? _GEN_5335 : _GEN_5029; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5353 = _T_1309 ? _GEN_5336 : _GEN_5030; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5354 = _T_1309 ? _GEN_5337 : _GEN_5031; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5355 = _T_1309 ? _GEN_5338 : _GEN_5032; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5356 = _T_1309 ? _GEN_5339 : _GEN_5033; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5357 = _T_1309 ? _GEN_5340 : _GEN_5034; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5358 = _T_1309 ? _GEN_5341 : _GEN_5035; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5359 = _T_1309 ? _GEN_5342 : _GEN_5036; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5360 = _T_1309 ? _GEN_5343 : _GEN_5037; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5361 = _T_1309 ? _GEN_5344 : _GEN_5038; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5362 = _T_1309 ? _GEN_5345 : _GEN_5039; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5363 = _T_1309 ? _GEN_5346 : _GEN_5040; // @[ISA.scala 361:117:@167708.16]
    assign _GEN_5364 = _T_1066 ? _GEN_5347 : _GEN_5024; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5365 = _T_1066 ? _GEN_5348 : _GEN_5025; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5366 = _T_1066 ? _GEN_5349 : _GEN_5026; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5367 = _T_1066 ? _GEN_5350 : _GEN_5027; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5368 = _T_1066 ? _GEN_5351 : _GEN_5028; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5369 = _T_1066 ? _GEN_5352 : _GEN_5029; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5370 = _T_1066 ? _GEN_5353 : _GEN_5030; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5371 = _T_1066 ? _GEN_5354 : _GEN_5031; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5372 = _T_1066 ? _GEN_5355 : _GEN_5032; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5373 = _T_1066 ? _GEN_5356 : _GEN_5033; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5374 = _T_1066 ? _GEN_5357 : _GEN_5034; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5375 = _T_1066 ? _GEN_5358 : _GEN_5035; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5376 = _T_1066 ? _GEN_5359 : _GEN_5036; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5377 = _T_1066 ? _GEN_5360 : _GEN_5037; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5378 = _T_1066 ? _GEN_5361 : _GEN_5038; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5379 = _T_1066 ? _GEN_5362 : _GEN_5039; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5380 = _T_1066 ? _GEN_5363 : _GEN_5040; // @[ISA.scala 360:109:@167536.14]
    assign _GEN_5381 = _T_823 ? _GEN_5364 : _GEN_5024; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5382 = _T_823 ? _GEN_5365 : _GEN_5025; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5383 = _T_823 ? _GEN_5366 : _GEN_5026; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5384 = _T_823 ? _GEN_5367 : _GEN_5027; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5385 = _T_823 ? _GEN_5368 : _GEN_5028; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5386 = _T_823 ? _GEN_5369 : _GEN_5029; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5387 = _T_823 ? _GEN_5370 : _GEN_5030; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5388 = _T_823 ? _GEN_5371 : _GEN_5031; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5389 = _T_823 ? _GEN_5372 : _GEN_5032; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5390 = _T_823 ? _GEN_5373 : _GEN_5033; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5391 = _T_823 ? _GEN_5374 : _GEN_5034; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5392 = _T_823 ? _GEN_5375 : _GEN_5035; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5393 = _T_823 ? _GEN_5376 : _GEN_5036; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5394 = _T_823 ? _GEN_5377 : _GEN_5037; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5395 = _T_823 ? _GEN_5378 : _GEN_5038; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5396 = _T_823 ? _GEN_5379 : _GEN_5039; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5397 = _T_823 ? _GEN_5380 : _GEN_5040; // @[ISA.scala 359:101:@167364.12]
    assign _GEN_5398 = _T_580 ? _GEN_5381 : _GEN_5024; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5399 = _T_580 ? _GEN_5382 : _GEN_5025; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5400 = _T_580 ? _GEN_5383 : _GEN_5026; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5401 = _T_580 ? _GEN_5384 : _GEN_5027; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5402 = _T_580 ? _GEN_5385 : _GEN_5028; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5403 = _T_580 ? _GEN_5386 : _GEN_5029; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5404 = _T_580 ? _GEN_5387 : _GEN_5030; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5405 = _T_580 ? _GEN_5388 : _GEN_5031; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5406 = _T_580 ? _GEN_5389 : _GEN_5032; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5407 = _T_580 ? _GEN_5390 : _GEN_5033; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5408 = _T_580 ? _GEN_5391 : _GEN_5034; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5409 = _T_580 ? _GEN_5392 : _GEN_5035; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5410 = _T_580 ? _GEN_5393 : _GEN_5036; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5411 = _T_580 ? _GEN_5394 : _GEN_5037; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5412 = _T_580 ? _GEN_5395 : _GEN_5038; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5413 = _T_580 ? _GEN_5396 : _GEN_5039; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5414 = _T_580 ? _GEN_5397 : _GEN_5040; // @[ISA.scala 358:93:@167192.10]
    assign _GEN_5415 = _T_337 ? _GEN_5398 : _GEN_5024; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5416 = _T_337 ? _GEN_5399 : _GEN_5025; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5417 = _T_337 ? _GEN_5400 : _GEN_5026; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5418 = _T_337 ? _GEN_5401 : _GEN_5027; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5419 = _T_337 ? _GEN_5402 : _GEN_5028; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5420 = _T_337 ? _GEN_5403 : _GEN_5029; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5421 = _T_337 ? _GEN_5404 : _GEN_5030; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5422 = _T_337 ? _GEN_5405 : _GEN_5031; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5423 = _T_337 ? _GEN_5406 : _GEN_5032; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5424 = _T_337 ? _GEN_5407 : _GEN_5033; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5425 = _T_337 ? _GEN_5408 : _GEN_5034; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5426 = _T_337 ? _GEN_5409 : _GEN_5035; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5427 = _T_337 ? _GEN_5410 : _GEN_5036; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5428 = _T_337 ? _GEN_5411 : _GEN_5037; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5429 = _T_337 ? _GEN_5412 : _GEN_5038; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5430 = _T_337 ? _GEN_5413 : _GEN_5039; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5431 = _T_337 ? _GEN_5414 : _GEN_5040; // @[ISA.scala 357:85:@167020.8]
    assign _GEN_5432 = _T_85 ? _GEN_5415 : _GEN_5024; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5433 = _T_85 ? _GEN_5416 : _GEN_5025; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5434 = _T_85 ? _GEN_5417 : _GEN_5026; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5435 = _T_85 ? _GEN_5418 : _GEN_5027; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5436 = _T_85 ? _GEN_5419 : _GEN_5028; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5437 = _T_85 ? _GEN_5420 : _GEN_5029; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5438 = _T_85 ? _GEN_5421 : _GEN_5030; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5439 = _T_85 ? _GEN_5422 : _GEN_5031; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5440 = _T_85 ? _GEN_5423 : _GEN_5032; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5441 = _T_85 ? _GEN_5424 : _GEN_5033; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5442 = _T_85 ? _GEN_5425 : _GEN_5034; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5443 = _T_85 ? _GEN_5426 : _GEN_5035; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5444 = _T_85 ? _GEN_5427 : _GEN_5036; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5445 = _T_85 ? _GEN_5428 : _GEN_5037; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5446 = _T_85 ? _GEN_5429 : _GEN_5038; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5447 = _T_85 ? _GEN_5430 : _GEN_5039; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5448 = _T_85 ? _GEN_5431 : _GEN_5040; // @[ISA.scala 356:44:@166848.6]
    assign _GEN_5714 = io_fromMemoryPort_sync ? 3'h2 : _GEN_5432; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5715 = io_fromMemoryPort_sync ? _GEN_4243 : _GEN_5433; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5716 = io_fromMemoryPort_sync ? 32'h0 : _GEN_5434; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5717 = io_fromMemoryPort_sync ? _GEN_4325 : _GEN_5435; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5718 = io_fromMemoryPort_sync ? 32'h1 : _GEN_5436; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5719 = io_fromMemoryPort_sync ? pcReg_signal_r : _GEN_5437; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5720 = io_fromMemoryPort_sync ? _GEN_352 : _GEN_5438; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5721 = io_fromMemoryPort_sync ? {{32'd0}, regfileWrite_signal_r_dstData} : _GEN_5439; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5722 = io_fromMemoryPort_sync ? _GEN_4243 : _GEN_5440; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5723 = io_fromMemoryPort_sync ? 32'h0 : _GEN_5441; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5724 = io_fromMemoryPort_sync ? _GEN_4325 : _GEN_5442; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5725 = io_fromMemoryPort_sync ? 32'h1 : _GEN_5443; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5726 = io_fromMemoryPort_sync ? 1'h0 : _GEN_5446; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5727 = io_fromMemoryPort_sync ? 1'h1 : _GEN_5447; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5728 = io_fromMemoryPort_sync ? 1'h0 : _GEN_5448; // @[ISA.scala 397:110:@178443.22]
    assign _GEN_5729 = _T_1793 ? _GEN_5714 : _GEN_5432; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5730 = _T_1793 ? _GEN_5715 : _GEN_5433; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5731 = _T_1793 ? _GEN_5716 : _GEN_5434; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5732 = _T_1793 ? _GEN_5717 : _GEN_5435; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5733 = _T_1793 ? _GEN_5718 : _GEN_5436; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5734 = _T_1793 ? _GEN_5719 : _GEN_5437; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5735 = _T_1793 ? _GEN_5720 : _GEN_5438; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5736 = _T_1793 ? _GEN_5721 : _GEN_5439; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5737 = _T_1793 ? _GEN_5722 : _GEN_5440; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5738 = _T_1793 ? _GEN_5723 : _GEN_5441; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5739 = _T_1793 ? _GEN_5724 : _GEN_5442; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5740 = _T_1793 ? _GEN_5725 : _GEN_5443; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5741 = _T_1793 ? _GEN_5726 : _GEN_5446; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5742 = _T_1793 ? _GEN_5727 : _GEN_5447; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5743 = _T_1793 ? _GEN_5728 : _GEN_5448; // @[ISA.scala 396:134:@178442.20]
    assign _GEN_5744 = _T_1552 ? _GEN_5729 : _GEN_5432; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5745 = _T_1552 ? _GEN_5730 : _GEN_5433; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5746 = _T_1552 ? _GEN_5731 : _GEN_5434; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5747 = _T_1552 ? _GEN_5732 : _GEN_5435; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5748 = _T_1552 ? _GEN_5733 : _GEN_5436; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5749 = _T_1552 ? _GEN_5734 : _GEN_5437; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5750 = _T_1552 ? _GEN_5735 : _GEN_5438; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5751 = _T_1552 ? _GEN_5736 : _GEN_5439; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5752 = _T_1552 ? _GEN_5737 : _GEN_5440; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5753 = _T_1552 ? _GEN_5738 : _GEN_5441; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5754 = _T_1552 ? _GEN_5739 : _GEN_5442; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5755 = _T_1552 ? _GEN_5740 : _GEN_5443; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5756 = _T_1552 ? _GEN_5741 : _GEN_5446; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5757 = _T_1552 ? _GEN_5742 : _GEN_5447; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5758 = _T_1552 ? _GEN_5743 : _GEN_5448; // @[ISA.scala 395:127:@178271.18]
    assign _GEN_5759 = _T_1309 ? _GEN_5744 : _GEN_5432; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5760 = _T_1309 ? _GEN_5745 : _GEN_5433; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5761 = _T_1309 ? _GEN_5746 : _GEN_5434; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5762 = _T_1309 ? _GEN_5747 : _GEN_5435; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5763 = _T_1309 ? _GEN_5748 : _GEN_5436; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5764 = _T_1309 ? _GEN_5749 : _GEN_5437; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5765 = _T_1309 ? _GEN_5750 : _GEN_5438; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5766 = _T_1309 ? _GEN_5751 : _GEN_5439; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5767 = _T_1309 ? _GEN_5752 : _GEN_5440; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5768 = _T_1309 ? _GEN_5753 : _GEN_5441; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5769 = _T_1309 ? _GEN_5754 : _GEN_5442; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5770 = _T_1309 ? _GEN_5755 : _GEN_5443; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5771 = _T_1309 ? _GEN_5756 : _GEN_5446; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5772 = _T_1309 ? _GEN_5757 : _GEN_5447; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5773 = _T_1309 ? _GEN_5758 : _GEN_5448; // @[ISA.scala 394:117:@178099.16]
    assign _GEN_5774 = _T_1066 ? _GEN_5759 : _GEN_5432; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5775 = _T_1066 ? _GEN_5760 : _GEN_5433; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5776 = _T_1066 ? _GEN_5761 : _GEN_5434; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5777 = _T_1066 ? _GEN_5762 : _GEN_5435; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5778 = _T_1066 ? _GEN_5763 : _GEN_5436; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5779 = _T_1066 ? _GEN_5764 : _GEN_5437; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5780 = _T_1066 ? _GEN_5765 : _GEN_5438; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5781 = _T_1066 ? _GEN_5766 : _GEN_5439; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5782 = _T_1066 ? _GEN_5767 : _GEN_5440; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5783 = _T_1066 ? _GEN_5768 : _GEN_5441; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5784 = _T_1066 ? _GEN_5769 : _GEN_5442; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5785 = _T_1066 ? _GEN_5770 : _GEN_5443; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5786 = _T_1066 ? _GEN_5771 : _GEN_5446; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5787 = _T_1066 ? _GEN_5772 : _GEN_5447; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5788 = _T_1066 ? _GEN_5773 : _GEN_5448; // @[ISA.scala 393:109:@177927.14]
    assign _GEN_5789 = _T_823 ? _GEN_5774 : _GEN_5432; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5790 = _T_823 ? _GEN_5775 : _GEN_5433; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5791 = _T_823 ? _GEN_5776 : _GEN_5434; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5792 = _T_823 ? _GEN_5777 : _GEN_5435; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5793 = _T_823 ? _GEN_5778 : _GEN_5436; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5794 = _T_823 ? _GEN_5779 : _GEN_5437; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5795 = _T_823 ? _GEN_5780 : _GEN_5438; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5796 = _T_823 ? _GEN_5781 : _GEN_5439; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5797 = _T_823 ? _GEN_5782 : _GEN_5440; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5798 = _T_823 ? _GEN_5783 : _GEN_5441; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5799 = _T_823 ? _GEN_5784 : _GEN_5442; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5800 = _T_823 ? _GEN_5785 : _GEN_5443; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5801 = _T_823 ? _GEN_5786 : _GEN_5446; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5802 = _T_823 ? _GEN_5787 : _GEN_5447; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5803 = _T_823 ? _GEN_5788 : _GEN_5448; // @[ISA.scala 392:101:@177755.12]
    assign _GEN_5804 = _T_580 ? _GEN_5789 : _GEN_5432; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5805 = _T_580 ? _GEN_5790 : _GEN_5433; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5806 = _T_580 ? _GEN_5791 : _GEN_5434; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5807 = _T_580 ? _GEN_5792 : _GEN_5435; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5808 = _T_580 ? _GEN_5793 : _GEN_5436; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5809 = _T_580 ? _GEN_5794 : _GEN_5437; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5810 = _T_580 ? _GEN_5795 : _GEN_5438; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5811 = _T_580 ? _GEN_5796 : _GEN_5439; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5812 = _T_580 ? _GEN_5797 : _GEN_5440; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5813 = _T_580 ? _GEN_5798 : _GEN_5441; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5814 = _T_580 ? _GEN_5799 : _GEN_5442; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5815 = _T_580 ? _GEN_5800 : _GEN_5443; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5816 = _T_580 ? _GEN_5801 : _GEN_5446; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5817 = _T_580 ? _GEN_5802 : _GEN_5447; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5818 = _T_580 ? _GEN_5803 : _GEN_5448; // @[ISA.scala 391:93:@177583.10]
    assign _GEN_5819 = _T_337 ? _GEN_5804 : _GEN_5432; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5820 = _T_337 ? _GEN_5805 : _GEN_5433; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5821 = _T_337 ? _GEN_5806 : _GEN_5434; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5822 = _T_337 ? _GEN_5807 : _GEN_5435; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5823 = _T_337 ? _GEN_5808 : _GEN_5436; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5824 = _T_337 ? _GEN_5809 : _GEN_5437; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5825 = _T_337 ? _GEN_5810 : _GEN_5438; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5826 = _T_337 ? _GEN_5811 : _GEN_5439; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5827 = _T_337 ? _GEN_5812 : _GEN_5440; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5828 = _T_337 ? _GEN_5813 : _GEN_5441; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5829 = _T_337 ? _GEN_5814 : _GEN_5442; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5830 = _T_337 ? _GEN_5815 : _GEN_5443; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5831 = _T_337 ? _GEN_5816 : _GEN_5446; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5832 = _T_337 ? _GEN_5817 : _GEN_5447; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5833 = _T_337 ? _GEN_5818 : _GEN_5448; // @[ISA.scala 390:85:@177411.8]
    assign _GEN_5834 = _T_85 ? _GEN_5819 : _GEN_5432; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5835 = _T_85 ? _GEN_5820 : _GEN_5433; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5836 = _T_85 ? _GEN_5821 : _GEN_5434; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5837 = _T_85 ? _GEN_5822 : _GEN_5435; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5838 = _T_85 ? _GEN_5823 : _GEN_5436; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5839 = _T_85 ? _GEN_5824 : _GEN_5437; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5840 = _T_85 ? _GEN_5825 : _GEN_5438; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5841 = _T_85 ? _GEN_5826 : _GEN_5439; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5842 = _T_85 ? _GEN_5827 : _GEN_5440; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5843 = _T_85 ? _GEN_5828 : _GEN_5441; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5844 = _T_85 ? _GEN_5829 : _GEN_5442; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5845 = _T_85 ? _GEN_5830 : _GEN_5443; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5846 = _T_85 ? _GEN_5831 : _GEN_5446; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5847 = _T_85 ? _GEN_5832 : _GEN_5447; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_5848 = _T_85 ? _GEN_5833 : _GEN_5448; // @[ISA.scala 389:44:@177239.6]
    assign _GEN_6038 = io_fromMemoryPort_sync ? 3'h4 : _GEN_5834; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6039 = io_fromMemoryPort_sync ? {{32'd0}, _T_223493} : _GEN_5835; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6040 = io_fromMemoryPort_sync ? 32'h0 : _GEN_5836; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6041 = io_fromMemoryPort_sync ? 32'h1 : _GEN_5837; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6042 = io_fromMemoryPort_sync ? 32'h1 : _GEN_5838; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6043 = io_fromMemoryPort_sync ? _T_223493 : _GEN_5839; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6044 = io_fromMemoryPort_sync ? _GEN_352 : _GEN_5840; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6045 = io_fromMemoryPort_sync ? {{32'd0}, _T_50} : _GEN_5841; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6046 = io_fromMemoryPort_sync ? {{32'd0}, _T_223493} : _GEN_5842; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6047 = io_fromMemoryPort_sync ? 32'h0 : _GEN_5843; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6048 = io_fromMemoryPort_sync ? 32'h1 : _GEN_5844; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6049 = io_fromMemoryPort_sync ? 32'h1 : _GEN_5845; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6050 = io_fromMemoryPort_sync ? _GEN_352 : _GEN_5444; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6051 = io_fromMemoryPort_sync ? {{32'd0}, _T_50} : _GEN_5445; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6052 = io_fromMemoryPort_sync ? 1'h0 : _GEN_5846; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6053 = io_fromMemoryPort_sync ? 1'h1 : _GEN_5847; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6054 = io_fromMemoryPort_sync ? 1'h1 : _GEN_5848; // @[ISA.scala 431:118:@187863.24]
    assign _GEN_6055 = _T_2036 ? _GEN_6038 : _GEN_5834; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6056 = _T_2036 ? _GEN_6039 : _GEN_5835; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6057 = _T_2036 ? _GEN_6040 : _GEN_5836; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6058 = _T_2036 ? _GEN_6041 : _GEN_5837; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6059 = _T_2036 ? _GEN_6042 : _GEN_5838; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6060 = _T_2036 ? _GEN_6043 : _GEN_5839; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6061 = _T_2036 ? _GEN_6044 : _GEN_5840; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6062 = _T_2036 ? _GEN_6045 : _GEN_5841; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6063 = _T_2036 ? _GEN_6046 : _GEN_5842; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6064 = _T_2036 ? _GEN_6047 : _GEN_5843; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6065 = _T_2036 ? _GEN_6048 : _GEN_5844; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6066 = _T_2036 ? _GEN_6049 : _GEN_5845; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6067 = _T_2036 ? _GEN_6050 : _GEN_5444; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6068 = _T_2036 ? _GEN_6051 : _GEN_5445; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6069 = _T_2036 ? _GEN_6052 : _GEN_5846; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6070 = _T_2036 ? _GEN_6053 : _GEN_5847; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6071 = _T_2036 ? _GEN_6054 : _GEN_5848; // @[ISA.scala 430:142:@187862.22]
    assign _GEN_6072 = _T_1795 ? _GEN_6055 : _GEN_5834; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6073 = _T_1795 ? _GEN_6056 : _GEN_5835; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6074 = _T_1795 ? _GEN_6057 : _GEN_5836; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6075 = _T_1795 ? _GEN_6058 : _GEN_5837; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6076 = _T_1795 ? _GEN_6059 : _GEN_5838; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6077 = _T_1795 ? _GEN_6060 : _GEN_5839; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6078 = _T_1795 ? _GEN_6061 : _GEN_5840; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6079 = _T_1795 ? _GEN_6062 : _GEN_5841; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6080 = _T_1795 ? _GEN_6063 : _GEN_5842; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6081 = _T_1795 ? _GEN_6064 : _GEN_5843; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6082 = _T_1795 ? _GEN_6065 : _GEN_5844; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6083 = _T_1795 ? _GEN_6066 : _GEN_5845; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6084 = _T_1795 ? _GEN_6067 : _GEN_5444; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6085 = _T_1795 ? _GEN_6068 : _GEN_5445; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6086 = _T_1795 ? _GEN_6069 : _GEN_5846; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6087 = _T_1795 ? _GEN_6070 : _GEN_5847; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6088 = _T_1795 ? _GEN_6071 : _GEN_5848; // @[ISA.scala 429:135:@187691.20]
    assign _GEN_6089 = _T_1552 ? _GEN_6072 : _GEN_5834; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6090 = _T_1552 ? _GEN_6073 : _GEN_5835; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6091 = _T_1552 ? _GEN_6074 : _GEN_5836; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6092 = _T_1552 ? _GEN_6075 : _GEN_5837; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6093 = _T_1552 ? _GEN_6076 : _GEN_5838; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6094 = _T_1552 ? _GEN_6077 : _GEN_5839; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6095 = _T_1552 ? _GEN_6078 : _GEN_5840; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6096 = _T_1552 ? _GEN_6079 : _GEN_5841; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6097 = _T_1552 ? _GEN_6080 : _GEN_5842; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6098 = _T_1552 ? _GEN_6081 : _GEN_5843; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6099 = _T_1552 ? _GEN_6082 : _GEN_5844; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6100 = _T_1552 ? _GEN_6083 : _GEN_5845; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6101 = _T_1552 ? _GEN_6084 : _GEN_5444; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6102 = _T_1552 ? _GEN_6085 : _GEN_5445; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6103 = _T_1552 ? _GEN_6086 : _GEN_5846; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6104 = _T_1552 ? _GEN_6087 : _GEN_5847; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6105 = _T_1552 ? _GEN_6088 : _GEN_5848; // @[ISA.scala 428:127:@187519.18]
    assign _GEN_6106 = _T_1309 ? _GEN_6089 : _GEN_5834; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6107 = _T_1309 ? _GEN_6090 : _GEN_5835; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6108 = _T_1309 ? _GEN_6091 : _GEN_5836; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6109 = _T_1309 ? _GEN_6092 : _GEN_5837; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6110 = _T_1309 ? _GEN_6093 : _GEN_5838; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6111 = _T_1309 ? _GEN_6094 : _GEN_5839; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6112 = _T_1309 ? _GEN_6095 : _GEN_5840; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6113 = _T_1309 ? _GEN_6096 : _GEN_5841; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6114 = _T_1309 ? _GEN_6097 : _GEN_5842; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6115 = _T_1309 ? _GEN_6098 : _GEN_5843; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6116 = _T_1309 ? _GEN_6099 : _GEN_5844; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6117 = _T_1309 ? _GEN_6100 : _GEN_5845; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6118 = _T_1309 ? _GEN_6101 : _GEN_5444; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6119 = _T_1309 ? _GEN_6102 : _GEN_5445; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6120 = _T_1309 ? _GEN_6103 : _GEN_5846; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6121 = _T_1309 ? _GEN_6104 : _GEN_5847; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6122 = _T_1309 ? _GEN_6105 : _GEN_5848; // @[ISA.scala 427:117:@187347.16]
    assign _GEN_6123 = _T_1066 ? _GEN_6106 : _GEN_5834; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6124 = _T_1066 ? _GEN_6107 : _GEN_5835; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6125 = _T_1066 ? _GEN_6108 : _GEN_5836; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6126 = _T_1066 ? _GEN_6109 : _GEN_5837; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6127 = _T_1066 ? _GEN_6110 : _GEN_5838; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6128 = _T_1066 ? _GEN_6111 : _GEN_5839; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6129 = _T_1066 ? _GEN_6112 : _GEN_5840; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6130 = _T_1066 ? _GEN_6113 : _GEN_5841; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6131 = _T_1066 ? _GEN_6114 : _GEN_5842; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6132 = _T_1066 ? _GEN_6115 : _GEN_5843; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6133 = _T_1066 ? _GEN_6116 : _GEN_5844; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6134 = _T_1066 ? _GEN_6117 : _GEN_5845; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6135 = _T_1066 ? _GEN_6118 : _GEN_5444; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6136 = _T_1066 ? _GEN_6119 : _GEN_5445; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6137 = _T_1066 ? _GEN_6120 : _GEN_5846; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6138 = _T_1066 ? _GEN_6121 : _GEN_5847; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6139 = _T_1066 ? _GEN_6122 : _GEN_5848; // @[ISA.scala 426:109:@187175.14]
    assign _GEN_6140 = _T_823 ? _GEN_6123 : _GEN_5834; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6141 = _T_823 ? _GEN_6124 : _GEN_5835; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6142 = _T_823 ? _GEN_6125 : _GEN_5836; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6143 = _T_823 ? _GEN_6126 : _GEN_5837; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6144 = _T_823 ? _GEN_6127 : _GEN_5838; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6145 = _T_823 ? _GEN_6128 : _GEN_5839; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6146 = _T_823 ? _GEN_6129 : _GEN_5840; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6147 = _T_823 ? _GEN_6130 : _GEN_5841; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6148 = _T_823 ? _GEN_6131 : _GEN_5842; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6149 = _T_823 ? _GEN_6132 : _GEN_5843; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6150 = _T_823 ? _GEN_6133 : _GEN_5844; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6151 = _T_823 ? _GEN_6134 : _GEN_5845; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6152 = _T_823 ? _GEN_6135 : _GEN_5444; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6153 = _T_823 ? _GEN_6136 : _GEN_5445; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6154 = _T_823 ? _GEN_6137 : _GEN_5846; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6155 = _T_823 ? _GEN_6138 : _GEN_5847; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6156 = _T_823 ? _GEN_6139 : _GEN_5848; // @[ISA.scala 425:101:@187003.12]
    assign _GEN_6157 = _T_580 ? _GEN_6140 : _GEN_5834; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6158 = _T_580 ? _GEN_6141 : _GEN_5835; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6159 = _T_580 ? _GEN_6142 : _GEN_5836; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6160 = _T_580 ? _GEN_6143 : _GEN_5837; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6161 = _T_580 ? _GEN_6144 : _GEN_5838; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6162 = _T_580 ? _GEN_6145 : _GEN_5839; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6163 = _T_580 ? _GEN_6146 : _GEN_5840; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6164 = _T_580 ? _GEN_6147 : _GEN_5841; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6165 = _T_580 ? _GEN_6148 : _GEN_5842; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6166 = _T_580 ? _GEN_6149 : _GEN_5843; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6167 = _T_580 ? _GEN_6150 : _GEN_5844; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6168 = _T_580 ? _GEN_6151 : _GEN_5845; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6169 = _T_580 ? _GEN_6152 : _GEN_5444; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6170 = _T_580 ? _GEN_6153 : _GEN_5445; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6171 = _T_580 ? _GEN_6154 : _GEN_5846; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6172 = _T_580 ? _GEN_6155 : _GEN_5847; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6173 = _T_580 ? _GEN_6156 : _GEN_5848; // @[ISA.scala 424:93:@186831.10]
    assign _GEN_6174 = _T_337 ? _GEN_6157 : _GEN_5834; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6175 = _T_337 ? _GEN_6158 : _GEN_5835; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6176 = _T_337 ? _GEN_6159 : _GEN_5836; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6177 = _T_337 ? _GEN_6160 : _GEN_5837; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6178 = _T_337 ? _GEN_6161 : _GEN_5838; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6179 = _T_337 ? _GEN_6162 : _GEN_5839; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6180 = _T_337 ? _GEN_6163 : _GEN_5840; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6181 = _T_337 ? _GEN_6164 : _GEN_5841; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6182 = _T_337 ? _GEN_6165 : _GEN_5842; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6183 = _T_337 ? _GEN_6166 : _GEN_5843; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6184 = _T_337 ? _GEN_6167 : _GEN_5844; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6185 = _T_337 ? _GEN_6168 : _GEN_5845; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6186 = _T_337 ? _GEN_6169 : _GEN_5444; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6187 = _T_337 ? _GEN_6170 : _GEN_5445; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6188 = _T_337 ? _GEN_6171 : _GEN_5846; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6189 = _T_337 ? _GEN_6172 : _GEN_5847; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6190 = _T_337 ? _GEN_6173 : _GEN_5848; // @[ISA.scala 423:85:@186659.8]
    assign _GEN_6191 = _T_85 ? _GEN_6174 : _GEN_5834; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6192 = _T_85 ? _GEN_6175 : _GEN_5835; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6193 = _T_85 ? _GEN_6176 : _GEN_5836; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6194 = _T_85 ? _GEN_6177 : _GEN_5837; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6195 = _T_85 ? _GEN_6178 : _GEN_5838; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6196 = _T_85 ? _GEN_6179 : _GEN_5839; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6197 = _T_85 ? _GEN_6180 : _GEN_5840; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6198 = _T_85 ? _GEN_6181 : _GEN_5841; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6199 = _T_85 ? _GEN_6182 : _GEN_5842; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6200 = _T_85 ? _GEN_6183 : _GEN_5843; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6201 = _T_85 ? _GEN_6184 : _GEN_5844; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6202 = _T_85 ? _GEN_6185 : _GEN_5845; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6203 = _T_85 ? _GEN_6186 : _GEN_5444; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6204 = _T_85 ? _GEN_6187 : _GEN_5445; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6205 = _T_85 ? _GEN_6188 : _GEN_5846; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6206 = _T_85 ? _GEN_6189 : _GEN_5847; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6207 = _T_85 ? _GEN_6190 : _GEN_5848; // @[ISA.scala 422:44:@186487.6]
    assign _GEN_6209 = reset ? 64'h0 : _GEN_6192; // @[ISA.scala 87:28:@18.4]
    assign _GEN_6215 = reset ? 64'h0 : _GEN_6198; // @[ISA.scala 87:28:@18.4]
    assign _GEN_6216 = reset ? 64'h0 : _GEN_6199; // @[ISA.scala 87:28:@18.4]
    assign _GEN_6224 = reset ? {{32'd0}, toRegsPort_r_dstData} : _GEN_6204; // @[ISA.scala 87:28:@18.4]
    assign io_fromMemoryPort_notify = fromMemoryPort_notify_r; // @[ISA.scala 465:34:@193602.4]
    assign io_toMemoryPort_notify = toMemoryPort_notify_r; // @[ISA.scala 466:32:@193603.4]
    assign io_toRegsPort_notify = toRegsPort_notify_r; // @[ISA.scala 467:30:@193604.4]
    assign io_toMemoryPort_addrIn = toMemoryPort_r_addrIn; // @[ISA.scala 468:25:@193608.4]
    assign io_toMemoryPort_dataIn = toMemoryPort_r_dataIn; // @[ISA.scala 468:25:@193607.4]
    assign io_toMemoryPort_mask = toMemoryPort_r_mask; // @[ISA.scala 468:25:@193606.4]
    assign io_toMemoryPort_req = toMemoryPort_r_req; // @[ISA.scala 468:25:@193605.4]
    assign io_toRegsPort_dst = toRegsPort_r_dst; // @[ISA.scala 469:23:@193610.4]
    assign io_toRegsPort_dstData = toRegsPort_r_dstData; // @[ISA.scala 469:23:@193609.4]
    `ifdef RANDOMIZE_GARBAGE_ASSIGN
    `define RANDOMIZE
    `endif
    `ifdef RANDOMIZE_INVALID_ASSIGN
    `define RANDOMIZE
    `endif
    `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
    `endif
    `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
    `endif
    `ifndef RANDOM
    `define RANDOM $random
    `endif
    `ifdef RANDOMIZE
    integer initvar;
    initial begin
    `ifdef INIT_RANDOM
    `INIT_RANDOM
    `endif
    `ifndef VERILATOR
    #0.002 begin end
    `endif
    `ifdef RANDOMIZE_REG_INIT
    _RAND_0 = {1{`RANDOM}};
    fromMemoryPort_notify_r = _RAND_0[0:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_1 = {1{`RANDOM}};
    toMemoryPort_notify_r = _RAND_1[0:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_2 = {1{`RANDOM}};
    toRegsPort_notify_r = _RAND_2[0:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_3 = {1{`RANDOM}};
    toMemoryPort_r_addrIn = _RAND_3[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_4 = {1{`RANDOM}};
    toMemoryPort_r_dataIn = _RAND_4[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_5 = {1{`RANDOM}};
    toMemoryPort_r_mask = _RAND_5[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_6 = {1{`RANDOM}};
    toMemoryPort_r_req = _RAND_6[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_7 = {1{`RANDOM}};
    toRegsPort_r_dst = _RAND_7[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_8 = {1{`RANDOM}};
    toRegsPort_r_dstData = _RAND_8[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_9 = {1{`RANDOM}};
    memoryAccess_signal_r_addrIn = _RAND_9[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_10 = {1{`RANDOM}};
    memoryAccess_signal_r_dataIn = _RAND_10[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_11 = {1{`RANDOM}};
    memoryAccess_signal_r_mask = _RAND_11[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_12 = {1{`RANDOM}};
    memoryAccess_signal_r_req = _RAND_12[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_13 = {1{`RANDOM}};
    pcReg_signal_r = _RAND_13[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_14 = {1{`RANDOM}};
    regfileWrite_signal_r_dst = _RAND_14[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_15 = {1{`RANDOM}};
    regfileWrite_signal_r_dstData = _RAND_15[31:0];
    `endif // RANDOMIZE_REG_INIT
    `ifdef RANDOMIZE_REG_INIT
    _RAND_16 = {1{`RANDOM}};
    state_r = _RAND_16[2:0];
    `endif // RANDOMIZE_REG_INIT
    end
    `endif
    // RANDOMIZE
    always @(posedge clock) begin
        if (reset) begin
            fromMemoryPort_notify_r <= 1'h0;
        end else begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    fromMemoryPort_notify_r <= 1'h0;
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1552) begin
                                                                                if (_T_1793) begin
                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                        fromMemoryPort_notify_r <= 1'h0;
                                                                                    end else begin
                                                                                        if (_T_85) begin
                                                                                            if (_T_337) begin
                                                                                                if (_T_580) begin
                                                                                                    if (_T_823) begin
                                                                                                        if (_T_1066) begin
                                                                                                            if (_T_1309) begin
                                                                                                                if (_T_1550) begin
                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                        fromMemoryPort_notify_r <= 1'h0;
                                                                                                                    end else begin
                                                                                                                        if (_T_85) begin
                                                                                                                            if (_T_337) begin
                                                                                                                                if (_T_580) begin
                                                                                                                                    if (_T_823) begin
                                                                                                                                        if (_T_1066) begin
                                                                                                                                            if (_T_1307) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_85) begin
                                                                                                                                                        if (_T_337) begin
                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                    if (_T_1064) begin
                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                            fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                        if (_T_821) begin
                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                                                        if (_T_578) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                                    if (_T_335) begin
                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                            fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                                                                        if (_T_823) begin
                                                                                                                                                                                                                                            if (_T_1066) begin
                                                                                                                                                                                                                                                if (_T_1309) begin
                                                                                                                                                                                                                                                    if (_T_1552) begin
                                                                                                                                                                                                                                                        if (_T_1795) begin
                                                                                                                                                                                                                                                            if (_T_2038) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_81) begin
                                                                                                                                                                                                                                                                        if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_66) begin
                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_62) begin
                                                                                                                                                                                                                                                                                        if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_47) begin
                                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                    if (_T_43) begin
                                                                                                                                                                                                                                                                                                        if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_43) begin
                                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_43) begin
                                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_43) begin
                                                                                                                                                                                                                                                                                                if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_19;
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_19;
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_47) begin
                                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_19;
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_19;
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_49;
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_49;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_62) begin
                                                                                                                                                                                                                                                                                if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_49;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_49;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_81) begin
                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_71;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_71;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_66) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_71;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_71;
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_81) begin
                                                                                                                                                                                                                                                                if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_105;
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_105;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_81) begin
                                                                                                                                                                                                                                                            if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_105;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_105;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                                                                                    if (_T_1066) begin
                                                                                                                                                                                                                                        if (_T_1309) begin
                                                                                                                                                                                                                                            if (_T_1552) begin
                                                                                                                                                                                                                                                if (_T_1795) begin
                                                                                                                                                                                                                                                    if (_T_2038) begin
                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                if (_T_335) begin
                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                        fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_127;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_341;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_341;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                    fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_341;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_341;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_341;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                        if (_T_335) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_341;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_341;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_341;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                    if (_T_578) begin
                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                            fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_670;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_670;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_670;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_670;
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                if (_T_578) begin
                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                        fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_670;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_670;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_670;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_670;
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                            if (_T_578) begin
                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                    fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_670;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_670;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_670;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_670;
                                                                                                                                                                                    end
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                            end
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                    if (_T_821) begin
                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                            fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                        end
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                if (_T_821) begin
                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                        fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                    end
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                        if (_T_580) begin
                                                                                                                                                                            if (_T_821) begin
                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                    fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                end else begin
                                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4163;
                                                                                                                                                                end
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_85) begin
                                                                                                                                                    if (_T_337) begin
                                                                                                                                                        if (_T_580) begin
                                                                                                                                                            if (_T_823) begin
                                                                                                                                                                if (_T_1064) begin
                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                        fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_85) begin
                                                                                                                                                if (_T_337) begin
                                                                                                                                                    if (_T_580) begin
                                                                                                                                                        if (_T_823) begin
                                                                                                                                                            if (_T_1064) begin
                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                    fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_337) begin
                                                                                                                                                if (_T_580) begin
                                                                                                                                                    if (_T_823) begin
                                                                                                                                                        if (_T_1064) begin
                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                                            end else begin
                                                                                                                                                                fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            fromMemoryPort_notify_r <= _GEN_4534;
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                        end
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    if (_T_85) begin
                                                                                                                        if (_T_337) begin
                                                                                                                            if (_T_580) begin
                                                                                                                                if (_T_823) begin
                                                                                                                                    if (_T_1066) begin
                                                                                                                                        if (_T_1307) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                            end else begin
                                                                                                                                                fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                    end
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1066) begin
                                                                                                                                    if (_T_1307) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                        end else begin
                                                                                                                                            fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1066) begin
                                                                                                                                if (_T_1307) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        fromMemoryPort_notify_r <= 1'h0;
                                                                                                                                    end else begin
                                                                                                                                        fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                fromMemoryPort_notify_r <= _GEN_4850;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                    end
                                                                                                end else begin
                                                                                                    fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                end
                                                                                            end else begin
                                                                                                fromMemoryPort_notify_r <= _GEN_5038;
                                                                                            end
                                                                                        end else begin
                                                                                            fromMemoryPort_notify_r <= _GEN_5038;
                                                                                        end
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1309) begin
                                                                                                            if (_T_1550) begin
                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                    fromMemoryPort_notify_r <= 1'h0;
                                                                                                                end else begin
                                                                                                                    fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                    end
                                                                                                end else begin
                                                                                                    fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                end
                                                                                            end else begin
                                                                                                fromMemoryPort_notify_r <= _GEN_5038;
                                                                                            end
                                                                                        end else begin
                                                                                            fromMemoryPort_notify_r <= _GEN_5038;
                                                                                        end
                                                                                    end else begin
                                                                                        fromMemoryPort_notify_r <= _GEN_5038;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1309) begin
                                                                                                        if (_T_1550) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                                                            end else begin
                                                                                                                fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                    end
                                                                                                end else begin
                                                                                                    fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                end
                                                                                            end else begin
                                                                                                fromMemoryPort_notify_r <= _GEN_5038;
                                                                                            end
                                                                                        end else begin
                                                                                            fromMemoryPort_notify_r <= _GEN_5038;
                                                                                        end
                                                                                    end else begin
                                                                                        fromMemoryPort_notify_r <= _GEN_5038;
                                                                                    end
                                                                                end else begin
                                                                                    fromMemoryPort_notify_r <= _GEN_5038;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1309) begin
                                                                                                    if (_T_1550) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            fromMemoryPort_notify_r <= 1'h0;
                                                                                                        end else begin
                                                                                                            fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                    end
                                                                                                end else begin
                                                                                                    fromMemoryPort_notify_r <= _GEN_5038;
                                                                                                end
                                                                                            end else begin
                                                                                                fromMemoryPort_notify_r <= _GEN_5038;
                                                                                            end
                                                                                        end else begin
                                                                                            fromMemoryPort_notify_r <= _GEN_5038;
                                                                                        end
                                                                                    end else begin
                                                                                        fromMemoryPort_notify_r <= _GEN_5038;
                                                                                    end
                                                                                end else begin
                                                                                    fromMemoryPort_notify_r <= _GEN_5038;
                                                                                end
                                                                            end else begin
                                                                                fromMemoryPort_notify_r <= _GEN_5038;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        fromMemoryPort_notify_r <= _GEN_5446;
                                                                    end
                                                                end else begin
                                                                    fromMemoryPort_notify_r <= _GEN_5446;
                                                                end
                                                            end else begin
                                                                fromMemoryPort_notify_r <= _GEN_5446;
                                                            end
                                                        end else begin
                                                            fromMemoryPort_notify_r <= _GEN_5446;
                                                        end
                                                    end else begin
                                                        fromMemoryPort_notify_r <= _GEN_5446;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1552) begin
                                                                            if (_T_1793) begin
                                                                                if (io_fromMemoryPort_sync) begin
                                                                                    fromMemoryPort_notify_r <= 1'h0;
                                                                                end else begin
                                                                                    fromMemoryPort_notify_r <= _GEN_5446;
                                                                                end
                                                                            end else begin
                                                                                fromMemoryPort_notify_r <= _GEN_5446;
                                                                            end
                                                                        end else begin
                                                                            fromMemoryPort_notify_r <= _GEN_5446;
                                                                        end
                                                                    end else begin
                                                                        fromMemoryPort_notify_r <= _GEN_5446;
                                                                    end
                                                                end else begin
                                                                    fromMemoryPort_notify_r <= _GEN_5446;
                                                                end
                                                            end else begin
                                                                fromMemoryPort_notify_r <= _GEN_5446;
                                                            end
                                                        end else begin
                                                            fromMemoryPort_notify_r <= _GEN_5446;
                                                        end
                                                    end else begin
                                                        fromMemoryPort_notify_r <= _GEN_5446;
                                                    end
                                                end else begin
                                                    fromMemoryPort_notify_r <= _GEN_5446;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1552) begin
                                                                        if (_T_1793) begin
                                                                            if (io_fromMemoryPort_sync) begin
                                                                                fromMemoryPort_notify_r <= 1'h0;
                                                                            end else begin
                                                                                fromMemoryPort_notify_r <= _GEN_5446;
                                                                            end
                                                                        end else begin
                                                                            fromMemoryPort_notify_r <= _GEN_5446;
                                                                        end
                                                                    end else begin
                                                                        fromMemoryPort_notify_r <= _GEN_5446;
                                                                    end
                                                                end else begin
                                                                    fromMemoryPort_notify_r <= _GEN_5446;
                                                                end
                                                            end else begin
                                                                fromMemoryPort_notify_r <= _GEN_5446;
                                                            end
                                                        end else begin
                                                            fromMemoryPort_notify_r <= _GEN_5446;
                                                        end
                                                    end else begin
                                                        fromMemoryPort_notify_r <= _GEN_5446;
                                                    end
                                                end else begin
                                                    fromMemoryPort_notify_r <= _GEN_5446;
                                                end
                                            end else begin
                                                fromMemoryPort_notify_r <= _GEN_5446;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1552) begin
                                                                    if (_T_1793) begin
                                                                        if (io_fromMemoryPort_sync) begin
                                                                            fromMemoryPort_notify_r <= 1'h0;
                                                                        end else begin
                                                                            fromMemoryPort_notify_r <= _GEN_5446;
                                                                        end
                                                                    end else begin
                                                                        fromMemoryPort_notify_r <= _GEN_5446;
                                                                    end
                                                                end else begin
                                                                    fromMemoryPort_notify_r <= _GEN_5446;
                                                                end
                                                            end else begin
                                                                fromMemoryPort_notify_r <= _GEN_5446;
                                                            end
                                                        end else begin
                                                            fromMemoryPort_notify_r <= _GEN_5446;
                                                        end
                                                    end else begin
                                                        fromMemoryPort_notify_r <= _GEN_5446;
                                                    end
                                                end else begin
                                                    fromMemoryPort_notify_r <= _GEN_5446;
                                                end
                                            end else begin
                                                fromMemoryPort_notify_r <= _GEN_5446;
                                            end
                                        end else begin
                                            fromMemoryPort_notify_r <= _GEN_5446;
                                        end
                                    end
                                end else begin
                                    fromMemoryPort_notify_r <= _GEN_5846;
                                end
                            end else begin
                                fromMemoryPort_notify_r <= _GEN_5846;
                            end
                        end else begin
                            fromMemoryPort_notify_r <= _GEN_5846;
                        end
                    end else begin
                        fromMemoryPort_notify_r <= _GEN_5846;
                    end
                end else begin
                    fromMemoryPort_notify_r <= _GEN_5846;
                end
            end else begin
                fromMemoryPort_notify_r <= _GEN_5846;
            end
        end
        if (reset) begin
            toMemoryPort_notify_r <= 1'h1;
        end else begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    toMemoryPort_notify_r <= 1'h1;
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1552) begin
                                                                                if (_T_1793) begin
                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                        toMemoryPort_notify_r <= 1'h1;
                                                                                    end else begin
                                                                                        if (_T_85) begin
                                                                                            if (_T_337) begin
                                                                                                if (_T_580) begin
                                                                                                    if (_T_823) begin
                                                                                                        if (_T_1066) begin
                                                                                                            if (_T_1309) begin
                                                                                                                if (_T_1550) begin
                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                        toMemoryPort_notify_r <= 1'h1;
                                                                                                                    end else begin
                                                                                                                        if (_T_85) begin
                                                                                                                            if (_T_337) begin
                                                                                                                                if (_T_580) begin
                                                                                                                                    if (_T_823) begin
                                                                                                                                        if (_T_1066) begin
                                                                                                                                            if (_T_1307) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_85) begin
                                                                                                                                                        if (_T_337) begin
                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                    if (_T_1064) begin
                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                            toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                        end else begin
                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                        if (_T_821) begin
                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                                                        if (_T_578) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                                    if (_T_335) begin
                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                            toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                                                                        if (_T_823) begin
                                                                                                                                                                                                                                            if (_T_1066) begin
                                                                                                                                                                                                                                                if (_T_1309) begin
                                                                                                                                                                                                                                                    if (_T_1552) begin
                                                                                                                                                                                                                                                        if (_T_1795) begin
                                                                                                                                                                                                                                                            if (_T_2038) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_81) begin
                                                                                                                                                                                                                                                                        if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_66) begin
                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_62) begin
                                                                                                                                                                                                                                                                                        if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_47) begin
                                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                    if (_T_43) begin
                                                                                                                                                                                                                                                                                                        if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_43) begin
                                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                        toMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_43) begin
                                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                        toMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_43) begin
                                                                                                                                                                                                                                                                                                if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                        toMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_20;
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_20;
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_47) begin
                                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_20;
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_20;
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                        toMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_50;
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_50;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_62) begin
                                                                                                                                                                                                                                                                                if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_50;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_50;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_81) begin
                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                        toMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_72;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_72;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_66) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_72;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_72;
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_81) begin
                                                                                                                                                                                                                                                                if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_106;
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_106;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_81) begin
                                                                                                                                                                                                                                                            if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_106;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_106;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                                                                                    if (_T_1066) begin
                                                                                                                                                                                                                                        if (_T_1309) begin
                                                                                                                                                                                                                                            if (_T_1552) begin
                                                                                                                                                                                                                                                if (_T_1795) begin
                                                                                                                                                                                                                                                    if (_T_2038) begin
                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                if (_T_335) begin
                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                        toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_128;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_342;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_342;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                    toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_342;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_342;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_342;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                        if (_T_335) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_342;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_342;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_342;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                    if (_T_578) begin
                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                            toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_671;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_671;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_671;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_671;
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                if (_T_578) begin
                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                        toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_671;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_671;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_671;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_671;
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                            if (_T_578) begin
                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                    toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_671;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_671;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_671;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_671;
                                                                                                                                                                                    end
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                            end
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                    if (_T_821) begin
                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                            toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                        end
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                if (_T_821) begin
                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                        toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                    end
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                        if (_T_580) begin
                                                                                                                                                                            if (_T_821) begin
                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                    toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_4164;
                                                                                                                                                                end
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_85) begin
                                                                                                                                                    if (_T_337) begin
                                                                                                                                                        if (_T_580) begin
                                                                                                                                                            if (_T_823) begin
                                                                                                                                                                if (_T_1064) begin
                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                        toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                    end else begin
                                                                                                                                                                        toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_85) begin
                                                                                                                                                if (_T_337) begin
                                                                                                                                                    if (_T_580) begin
                                                                                                                                                        if (_T_823) begin
                                                                                                                                                            if (_T_1064) begin
                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                    toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                                end else begin
                                                                                                                                                                    toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_337) begin
                                                                                                                                                if (_T_580) begin
                                                                                                                                                    if (_T_823) begin
                                                                                                                                                        if (_T_1064) begin
                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                                                                                                            end else begin
                                                                                                                                                                toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            toMemoryPort_notify_r <= _GEN_4535;
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                        end
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    if (_T_85) begin
                                                                                                                        if (_T_337) begin
                                                                                                                            if (_T_580) begin
                                                                                                                                if (_T_823) begin
                                                                                                                                    if (_T_1066) begin
                                                                                                                                        if (_T_1307) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                                                                                            end else begin
                                                                                                                                                toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                    end
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1066) begin
                                                                                                                                    if (_T_1307) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            toMemoryPort_notify_r <= 1'h1;
                                                                                                                                        end else begin
                                                                                                                                            toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1066) begin
                                                                                                                                if (_T_1307) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        toMemoryPort_notify_r <= 1'h1;
                                                                                                                                    end else begin
                                                                                                                                        toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toMemoryPort_notify_r <= _GEN_4851;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toMemoryPort_notify_r <= _GEN_4851;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_notify_r <= _GEN_5039;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_notify_r <= _GEN_5039;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_notify_r <= _GEN_5039;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_notify_r <= _GEN_5039;
                                                                                        end
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1309) begin
                                                                                                            if (_T_1550) begin
                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                    toMemoryPort_notify_r <= 1'h1;
                                                                                                                end else begin
                                                                                                                    toMemoryPort_notify_r <= _GEN_5039;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toMemoryPort_notify_r <= _GEN_5039;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            toMemoryPort_notify_r <= _GEN_5039;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_notify_r <= _GEN_5039;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_notify_r <= _GEN_5039;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_notify_r <= _GEN_5039;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_notify_r <= _GEN_5039;
                                                                                        end
                                                                                    end else begin
                                                                                        toMemoryPort_notify_r <= _GEN_5039;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1309) begin
                                                                                                        if (_T_1550) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                                                            end else begin
                                                                                                                toMemoryPort_notify_r <= _GEN_5039;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            toMemoryPort_notify_r <= _GEN_5039;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_notify_r <= _GEN_5039;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_notify_r <= _GEN_5039;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_notify_r <= _GEN_5039;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_notify_r <= _GEN_5039;
                                                                                        end
                                                                                    end else begin
                                                                                        toMemoryPort_notify_r <= _GEN_5039;
                                                                                    end
                                                                                end else begin
                                                                                    toMemoryPort_notify_r <= _GEN_5039;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1309) begin
                                                                                                    if (_T_1550) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            toMemoryPort_notify_r <= 1'h1;
                                                                                                        end else begin
                                                                                                            toMemoryPort_notify_r <= _GEN_5039;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_notify_r <= _GEN_5039;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_notify_r <= _GEN_5039;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_notify_r <= _GEN_5039;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_notify_r <= _GEN_5039;
                                                                                        end
                                                                                    end else begin
                                                                                        toMemoryPort_notify_r <= _GEN_5039;
                                                                                    end
                                                                                end else begin
                                                                                    toMemoryPort_notify_r <= _GEN_5039;
                                                                                end
                                                                            end else begin
                                                                                toMemoryPort_notify_r <= _GEN_5039;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_notify_r <= _GEN_5447;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_notify_r <= _GEN_5447;
                                                                end
                                                            end else begin
                                                                toMemoryPort_notify_r <= _GEN_5447;
                                                            end
                                                        end else begin
                                                            toMemoryPort_notify_r <= _GEN_5447;
                                                        end
                                                    end else begin
                                                        toMemoryPort_notify_r <= _GEN_5447;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1552) begin
                                                                            if (_T_1793) begin
                                                                                if (io_fromMemoryPort_sync) begin
                                                                                    toMemoryPort_notify_r <= 1'h1;
                                                                                end else begin
                                                                                    toMemoryPort_notify_r <= _GEN_5447;
                                                                                end
                                                                            end else begin
                                                                                toMemoryPort_notify_r <= _GEN_5447;
                                                                            end
                                                                        end else begin
                                                                            toMemoryPort_notify_r <= _GEN_5447;
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_notify_r <= _GEN_5447;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_notify_r <= _GEN_5447;
                                                                end
                                                            end else begin
                                                                toMemoryPort_notify_r <= _GEN_5447;
                                                            end
                                                        end else begin
                                                            toMemoryPort_notify_r <= _GEN_5447;
                                                        end
                                                    end else begin
                                                        toMemoryPort_notify_r <= _GEN_5447;
                                                    end
                                                end else begin
                                                    toMemoryPort_notify_r <= _GEN_5447;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1552) begin
                                                                        if (_T_1793) begin
                                                                            if (io_fromMemoryPort_sync) begin
                                                                                toMemoryPort_notify_r <= 1'h1;
                                                                            end else begin
                                                                                toMemoryPort_notify_r <= _GEN_5447;
                                                                            end
                                                                        end else begin
                                                                            toMemoryPort_notify_r <= _GEN_5447;
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_notify_r <= _GEN_5447;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_notify_r <= _GEN_5447;
                                                                end
                                                            end else begin
                                                                toMemoryPort_notify_r <= _GEN_5447;
                                                            end
                                                        end else begin
                                                            toMemoryPort_notify_r <= _GEN_5447;
                                                        end
                                                    end else begin
                                                        toMemoryPort_notify_r <= _GEN_5447;
                                                    end
                                                end else begin
                                                    toMemoryPort_notify_r <= _GEN_5447;
                                                end
                                            end else begin
                                                toMemoryPort_notify_r <= _GEN_5447;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1552) begin
                                                                    if (_T_1793) begin
                                                                        if (io_fromMemoryPort_sync) begin
                                                                            toMemoryPort_notify_r <= 1'h1;
                                                                        end else begin
                                                                            toMemoryPort_notify_r <= _GEN_5447;
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_notify_r <= _GEN_5447;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_notify_r <= _GEN_5447;
                                                                end
                                                            end else begin
                                                                toMemoryPort_notify_r <= _GEN_5447;
                                                            end
                                                        end else begin
                                                            toMemoryPort_notify_r <= _GEN_5447;
                                                        end
                                                    end else begin
                                                        toMemoryPort_notify_r <= _GEN_5447;
                                                    end
                                                end else begin
                                                    toMemoryPort_notify_r <= _GEN_5447;
                                                end
                                            end else begin
                                                toMemoryPort_notify_r <= _GEN_5447;
                                            end
                                        end else begin
                                            toMemoryPort_notify_r <= _GEN_5447;
                                        end
                                    end
                                end else begin
                                    toMemoryPort_notify_r <= _GEN_5847;
                                end
                            end else begin
                                toMemoryPort_notify_r <= _GEN_5847;
                            end
                        end else begin
                            toMemoryPort_notify_r <= _GEN_5847;
                        end
                    end else begin
                        toMemoryPort_notify_r <= _GEN_5847;
                    end
                end else begin
                    toMemoryPort_notify_r <= _GEN_5847;
                end
            end else begin
                toMemoryPort_notify_r <= _GEN_5847;
            end
        end
        if (reset) begin
            toRegsPort_notify_r <= 1'h0;
        end else begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    toRegsPort_notify_r <= 1'h1;
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1552) begin
                                                                                if (_T_1793) begin
                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                        toRegsPort_notify_r <= 1'h0;
                                                                                    end else begin
                                                                                        if (_T_85) begin
                                                                                            if (_T_337) begin
                                                                                                if (_T_580) begin
                                                                                                    if (_T_823) begin
                                                                                                        if (_T_1066) begin
                                                                                                            if (_T_1309) begin
                                                                                                                if (_T_1550) begin
                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                        toRegsPort_notify_r <= 1'h1;
                                                                                                                    end else begin
                                                                                                                        if (_T_85) begin
                                                                                                                            if (_T_337) begin
                                                                                                                                if (_T_580) begin
                                                                                                                                    if (_T_823) begin
                                                                                                                                        if (_T_1066) begin
                                                                                                                                            if (_T_1307) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    toRegsPort_notify_r <= 1'h1;
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_85) begin
                                                                                                                                                        if (_T_337) begin
                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                    if (_T_1064) begin
                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                            toRegsPort_notify_r <= 1'h1;
                                                                                                                                                                        end else begin
                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                        if (_T_821) begin
                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                                                        if (_T_578) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                                    if (_T_335) begin
                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                            toRegsPort_notify_r <= 1'h1;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                                                                        if (_T_823) begin
                                                                                                                                                                                                                                            if (_T_1066) begin
                                                                                                                                                                                                                                                if (_T_1309) begin
                                                                                                                                                                                                                                                    if (_T_1552) begin
                                                                                                                                                                                                                                                        if (_T_1795) begin
                                                                                                                                                                                                                                                            if (_T_2038) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_81) begin
                                                                                                                                                                                                                                                                        if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_66) begin
                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    toRegsPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_62) begin
                                                                                                                                                                                                                                                                                        if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                            toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_47) begin
                                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                    toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                    if (_T_43) begin
                                                                                                                                                                                                                                                                                                        if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                            toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_43) begin
                                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                        toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_43) begin
                                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                        toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_43) begin
                                                                                                                                                                                                                                                                                                if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                    toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                        toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_21;
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_21;
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_47) begin
                                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                            toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_21;
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_21;
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                toRegsPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                        toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_51;
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_51;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_62) begin
                                                                                                                                                                                                                                                                                if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_51;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_51;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_81) begin
                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                        toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                toRegsPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_73;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_73;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_66) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            toRegsPort_notify_r <= 1'h1;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_73;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_73;
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_81) begin
                                                                                                                                                                                                                                                                if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_107;
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_107;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_81) begin
                                                                                                                                                                                                                                                            if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_107;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_107;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                                                                                    if (_T_1066) begin
                                                                                                                                                                                                                                        if (_T_1309) begin
                                                                                                                                                                                                                                            if (_T_1552) begin
                                                                                                                                                                                                                                                if (_T_1795) begin
                                                                                                                                                                                                                                                    if (_T_2038) begin
                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                            toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                if (_T_335) begin
                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                        toRegsPort_notify_r <= 1'h1;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_129;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_343;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_343;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                    toRegsPort_notify_r <= 1'h1;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_343;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_343;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_343;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                        if (_T_335) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                toRegsPort_notify_r <= 1'h1;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_343;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_343;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_343;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                    if (_T_578) begin
                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                            toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_672;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_672;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_672;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_672;
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                if (_T_578) begin
                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                        toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_672;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_672;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_672;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_672;
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                            if (_T_578) begin
                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                    toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_672;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toRegsPort_notify_r <= _GEN_672;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_672;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_672;
                                                                                                                                                                                    end
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                            end
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                    if (_T_821) begin
                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                            toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                        end
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                if (_T_821) begin
                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                        toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                    end
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                        if (_T_580) begin
                                                                                                                                                                            if (_T_821) begin
                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                    toRegsPort_notify_r <= 1'h0;
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    toRegsPort_notify_r <= _GEN_4165;
                                                                                                                                                                end
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_85) begin
                                                                                                                                                    if (_T_337) begin
                                                                                                                                                        if (_T_580) begin
                                                                                                                                                            if (_T_823) begin
                                                                                                                                                                if (_T_1064) begin
                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                        toRegsPort_notify_r <= 1'h1;
                                                                                                                                                                    end else begin
                                                                                                                                                                        toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_85) begin
                                                                                                                                                if (_T_337) begin
                                                                                                                                                    if (_T_580) begin
                                                                                                                                                        if (_T_823) begin
                                                                                                                                                            if (_T_1064) begin
                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                    toRegsPort_notify_r <= 1'h1;
                                                                                                                                                                end else begin
                                                                                                                                                                    toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_337) begin
                                                                                                                                                if (_T_580) begin
                                                                                                                                                    if (_T_823) begin
                                                                                                                                                        if (_T_1064) begin
                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                toRegsPort_notify_r <= 1'h1;
                                                                                                                                                            end else begin
                                                                                                                                                                toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            toRegsPort_notify_r <= _GEN_4536;
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toRegsPort_notify_r <= _GEN_4852;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toRegsPort_notify_r <= _GEN_4852;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toRegsPort_notify_r <= _GEN_4852;
                                                                                                                        end
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    if (_T_85) begin
                                                                                                                        if (_T_337) begin
                                                                                                                            if (_T_580) begin
                                                                                                                                if (_T_823) begin
                                                                                                                                    if (_T_1066) begin
                                                                                                                                        if (_T_1307) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                toRegsPort_notify_r <= 1'h1;
                                                                                                                                            end else begin
                                                                                                                                                toRegsPort_notify_r <= _GEN_4852;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            toRegsPort_notify_r <= _GEN_4852;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        toRegsPort_notify_r <= _GEN_4852;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toRegsPort_notify_r <= _GEN_4852;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toRegsPort_notify_r <= _GEN_4852;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toRegsPort_notify_r <= _GEN_4852;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toRegsPort_notify_r <= _GEN_4852;
                                                                                                                    end
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1066) begin
                                                                                                                                    if (_T_1307) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            toRegsPort_notify_r <= 1'h1;
                                                                                                                                        end else begin
                                                                                                                                            toRegsPort_notify_r <= _GEN_4852;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        toRegsPort_notify_r <= _GEN_4852;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toRegsPort_notify_r <= _GEN_4852;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toRegsPort_notify_r <= _GEN_4852;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toRegsPort_notify_r <= _GEN_4852;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toRegsPort_notify_r <= _GEN_4852;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toRegsPort_notify_r <= _GEN_4852;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1066) begin
                                                                                                                                if (_T_1307) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        toRegsPort_notify_r <= 1'h1;
                                                                                                                                    end else begin
                                                                                                                                        toRegsPort_notify_r <= _GEN_4852;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toRegsPort_notify_r <= _GEN_4852;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toRegsPort_notify_r <= _GEN_4852;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toRegsPort_notify_r <= _GEN_4852;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toRegsPort_notify_r <= _GEN_4852;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toRegsPort_notify_r <= _GEN_4852;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toRegsPort_notify_r <= _GEN_4852;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toRegsPort_notify_r <= _GEN_5040;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toRegsPort_notify_r <= _GEN_5040;
                                                                                                end
                                                                                            end else begin
                                                                                                toRegsPort_notify_r <= _GEN_5040;
                                                                                            end
                                                                                        end else begin
                                                                                            toRegsPort_notify_r <= _GEN_5040;
                                                                                        end
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1309) begin
                                                                                                            if (_T_1550) begin
                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                    toRegsPort_notify_r <= 1'h1;
                                                                                                                end else begin
                                                                                                                    toRegsPort_notify_r <= _GEN_5040;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toRegsPort_notify_r <= _GEN_5040;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            toRegsPort_notify_r <= _GEN_5040;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toRegsPort_notify_r <= _GEN_5040;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toRegsPort_notify_r <= _GEN_5040;
                                                                                                end
                                                                                            end else begin
                                                                                                toRegsPort_notify_r <= _GEN_5040;
                                                                                            end
                                                                                        end else begin
                                                                                            toRegsPort_notify_r <= _GEN_5040;
                                                                                        end
                                                                                    end else begin
                                                                                        toRegsPort_notify_r <= _GEN_5040;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1309) begin
                                                                                                        if (_T_1550) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                toRegsPort_notify_r <= 1'h1;
                                                                                                            end else begin
                                                                                                                toRegsPort_notify_r <= _GEN_5040;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            toRegsPort_notify_r <= _GEN_5040;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toRegsPort_notify_r <= _GEN_5040;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toRegsPort_notify_r <= _GEN_5040;
                                                                                                end
                                                                                            end else begin
                                                                                                toRegsPort_notify_r <= _GEN_5040;
                                                                                            end
                                                                                        end else begin
                                                                                            toRegsPort_notify_r <= _GEN_5040;
                                                                                        end
                                                                                    end else begin
                                                                                        toRegsPort_notify_r <= _GEN_5040;
                                                                                    end
                                                                                end else begin
                                                                                    toRegsPort_notify_r <= _GEN_5040;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1309) begin
                                                                                                    if (_T_1550) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            toRegsPort_notify_r <= 1'h1;
                                                                                                        end else begin
                                                                                                            toRegsPort_notify_r <= _GEN_5040;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toRegsPort_notify_r <= _GEN_5040;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toRegsPort_notify_r <= _GEN_5040;
                                                                                                end
                                                                                            end else begin
                                                                                                toRegsPort_notify_r <= _GEN_5040;
                                                                                            end
                                                                                        end else begin
                                                                                            toRegsPort_notify_r <= _GEN_5040;
                                                                                        end
                                                                                    end else begin
                                                                                        toRegsPort_notify_r <= _GEN_5040;
                                                                                    end
                                                                                end else begin
                                                                                    toRegsPort_notify_r <= _GEN_5040;
                                                                                end
                                                                            end else begin
                                                                                toRegsPort_notify_r <= _GEN_5040;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        toRegsPort_notify_r <= _GEN_5448;
                                                                    end
                                                                end else begin
                                                                    toRegsPort_notify_r <= _GEN_5448;
                                                                end
                                                            end else begin
                                                                toRegsPort_notify_r <= _GEN_5448;
                                                            end
                                                        end else begin
                                                            toRegsPort_notify_r <= _GEN_5448;
                                                        end
                                                    end else begin
                                                        toRegsPort_notify_r <= _GEN_5448;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1552) begin
                                                                            if (_T_1793) begin
                                                                                if (io_fromMemoryPort_sync) begin
                                                                                    toRegsPort_notify_r <= 1'h0;
                                                                                end else begin
                                                                                    toRegsPort_notify_r <= _GEN_5448;
                                                                                end
                                                                            end else begin
                                                                                toRegsPort_notify_r <= _GEN_5448;
                                                                            end
                                                                        end else begin
                                                                            toRegsPort_notify_r <= _GEN_5448;
                                                                        end
                                                                    end else begin
                                                                        toRegsPort_notify_r <= _GEN_5448;
                                                                    end
                                                                end else begin
                                                                    toRegsPort_notify_r <= _GEN_5448;
                                                                end
                                                            end else begin
                                                                toRegsPort_notify_r <= _GEN_5448;
                                                            end
                                                        end else begin
                                                            toRegsPort_notify_r <= _GEN_5448;
                                                        end
                                                    end else begin
                                                        toRegsPort_notify_r <= _GEN_5448;
                                                    end
                                                end else begin
                                                    toRegsPort_notify_r <= _GEN_5448;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1552) begin
                                                                        if (_T_1793) begin
                                                                            if (io_fromMemoryPort_sync) begin
                                                                                toRegsPort_notify_r <= 1'h0;
                                                                            end else begin
                                                                                toRegsPort_notify_r <= _GEN_5448;
                                                                            end
                                                                        end else begin
                                                                            toRegsPort_notify_r <= _GEN_5448;
                                                                        end
                                                                    end else begin
                                                                        toRegsPort_notify_r <= _GEN_5448;
                                                                    end
                                                                end else begin
                                                                    toRegsPort_notify_r <= _GEN_5448;
                                                                end
                                                            end else begin
                                                                toRegsPort_notify_r <= _GEN_5448;
                                                            end
                                                        end else begin
                                                            toRegsPort_notify_r <= _GEN_5448;
                                                        end
                                                    end else begin
                                                        toRegsPort_notify_r <= _GEN_5448;
                                                    end
                                                end else begin
                                                    toRegsPort_notify_r <= _GEN_5448;
                                                end
                                            end else begin
                                                toRegsPort_notify_r <= _GEN_5448;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1552) begin
                                                                    if (_T_1793) begin
                                                                        if (io_fromMemoryPort_sync) begin
                                                                            toRegsPort_notify_r <= 1'h0;
                                                                        end else begin
                                                                            toRegsPort_notify_r <= _GEN_5448;
                                                                        end
                                                                    end else begin
                                                                        toRegsPort_notify_r <= _GEN_5448;
                                                                    end
                                                                end else begin
                                                                    toRegsPort_notify_r <= _GEN_5448;
                                                                end
                                                            end else begin
                                                                toRegsPort_notify_r <= _GEN_5448;
                                                            end
                                                        end else begin
                                                            toRegsPort_notify_r <= _GEN_5448;
                                                        end
                                                    end else begin
                                                        toRegsPort_notify_r <= _GEN_5448;
                                                    end
                                                end else begin
                                                    toRegsPort_notify_r <= _GEN_5448;
                                                end
                                            end else begin
                                                toRegsPort_notify_r <= _GEN_5448;
                                            end
                                        end else begin
                                            toRegsPort_notify_r <= _GEN_5448;
                                        end
                                    end
                                end else begin
                                    toRegsPort_notify_r <= _GEN_5848;
                                end
                            end else begin
                                toRegsPort_notify_r <= _GEN_5848;
                            end
                        end else begin
                            toRegsPort_notify_r <= _GEN_5848;
                        end
                    end else begin
                        toRegsPort_notify_r <= _GEN_5848;
                    end
                end else begin
                    toRegsPort_notify_r <= _GEN_5848;
                end
            end else begin
                toRegsPort_notify_r <= _GEN_5848;
            end
        end
        toMemoryPort_r_addrIn <= _GEN_6216[31:0];
        if (reset) begin
            toMemoryPort_r_dataIn <= 32'h0;
        end else begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    toMemoryPort_r_dataIn <= 32'h0;
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1552) begin
                                                                                if (_T_1793) begin
                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                        toMemoryPort_r_dataIn <= 32'h0;
                                                                                    end else begin
                                                                                        if (_T_85) begin
                                                                                            if (_T_337) begin
                                                                                                if (_T_580) begin
                                                                                                    if (_T_823) begin
                                                                                                        if (_T_1066) begin
                                                                                                            if (_T_1309) begin
                                                                                                                if (_T_1550) begin
                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                        toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                    end else begin
                                                                                                                        if (_T_85) begin
                                                                                                                            if (_T_337) begin
                                                                                                                                if (_T_580) begin
                                                                                                                                    if (_T_823) begin
                                                                                                                                        if (_T_1066) begin
                                                                                                                                            if (_T_1307) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_85) begin
                                                                                                                                                        if (_T_337) begin
                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                    if (_T_1064) begin
                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                            toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                        if (_T_821) begin
                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                if (_T_8209) begin
                                                                                                                                                                                                    toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_8217) begin
                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_01;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_8229) begin
                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_02;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_8246) begin
                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_03;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_8268) begin
                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_04;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_8295) begin
                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_05;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_8327) begin
                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_06;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_8364) begin
                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_07;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                if (_T_8406) begin
                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_08;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    if (_T_8453) begin
                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_09;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        if (_T_8505) begin
                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_10;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            if (_T_8562) begin
                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_11;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                if (_T_8624) begin
                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_12;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    if (_T_8691) begin
                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_13;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_8763) begin
                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_14;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_8840) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_15;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_8922) begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_16;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_9009) begin
                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_17;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_9101) begin
                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_18;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_9198) begin
                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_19;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_9300) begin
                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_20;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_9407) begin
                                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_21;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_9519) begin
                                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_22;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_9636) begin
                                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_23;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_9758) begin
                                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_24;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                    if (_T_9885) begin
                                                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_25;
                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                        if (_T_10017) begin
                                                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_26;
                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                            if (_T_10154) begin
                                                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_27;
                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                if (_T_10296) begin
                                                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_28;
                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                    if (_T_10443) begin
                                                                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_29;
                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                        if (_T_10595) begin
                                                                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_30;
                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_31;
                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                                                        if (_T_578) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                                    if (_T_335) begin
                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                                                                        if (_T_823) begin
                                                                                                                                                                                                                                            if (_T_1066) begin
                                                                                                                                                                                                                                                if (_T_1309) begin
                                                                                                                                                                                                                                                    if (_T_1552) begin
                                                                                                                                                                                                                                                        if (_T_1795) begin
                                                                                                                                                                                                                                                            if (_T_2038) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_66) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_47) begin
                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_66) begin
                                                                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_47) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_66) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_46;
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_46;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_46;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_46;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                                                                                    if (_T_1066) begin
                                                                                                                                                                                                                                        if (_T_1309) begin
                                                                                                                                                                                                                                            if (_T_1552) begin
                                                                                                                                                                                                                                                if (_T_1795) begin
                                                                                                                                                                                                                                                    if (_T_2038) begin
                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                if (_T_335) begin
                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_100;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_338;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_338;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_338;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_338;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_338;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                        if (_T_335) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_338;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_338;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_338;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                    if (_T_578) begin
                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                            toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_665;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_665;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_665;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_665;
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                if (_T_578) begin
                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                        toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_665;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_665;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_665;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_665;
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                            if (_T_578) begin
                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                    toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_665;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_665;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_665;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_665;
                                                                                                                                                                                    end
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                            end
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                    if (_T_821) begin
                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                            if (_T_8209) begin
                                                                                                                                                                                                toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_8217) begin
                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_01;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_8229) begin
                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_02;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_8246) begin
                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_03;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_8268) begin
                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_04;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_8295) begin
                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_05;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_8327) begin
                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_06;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_8364) begin
                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_07;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_8406) begin
                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_08;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                if (_T_8453) begin
                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_09;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    if (_T_8505) begin
                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_10;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        if (_T_8562) begin
                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_11;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            if (_T_8624) begin
                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_12;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                if (_T_8691) begin
                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_13;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    if (_T_8763) begin
                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_14;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_8840) begin
                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_15;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_8922) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_16;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_9009) begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_17;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_9101) begin
                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_18;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_9198) begin
                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_19;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_9300) begin
                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_20;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_9407) begin
                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_21;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_9519) begin
                                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_22;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_9636) begin
                                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_23;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_9758) begin
                                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_24;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_9885) begin
                                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_25;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                    if (_T_10017) begin
                                                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_26;
                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                        if (_T_10154) begin
                                                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_27;
                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                            if (_T_10296) begin
                                                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_28;
                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                if (_T_10443) begin
                                                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_29;
                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                    if (_T_10595) begin
                                                                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_30;
                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_31;
                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                        end
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                if (_T_821) begin
                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                        if (_T_8209) begin
                                                                                                                                                                                            toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_8217) begin
                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_01;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_8229) begin
                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_02;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_8246) begin
                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_03;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_8268) begin
                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_04;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_8295) begin
                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_05;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_8327) begin
                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_06;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_8364) begin
                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_07;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_8406) begin
                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_08;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_8453) begin
                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_09;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                if (_T_8505) begin
                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_10;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    if (_T_8562) begin
                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_11;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        if (_T_8624) begin
                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_12;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            if (_T_8691) begin
                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_13;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                if (_T_8763) begin
                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_14;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    if (_T_8840) begin
                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_15;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_8922) begin
                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_16;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_9009) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_17;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_9101) begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_18;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_9198) begin
                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_19;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_9300) begin
                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_20;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_9407) begin
                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_21;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_9519) begin
                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_22;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_9636) begin
                                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_23;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_9758) begin
                                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_24;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_9885) begin
                                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_25;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_10017) begin
                                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_26;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                    if (_T_10154) begin
                                                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_27;
                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                        if (_T_10296) begin
                                                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_28;
                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                            if (_T_10443) begin
                                                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_29;
                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                if (_T_10595) begin
                                                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_30;
                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_31;
                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                    end
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                        if (_T_580) begin
                                                                                                                                                                            if (_T_821) begin
                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                    if (_T_8209) begin
                                                                                                                                                                                        toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_8217) begin
                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_01;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_8229) begin
                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_02;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_8246) begin
                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_03;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_8268) begin
                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_04;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_8295) begin
                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_05;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_8327) begin
                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_06;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_8364) begin
                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_07;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_8406) begin
                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_08;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_8453) begin
                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_09;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_8505) begin
                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_10;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                if (_T_8562) begin
                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_11;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    if (_T_8624) begin
                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_12;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        if (_T_8691) begin
                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_13;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            if (_T_8763) begin
                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_14;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                if (_T_8840) begin
                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_15;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    if (_T_8922) begin
                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_16;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_9009) begin
                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_17;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_9101) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_18;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_9198) begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_19;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_9300) begin
                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_20;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_9407) begin
                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_21;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_9519) begin
                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_22;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_9636) begin
                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_23;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_9758) begin
                                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_24;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_9885) begin
                                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_25;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_10017) begin
                                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_26;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_10154) begin
                                                                                                                                                                                                                                                                                                    toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_27;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                    if (_T_10296) begin
                                                                                                                                                                                                                                                                                                        toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_28;
                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                        if (_T_10443) begin
                                                                                                                                                                                                                                                                                                            toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_29;
                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                            if (_T_10595) begin
                                                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_30;
                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                toMemoryPort_r_dataIn <= io_fromRegsPort_reg_file_31;
                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4160;
                                                                                                                                                                end
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_85) begin
                                                                                                                                                    if (_T_337) begin
                                                                                                                                                        if (_T_580) begin
                                                                                                                                                            if (_T_823) begin
                                                                                                                                                                if (_T_1064) begin
                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                        toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_85) begin
                                                                                                                                                if (_T_337) begin
                                                                                                                                                    if (_T_580) begin
                                                                                                                                                        if (_T_823) begin
                                                                                                                                                            if (_T_1064) begin
                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                    toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_337) begin
                                                                                                                                                if (_T_580) begin
                                                                                                                                                    if (_T_823) begin
                                                                                                                                                        if (_T_1064) begin
                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                                            end else begin
                                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4531;
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                        end
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    if (_T_85) begin
                                                                                                                        if (_T_337) begin
                                                                                                                            if (_T_580) begin
                                                                                                                                if (_T_823) begin
                                                                                                                                    if (_T_1066) begin
                                                                                                                                        if (_T_1307) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                            end else begin
                                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                    end
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1066) begin
                                                                                                                                    if (_T_1307) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                        end else begin
                                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1066) begin
                                                                                                                                if (_T_1307) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                                    end else begin
                                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toMemoryPort_r_dataIn <= _GEN_4845;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                        end
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1309) begin
                                                                                                            if (_T_1550) begin
                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                    toMemoryPort_r_dataIn <= 32'h0;
                                                                                                                end else begin
                                                                                                                    toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                        end
                                                                                    end else begin
                                                                                        toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1309) begin
                                                                                                        if (_T_1550) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                toMemoryPort_r_dataIn <= 32'h0;
                                                                                                            end else begin
                                                                                                                toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                        end
                                                                                    end else begin
                                                                                        toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                    end
                                                                                end else begin
                                                                                    toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1309) begin
                                                                                                    if (_T_1550) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            toMemoryPort_r_dataIn <= 32'h0;
                                                                                                        end else begin
                                                                                                            toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                        end
                                                                                    end else begin
                                                                                        toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                    end
                                                                                end else begin
                                                                                    toMemoryPort_r_dataIn <= _GEN_5033;
                                                                                end
                                                                            end else begin
                                                                                toMemoryPort_r_dataIn <= _GEN_5033;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_r_dataIn <= _GEN_5441;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_r_dataIn <= _GEN_5441;
                                                                end
                                                            end else begin
                                                                toMemoryPort_r_dataIn <= _GEN_5441;
                                                            end
                                                        end else begin
                                                            toMemoryPort_r_dataIn <= _GEN_5441;
                                                        end
                                                    end else begin
                                                        toMemoryPort_r_dataIn <= _GEN_5441;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1552) begin
                                                                            if (_T_1793) begin
                                                                                if (io_fromMemoryPort_sync) begin
                                                                                    toMemoryPort_r_dataIn <= 32'h0;
                                                                                end else begin
                                                                                    toMemoryPort_r_dataIn <= _GEN_5441;
                                                                                end
                                                                            end else begin
                                                                                toMemoryPort_r_dataIn <= _GEN_5441;
                                                                            end
                                                                        end else begin
                                                                            toMemoryPort_r_dataIn <= _GEN_5441;
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_r_dataIn <= _GEN_5441;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_r_dataIn <= _GEN_5441;
                                                                end
                                                            end else begin
                                                                toMemoryPort_r_dataIn <= _GEN_5441;
                                                            end
                                                        end else begin
                                                            toMemoryPort_r_dataIn <= _GEN_5441;
                                                        end
                                                    end else begin
                                                        toMemoryPort_r_dataIn <= _GEN_5441;
                                                    end
                                                end else begin
                                                    toMemoryPort_r_dataIn <= _GEN_5441;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1552) begin
                                                                        if (_T_1793) begin
                                                                            if (io_fromMemoryPort_sync) begin
                                                                                toMemoryPort_r_dataIn <= 32'h0;
                                                                            end else begin
                                                                                toMemoryPort_r_dataIn <= _GEN_5441;
                                                                            end
                                                                        end else begin
                                                                            toMemoryPort_r_dataIn <= _GEN_5441;
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_r_dataIn <= _GEN_5441;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_r_dataIn <= _GEN_5441;
                                                                end
                                                            end else begin
                                                                toMemoryPort_r_dataIn <= _GEN_5441;
                                                            end
                                                        end else begin
                                                            toMemoryPort_r_dataIn <= _GEN_5441;
                                                        end
                                                    end else begin
                                                        toMemoryPort_r_dataIn <= _GEN_5441;
                                                    end
                                                end else begin
                                                    toMemoryPort_r_dataIn <= _GEN_5441;
                                                end
                                            end else begin
                                                toMemoryPort_r_dataIn <= _GEN_5441;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1552) begin
                                                                    if (_T_1793) begin
                                                                        if (io_fromMemoryPort_sync) begin
                                                                            toMemoryPort_r_dataIn <= 32'h0;
                                                                        end else begin
                                                                            toMemoryPort_r_dataIn <= _GEN_5441;
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_r_dataIn <= _GEN_5441;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_r_dataIn <= _GEN_5441;
                                                                end
                                                            end else begin
                                                                toMemoryPort_r_dataIn <= _GEN_5441;
                                                            end
                                                        end else begin
                                                            toMemoryPort_r_dataIn <= _GEN_5441;
                                                        end
                                                    end else begin
                                                        toMemoryPort_r_dataIn <= _GEN_5441;
                                                    end
                                                end else begin
                                                    toMemoryPort_r_dataIn <= _GEN_5441;
                                                end
                                            end else begin
                                                toMemoryPort_r_dataIn <= _GEN_5441;
                                            end
                                        end else begin
                                            toMemoryPort_r_dataIn <= _GEN_5441;
                                        end
                                    end
                                end else begin
                                    toMemoryPort_r_dataIn <= _GEN_5843;
                                end
                            end else begin
                                toMemoryPort_r_dataIn <= _GEN_5843;
                            end
                        end else begin
                            toMemoryPort_r_dataIn <= _GEN_5843;
                        end
                    end else begin
                        toMemoryPort_r_dataIn <= _GEN_5843;
                    end
                end else begin
                    toMemoryPort_r_dataIn <= _GEN_5843;
                end
            end else begin
                toMemoryPort_r_dataIn <= _GEN_5843;
            end
        end
        if (reset) begin
            toMemoryPort_r_mask <= 32'h1;
        end else begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    toMemoryPort_r_mask <= 32'h1;
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1552) begin
                                                                                if (_T_1793) begin
                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                        if (_T_228862) begin
                                                                                            toMemoryPort_r_mask <= 32'h3;
                                                                                        end else begin
                                                                                            if (_T_228877) begin
                                                                                                toMemoryPort_r_mask <= 32'h2;
                                                                                            end else begin
                                                                                                if (_T_228892) begin
                                                                                                    toMemoryPort_r_mask <= 32'h1;
                                                                                                end else begin
                                                                                                    if (_T_228911) begin
                                                                                                        toMemoryPort_r_mask <= 32'h5;
                                                                                                    end else begin
                                                                                                        if (_T_228934) begin
                                                                                                            toMemoryPort_r_mask <= 32'h4;
                                                                                                        end else begin
                                                                                                            toMemoryPort_r_mask <= 32'h0;
                                                                                                        end
                                                                                                    end
                                                                                                end
                                                                                            end
                                                                                        end
                                                                                    end else begin
                                                                                        if (_T_85) begin
                                                                                            if (_T_337) begin
                                                                                                if (_T_580) begin
                                                                                                    if (_T_823) begin
                                                                                                        if (_T_1066) begin
                                                                                                            if (_T_1309) begin
                                                                                                                if (_T_1550) begin
                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                        toMemoryPort_r_mask <= 32'h1;
                                                                                                                    end else begin
                                                                                                                        if (_T_85) begin
                                                                                                                            if (_T_337) begin
                                                                                                                                if (_T_580) begin
                                                                                                                                    if (_T_823) begin
                                                                                                                                        if (_T_1066) begin
                                                                                                                                            if (_T_1307) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_85) begin
                                                                                                                                                        if (_T_337) begin
                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                    if (_T_1064) begin
                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                            toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                        end else begin
                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                        if (_T_821) begin
                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                if (_T_228862) begin
                                                                                                                                                                                                    toMemoryPort_r_mask <= 32'h3;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_228877) begin
                                                                                                                                                                                                        toMemoryPort_r_mask <= 32'h2;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_228892) begin
                                                                                                                                                                                                            toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_228911) begin
                                                                                                                                                                                                                toMemoryPort_r_mask <= 32'h5;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_228934) begin
                                                                                                                                                                                                                    toMemoryPort_r_mask <= 32'h4;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    toMemoryPort_r_mask <= 32'h0;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                                                        if (_T_578) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                                    if (_T_335) begin
                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                            toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                                                                        if (_T_823) begin
                                                                                                                                                                                                                                            if (_T_1066) begin
                                                                                                                                                                                                                                                if (_T_1309) begin
                                                                                                                                                                                                                                                    if (_T_1552) begin
                                                                                                                                                                                                                                                        if (_T_1795) begin
                                                                                                                                                                                                                                                            if (_T_2038) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_66) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_47) begin
                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_66) begin
                                                                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                        toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_47) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_66) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_47;
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_47;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_47;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_47;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                                                                                    if (_T_1066) begin
                                                                                                                                                                                                                                        if (_T_1309) begin
                                                                                                                                                                                                                                            if (_T_1552) begin
                                                                                                                                                                                                                                                if (_T_1795) begin
                                                                                                                                                                                                                                                    if (_T_2038) begin
                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                            toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                if (_T_335) begin
                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                        toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_101;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_339;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_339;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                    toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_339;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_339;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_339;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                        if (_T_335) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_339;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_339;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_339;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                    if (_T_578) begin
                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                            toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_666;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_666;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_666;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_666;
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                if (_T_578) begin
                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                        toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_666;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_666;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_666;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_666;
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                            if (_T_578) begin
                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                    toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_666;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_666;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_666;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_666;
                                                                                                                                                                                    end
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                            end
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                    if (_T_821) begin
                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                            if (_T_228862) begin
                                                                                                                                                                                                toMemoryPort_r_mask <= 32'h3;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_228877) begin
                                                                                                                                                                                                    toMemoryPort_r_mask <= 32'h2;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_228892) begin
                                                                                                                                                                                                        toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_228911) begin
                                                                                                                                                                                                            toMemoryPort_r_mask <= 32'h5;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_228934) begin
                                                                                                                                                                                                                toMemoryPort_r_mask <= 32'h4;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_r_mask <= 32'h0;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                        end
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                if (_T_821) begin
                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                        if (_T_228862) begin
                                                                                                                                                                                            toMemoryPort_r_mask <= 32'h3;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_228877) begin
                                                                                                                                                                                                toMemoryPort_r_mask <= 32'h2;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_228892) begin
                                                                                                                                                                                                    toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_228911) begin
                                                                                                                                                                                                        toMemoryPort_r_mask <= 32'h5;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_228934) begin
                                                                                                                                                                                                            toMemoryPort_r_mask <= 32'h4;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_r_mask <= 32'h0;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                    end
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                        if (_T_580) begin
                                                                                                                                                                            if (_T_821) begin
                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_4325;
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_4161;
                                                                                                                                                                end
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_85) begin
                                                                                                                                                    if (_T_337) begin
                                                                                                                                                        if (_T_580) begin
                                                                                                                                                            if (_T_823) begin
                                                                                                                                                                if (_T_1064) begin
                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                        toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                    end else begin
                                                                                                                                                                        toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_85) begin
                                                                                                                                                if (_T_337) begin
                                                                                                                                                    if (_T_580) begin
                                                                                                                                                        if (_T_823) begin
                                                                                                                                                            if (_T_1064) begin
                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                    toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                                end else begin
                                                                                                                                                                    toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_337) begin
                                                                                                                                                if (_T_580) begin
                                                                                                                                                    if (_T_823) begin
                                                                                                                                                        if (_T_1064) begin
                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                toMemoryPort_r_mask <= 32'h1;
                                                                                                                                                            end else begin
                                                                                                                                                                toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            toMemoryPort_r_mask <= _GEN_4532;
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                        end
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    if (_T_85) begin
                                                                                                                        if (_T_337) begin
                                                                                                                            if (_T_580) begin
                                                                                                                                if (_T_823) begin
                                                                                                                                    if (_T_1066) begin
                                                                                                                                        if (_T_1307) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                toMemoryPort_r_mask <= 32'h1;
                                                                                                                                            end else begin
                                                                                                                                                toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                    end
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1066) begin
                                                                                                                                    if (_T_1307) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            toMemoryPort_r_mask <= 32'h1;
                                                                                                                                        end else begin
                                                                                                                                            toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1066) begin
                                                                                                                                if (_T_1307) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        toMemoryPort_r_mask <= 32'h1;
                                                                                                                                    end else begin
                                                                                                                                        toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toMemoryPort_r_mask <= _GEN_4846;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toMemoryPort_r_mask <= _GEN_4846;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_r_mask <= _GEN_5034;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_r_mask <= _GEN_5034;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_r_mask <= _GEN_5034;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_r_mask <= _GEN_5034;
                                                                                        end
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1309) begin
                                                                                                            if (_T_1550) begin
                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                    toMemoryPort_r_mask <= 32'h1;
                                                                                                                end else begin
                                                                                                                    toMemoryPort_r_mask <= _GEN_5034;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toMemoryPort_r_mask <= _GEN_5034;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            toMemoryPort_r_mask <= _GEN_5034;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_r_mask <= _GEN_5034;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_r_mask <= _GEN_5034;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_r_mask <= _GEN_5034;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_r_mask <= _GEN_5034;
                                                                                        end
                                                                                    end else begin
                                                                                        toMemoryPort_r_mask <= _GEN_5034;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1309) begin
                                                                                                        if (_T_1550) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                toMemoryPort_r_mask <= 32'h1;
                                                                                                            end else begin
                                                                                                                toMemoryPort_r_mask <= _GEN_5034;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            toMemoryPort_r_mask <= _GEN_5034;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_r_mask <= _GEN_5034;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_r_mask <= _GEN_5034;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_r_mask <= _GEN_5034;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_r_mask <= _GEN_5034;
                                                                                        end
                                                                                    end else begin
                                                                                        toMemoryPort_r_mask <= _GEN_5034;
                                                                                    end
                                                                                end else begin
                                                                                    toMemoryPort_r_mask <= _GEN_5034;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1309) begin
                                                                                                    if (_T_1550) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            toMemoryPort_r_mask <= 32'h1;
                                                                                                        end else begin
                                                                                                            toMemoryPort_r_mask <= _GEN_5034;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_r_mask <= _GEN_5034;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_r_mask <= _GEN_5034;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_r_mask <= _GEN_5034;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_r_mask <= _GEN_5034;
                                                                                        end
                                                                                    end else begin
                                                                                        toMemoryPort_r_mask <= _GEN_5034;
                                                                                    end
                                                                                end else begin
                                                                                    toMemoryPort_r_mask <= _GEN_5034;
                                                                                end
                                                                            end else begin
                                                                                toMemoryPort_r_mask <= _GEN_5034;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_r_mask <= _GEN_5442;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_r_mask <= _GEN_5442;
                                                                end
                                                            end else begin
                                                                toMemoryPort_r_mask <= _GEN_5442;
                                                            end
                                                        end else begin
                                                            toMemoryPort_r_mask <= _GEN_5442;
                                                        end
                                                    end else begin
                                                        toMemoryPort_r_mask <= _GEN_5442;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1552) begin
                                                                            if (_T_1793) begin
                                                                                if (io_fromMemoryPort_sync) begin
                                                                                    toMemoryPort_r_mask <= _GEN_4325;
                                                                                end else begin
                                                                                    toMemoryPort_r_mask <= _GEN_5442;
                                                                                end
                                                                            end else begin
                                                                                toMemoryPort_r_mask <= _GEN_5442;
                                                                            end
                                                                        end else begin
                                                                            toMemoryPort_r_mask <= _GEN_5442;
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_r_mask <= _GEN_5442;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_r_mask <= _GEN_5442;
                                                                end
                                                            end else begin
                                                                toMemoryPort_r_mask <= _GEN_5442;
                                                            end
                                                        end else begin
                                                            toMemoryPort_r_mask <= _GEN_5442;
                                                        end
                                                    end else begin
                                                        toMemoryPort_r_mask <= _GEN_5442;
                                                    end
                                                end else begin
                                                    toMemoryPort_r_mask <= _GEN_5442;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1552) begin
                                                                        if (_T_1793) begin
                                                                            if (io_fromMemoryPort_sync) begin
                                                                                toMemoryPort_r_mask <= _GEN_4325;
                                                                            end else begin
                                                                                toMemoryPort_r_mask <= _GEN_5442;
                                                                            end
                                                                        end else begin
                                                                            toMemoryPort_r_mask <= _GEN_5442;
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_r_mask <= _GEN_5442;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_r_mask <= _GEN_5442;
                                                                end
                                                            end else begin
                                                                toMemoryPort_r_mask <= _GEN_5442;
                                                            end
                                                        end else begin
                                                            toMemoryPort_r_mask <= _GEN_5442;
                                                        end
                                                    end else begin
                                                        toMemoryPort_r_mask <= _GEN_5442;
                                                    end
                                                end else begin
                                                    toMemoryPort_r_mask <= _GEN_5442;
                                                end
                                            end else begin
                                                toMemoryPort_r_mask <= _GEN_5442;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1552) begin
                                                                    if (_T_1793) begin
                                                                        if (io_fromMemoryPort_sync) begin
                                                                            toMemoryPort_r_mask <= _GEN_4325;
                                                                        end else begin
                                                                            toMemoryPort_r_mask <= _GEN_5442;
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_r_mask <= _GEN_5442;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_r_mask <= _GEN_5442;
                                                                end
                                                            end else begin
                                                                toMemoryPort_r_mask <= _GEN_5442;
                                                            end
                                                        end else begin
                                                            toMemoryPort_r_mask <= _GEN_5442;
                                                        end
                                                    end else begin
                                                        toMemoryPort_r_mask <= _GEN_5442;
                                                    end
                                                end else begin
                                                    toMemoryPort_r_mask <= _GEN_5442;
                                                end
                                            end else begin
                                                toMemoryPort_r_mask <= _GEN_5442;
                                            end
                                        end else begin
                                            toMemoryPort_r_mask <= _GEN_5442;
                                        end
                                    end
                                end else begin
                                    toMemoryPort_r_mask <= _GEN_5844;
                                end
                            end else begin
                                toMemoryPort_r_mask <= _GEN_5844;
                            end
                        end else begin
                            toMemoryPort_r_mask <= _GEN_5844;
                        end
                    end else begin
                        toMemoryPort_r_mask <= _GEN_5844;
                    end
                end else begin
                    toMemoryPort_r_mask <= _GEN_5844;
                end
            end else begin
                toMemoryPort_r_mask <= _GEN_5844;
            end
        end
        if (reset) begin
            toMemoryPort_r_req <= 32'h1;
        end else begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    toMemoryPort_r_req <= 32'h1;
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1552) begin
                                                                                if (_T_1793) begin
                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                        toMemoryPort_r_req <= 32'h1;
                                                                                    end else begin
                                                                                        if (_T_85) begin
                                                                                            if (_T_337) begin
                                                                                                if (_T_580) begin
                                                                                                    if (_T_823) begin
                                                                                                        if (_T_1066) begin
                                                                                                            if (_T_1309) begin
                                                                                                                if (_T_1550) begin
                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                        toMemoryPort_r_req <= 32'h1;
                                                                                                                    end else begin
                                                                                                                        if (_T_85) begin
                                                                                                                            if (_T_337) begin
                                                                                                                                if (_T_580) begin
                                                                                                                                    if (_T_823) begin
                                                                                                                                        if (_T_1066) begin
                                                                                                                                            if (_T_1307) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    toMemoryPort_r_req <= 32'h1;
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_85) begin
                                                                                                                                                        if (_T_337) begin
                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                    if (_T_1064) begin
                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                            toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                        end else begin
                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                        if (_T_821) begin
                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                toMemoryPort_r_req <= 32'h2;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                                                        if (_T_578) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                                    if (_T_335) begin
                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                            toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                                                                        if (_T_823) begin
                                                                                                                                                                                                                                            if (_T_1066) begin
                                                                                                                                                                                                                                                if (_T_1309) begin
                                                                                                                                                                                                                                                    if (_T_1552) begin
                                                                                                                                                                                                                                                        if (_T_1795) begin
                                                                                                                                                                                                                                                            if (_T_2038) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_66) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_47) begin
                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_66) begin
                                                                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                        toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_47) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_66) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_48;
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_48;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_48;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_48;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                                                                                    if (_T_1066) begin
                                                                                                                                                                                                                                        if (_T_1309) begin
                                                                                                                                                                                                                                            if (_T_1552) begin
                                                                                                                                                                                                                                                if (_T_1795) begin
                                                                                                                                                                                                                                                    if (_T_2038) begin
                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                            toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                if (_T_335) begin
                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                        toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_102;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_340;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_340;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                    toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_340;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_340;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_340;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                        if (_T_335) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_340;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_340;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_340;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                    if (_T_578) begin
                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                            toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_667;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_667;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_667;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_667;
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                if (_T_578) begin
                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                        toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_667;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_667;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_667;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_667;
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                            if (_T_578) begin
                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                    toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_667;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                toMemoryPort_r_req <= _GEN_667;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_667;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_667;
                                                                                                                                                                                    end
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                            end
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                    if (_T_821) begin
                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                            toMemoryPort_r_req <= 32'h2;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                        end
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                if (_T_821) begin
                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                        toMemoryPort_r_req <= 32'h2;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                    end
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                        if (_T_580) begin
                                                                                                                                                                            if (_T_821) begin
                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                    toMemoryPort_r_req <= 32'h2;
                                                                                                                                                                                end else begin
                                                                                                                                                                                    toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    toMemoryPort_r_req <= _GEN_4162;
                                                                                                                                                                end
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_85) begin
                                                                                                                                                    if (_T_337) begin
                                                                                                                                                        if (_T_580) begin
                                                                                                                                                            if (_T_823) begin
                                                                                                                                                                if (_T_1064) begin
                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                        toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                    end else begin
                                                                                                                                                                        toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_85) begin
                                                                                                                                                if (_T_337) begin
                                                                                                                                                    if (_T_580) begin
                                                                                                                                                        if (_T_823) begin
                                                                                                                                                            if (_T_1064) begin
                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                    toMemoryPort_r_req <= 32'h1;
                                                                                                                                                                end else begin
                                                                                                                                                                    toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_337) begin
                                                                                                                                                if (_T_580) begin
                                                                                                                                                    if (_T_823) begin
                                                                                                                                                        if (_T_1064) begin
                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                toMemoryPort_r_req <= 32'h1;
                                                                                                                                                            end else begin
                                                                                                                                                                toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            toMemoryPort_r_req <= _GEN_4533;
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_r_req <= _GEN_4847;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_r_req <= _GEN_4847;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_r_req <= _GEN_4847;
                                                                                                                        end
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    if (_T_85) begin
                                                                                                                        if (_T_337) begin
                                                                                                                            if (_T_580) begin
                                                                                                                                if (_T_823) begin
                                                                                                                                    if (_T_1066) begin
                                                                                                                                        if (_T_1307) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                toMemoryPort_r_req <= 32'h1;
                                                                                                                                            end else begin
                                                                                                                                                toMemoryPort_r_req <= _GEN_4847;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            toMemoryPort_r_req <= _GEN_4847;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        toMemoryPort_r_req <= _GEN_4847;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_r_req <= _GEN_4847;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_r_req <= _GEN_4847;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_r_req <= _GEN_4847;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toMemoryPort_r_req <= _GEN_4847;
                                                                                                                    end
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1066) begin
                                                                                                                                    if (_T_1307) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            toMemoryPort_r_req <= 32'h1;
                                                                                                                                        end else begin
                                                                                                                                            toMemoryPort_r_req <= _GEN_4847;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        toMemoryPort_r_req <= _GEN_4847;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_r_req <= _GEN_4847;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_r_req <= _GEN_4847;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_r_req <= _GEN_4847;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toMemoryPort_r_req <= _GEN_4847;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toMemoryPort_r_req <= _GEN_4847;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1066) begin
                                                                                                                                if (_T_1307) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        toMemoryPort_r_req <= 32'h1;
                                                                                                                                    end else begin
                                                                                                                                        toMemoryPort_r_req <= _GEN_4847;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toMemoryPort_r_req <= _GEN_4847;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toMemoryPort_r_req <= _GEN_4847;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toMemoryPort_r_req <= _GEN_4847;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toMemoryPort_r_req <= _GEN_4847;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toMemoryPort_r_req <= _GEN_4847;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toMemoryPort_r_req <= _GEN_4847;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_r_req <= _GEN_5035;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_r_req <= _GEN_5035;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_r_req <= _GEN_5035;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_r_req <= _GEN_5035;
                                                                                        end
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1309) begin
                                                                                                            if (_T_1550) begin
                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                    toMemoryPort_r_req <= 32'h1;
                                                                                                                end else begin
                                                                                                                    toMemoryPort_r_req <= _GEN_5035;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toMemoryPort_r_req <= _GEN_5035;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            toMemoryPort_r_req <= _GEN_5035;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_r_req <= _GEN_5035;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_r_req <= _GEN_5035;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_r_req <= _GEN_5035;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_r_req <= _GEN_5035;
                                                                                        end
                                                                                    end else begin
                                                                                        toMemoryPort_r_req <= _GEN_5035;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1309) begin
                                                                                                        if (_T_1550) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                toMemoryPort_r_req <= 32'h1;
                                                                                                            end else begin
                                                                                                                toMemoryPort_r_req <= _GEN_5035;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            toMemoryPort_r_req <= _GEN_5035;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_r_req <= _GEN_5035;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_r_req <= _GEN_5035;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_r_req <= _GEN_5035;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_r_req <= _GEN_5035;
                                                                                        end
                                                                                    end else begin
                                                                                        toMemoryPort_r_req <= _GEN_5035;
                                                                                    end
                                                                                end else begin
                                                                                    toMemoryPort_r_req <= _GEN_5035;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1309) begin
                                                                                                    if (_T_1550) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            toMemoryPort_r_req <= 32'h1;
                                                                                                        end else begin
                                                                                                            toMemoryPort_r_req <= _GEN_5035;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toMemoryPort_r_req <= _GEN_5035;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toMemoryPort_r_req <= _GEN_5035;
                                                                                                end
                                                                                            end else begin
                                                                                                toMemoryPort_r_req <= _GEN_5035;
                                                                                            end
                                                                                        end else begin
                                                                                            toMemoryPort_r_req <= _GEN_5035;
                                                                                        end
                                                                                    end else begin
                                                                                        toMemoryPort_r_req <= _GEN_5035;
                                                                                    end
                                                                                end else begin
                                                                                    toMemoryPort_r_req <= _GEN_5035;
                                                                                end
                                                                            end else begin
                                                                                toMemoryPort_r_req <= _GEN_5035;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_r_req <= _GEN_5443;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_r_req <= _GEN_5443;
                                                                end
                                                            end else begin
                                                                toMemoryPort_r_req <= _GEN_5443;
                                                            end
                                                        end else begin
                                                            toMemoryPort_r_req <= _GEN_5443;
                                                        end
                                                    end else begin
                                                        toMemoryPort_r_req <= _GEN_5443;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1552) begin
                                                                            if (_T_1793) begin
                                                                                if (io_fromMemoryPort_sync) begin
                                                                                    toMemoryPort_r_req <= 32'h1;
                                                                                end else begin
                                                                                    toMemoryPort_r_req <= _GEN_5443;
                                                                                end
                                                                            end else begin
                                                                                toMemoryPort_r_req <= _GEN_5443;
                                                                            end
                                                                        end else begin
                                                                            toMemoryPort_r_req <= _GEN_5443;
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_r_req <= _GEN_5443;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_r_req <= _GEN_5443;
                                                                end
                                                            end else begin
                                                                toMemoryPort_r_req <= _GEN_5443;
                                                            end
                                                        end else begin
                                                            toMemoryPort_r_req <= _GEN_5443;
                                                        end
                                                    end else begin
                                                        toMemoryPort_r_req <= _GEN_5443;
                                                    end
                                                end else begin
                                                    toMemoryPort_r_req <= _GEN_5443;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1552) begin
                                                                        if (_T_1793) begin
                                                                            if (io_fromMemoryPort_sync) begin
                                                                                toMemoryPort_r_req <= 32'h1;
                                                                            end else begin
                                                                                toMemoryPort_r_req <= _GEN_5443;
                                                                            end
                                                                        end else begin
                                                                            toMemoryPort_r_req <= _GEN_5443;
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_r_req <= _GEN_5443;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_r_req <= _GEN_5443;
                                                                end
                                                            end else begin
                                                                toMemoryPort_r_req <= _GEN_5443;
                                                            end
                                                        end else begin
                                                            toMemoryPort_r_req <= _GEN_5443;
                                                        end
                                                    end else begin
                                                        toMemoryPort_r_req <= _GEN_5443;
                                                    end
                                                end else begin
                                                    toMemoryPort_r_req <= _GEN_5443;
                                                end
                                            end else begin
                                                toMemoryPort_r_req <= _GEN_5443;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1552) begin
                                                                    if (_T_1793) begin
                                                                        if (io_fromMemoryPort_sync) begin
                                                                            toMemoryPort_r_req <= 32'h1;
                                                                        end else begin
                                                                            toMemoryPort_r_req <= _GEN_5443;
                                                                        end
                                                                    end else begin
                                                                        toMemoryPort_r_req <= _GEN_5443;
                                                                    end
                                                                end else begin
                                                                    toMemoryPort_r_req <= _GEN_5443;
                                                                end
                                                            end else begin
                                                                toMemoryPort_r_req <= _GEN_5443;
                                                            end
                                                        end else begin
                                                            toMemoryPort_r_req <= _GEN_5443;
                                                        end
                                                    end else begin
                                                        toMemoryPort_r_req <= _GEN_5443;
                                                    end
                                                end else begin
                                                    toMemoryPort_r_req <= _GEN_5443;
                                                end
                                            end else begin
                                                toMemoryPort_r_req <= _GEN_5443;
                                            end
                                        end else begin
                                            toMemoryPort_r_req <= _GEN_5443;
                                        end
                                    end
                                end else begin
                                    toMemoryPort_r_req <= _GEN_5845;
                                end
                            end else begin
                                toMemoryPort_r_req <= _GEN_5845;
                            end
                        end else begin
                            toMemoryPort_r_req <= _GEN_5845;
                        end
                    end else begin
                        toMemoryPort_r_req <= _GEN_5845;
                    end
                end else begin
                    toMemoryPort_r_req <= _GEN_5845;
                end
            end else begin
                toMemoryPort_r_req <= _GEN_5845;
            end
        end
        if (!(reset)) begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    if (_T_2328) begin
                                                        toRegsPort_r_dst <= _T_2333;
                                                    end else begin
                                                        toRegsPort_r_dst <= 32'h0;
                                                    end
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1550) begin
                                                                                if (io_fromMemoryPort_sync) begin
                                                                                    if (_T_2328) begin
                                                                                        toRegsPort_r_dst <= _T_2333;
                                                                                    end else begin
                                                                                        toRegsPort_r_dst <= 32'h0;
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1307) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                if (_T_2328) begin
                                                                                                                    toRegsPort_r_dst <= _T_2333;
                                                                                                                end else begin
                                                                                                                    toRegsPort_r_dst <= 32'h0;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1064) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        if (_T_2328) begin
                                                                                                                                            toRegsPort_r_dst <= _T_2333;
                                                                                                                                        end else begin
                                                                                                                                            toRegsPort_r_dst <= 32'h0;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_335) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    toRegsPort_r_dst <= _GEN_352;
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_66) begin
                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                            toRegsPort_r_dst <= regfileWrite_signal_r_dst;
                                                                                                                                                        end
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_66) begin
                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                        toRegsPort_r_dst <= regfileWrite_signal_r_dst;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_66) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    toRegsPort_r_dst <= regfileWrite_signal_r_dst;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    if (_T_85) begin
                                                                                                                                        if (_T_335) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                toRegsPort_r_dst <= _GEN_352;
                                                                                                                                            end else begin
                                                                                                                                                if (_T_66) begin
                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                        toRegsPort_r_dst <= regfileWrite_signal_r_dst;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            toRegsPort_r_dst <= _GEN_103;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        toRegsPort_r_dst <= _GEN_103;
                                                                                                                                    end
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                if (_T_85) begin
                                                                                                                                    if (_T_335) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            toRegsPort_r_dst <= _GEN_352;
                                                                                                                                        end else begin
                                                                                                                                            toRegsPort_r_dst <= _GEN_103;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        toRegsPort_r_dst <= _GEN_103;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toRegsPort_r_dst <= _GEN_103;
                                                                                                                                end
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            if (_T_85) begin
                                                                                                                                if (_T_335) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        toRegsPort_r_dst <= _GEN_352;
                                                                                                                                    end else begin
                                                                                                                                        toRegsPort_r_dst <= _GEN_103;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    toRegsPort_r_dst <= _GEN_103;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toRegsPort_r_dst <= _GEN_103;
                                                                                                                            end
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toRegsPort_r_dst <= _GEN_668;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toRegsPort_r_dst <= _GEN_668;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1064) begin
                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                    toRegsPort_r_dst <= _GEN_352;
                                                                                                                                end else begin
                                                                                                                                    toRegsPort_r_dst <= _GEN_668;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                toRegsPort_r_dst <= _GEN_668;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toRegsPort_r_dst <= _GEN_668;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toRegsPort_r_dst <= _GEN_668;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toRegsPort_r_dst <= _GEN_668;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toRegsPort_r_dst <= _GEN_668;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        if (_T_85) begin
                                                                                                            if (_T_337) begin
                                                                                                                if (_T_580) begin
                                                                                                                    if (_T_823) begin
                                                                                                                        if (_T_1064) begin
                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                toRegsPort_r_dst <= _GEN_352;
                                                                                                                            end else begin
                                                                                                                                toRegsPort_r_dst <= _GEN_668;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            toRegsPort_r_dst <= _GEN_668;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toRegsPort_r_dst <= _GEN_668;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toRegsPort_r_dst <= _GEN_668;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toRegsPort_r_dst <= _GEN_668;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            toRegsPort_r_dst <= _GEN_668;
                                                                                                        end
                                                                                                    end
                                                                                                end else begin
                                                                                                    if (_T_85) begin
                                                                                                        if (_T_337) begin
                                                                                                            if (_T_580) begin
                                                                                                                if (_T_823) begin
                                                                                                                    if (_T_1064) begin
                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                            toRegsPort_r_dst <= _GEN_352;
                                                                                                                        end else begin
                                                                                                                            toRegsPort_r_dst <= _GEN_668;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        toRegsPort_r_dst <= _GEN_668;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    toRegsPort_r_dst <= _GEN_668;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                toRegsPort_r_dst <= _GEN_668;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            toRegsPort_r_dst <= _GEN_668;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toRegsPort_r_dst <= _GEN_668;
                                                                                                    end
                                                                                                end
                                                                                            end else begin
                                                                                                toRegsPort_r_dst <= _GEN_4848;
                                                                                            end
                                                                                        end else begin
                                                                                            toRegsPort_r_dst <= _GEN_4848;
                                                                                        end
                                                                                    end else begin
                                                                                        toRegsPort_r_dst <= _GEN_4848;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1307) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            toRegsPort_r_dst <= _GEN_352;
                                                                                                        end else begin
                                                                                                            toRegsPort_r_dst <= _GEN_4848;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        toRegsPort_r_dst <= _GEN_4848;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toRegsPort_r_dst <= _GEN_4848;
                                                                                                end
                                                                                            end else begin
                                                                                                toRegsPort_r_dst <= _GEN_4848;
                                                                                            end
                                                                                        end else begin
                                                                                            toRegsPort_r_dst <= _GEN_4848;
                                                                                        end
                                                                                    end else begin
                                                                                        toRegsPort_r_dst <= _GEN_4848;
                                                                                    end
                                                                                end else begin
                                                                                    toRegsPort_r_dst <= _GEN_4848;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1307) begin
                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                        toRegsPort_r_dst <= _GEN_352;
                                                                                                    end else begin
                                                                                                        toRegsPort_r_dst <= _GEN_4848;
                                                                                                    end
                                                                                                end else begin
                                                                                                    toRegsPort_r_dst <= _GEN_4848;
                                                                                                end
                                                                                            end else begin
                                                                                                toRegsPort_r_dst <= _GEN_4848;
                                                                                            end
                                                                                        end else begin
                                                                                            toRegsPort_r_dst <= _GEN_4848;
                                                                                        end
                                                                                    end else begin
                                                                                        toRegsPort_r_dst <= _GEN_4848;
                                                                                    end
                                                                                end else begin
                                                                                    toRegsPort_r_dst <= _GEN_4848;
                                                                                end
                                                                            end else begin
                                                                                toRegsPort_r_dst <= _GEN_4848;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        if (_T_85) begin
                                                                            if (_T_337) begin
                                                                                if (_T_580) begin
                                                                                    if (_T_823) begin
                                                                                        if (_T_1066) begin
                                                                                            if (_T_1307) begin
                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                    toRegsPort_r_dst <= _GEN_352;
                                                                                                end else begin
                                                                                                    toRegsPort_r_dst <= _GEN_4848;
                                                                                                end
                                                                                            end else begin
                                                                                                toRegsPort_r_dst <= _GEN_4848;
                                                                                            end
                                                                                        end else begin
                                                                                            toRegsPort_r_dst <= _GEN_4848;
                                                                                        end
                                                                                    end else begin
                                                                                        toRegsPort_r_dst <= _GEN_4848;
                                                                                    end
                                                                                end else begin
                                                                                    toRegsPort_r_dst <= _GEN_4848;
                                                                                end
                                                                            end else begin
                                                                                toRegsPort_r_dst <= _GEN_4848;
                                                                            end
                                                                        end else begin
                                                                            toRegsPort_r_dst <= _GEN_4848;
                                                                        end
                                                                    end
                                                                end else begin
                                                                    toRegsPort_r_dst <= _GEN_5036;
                                                                end
                                                            end else begin
                                                                toRegsPort_r_dst <= _GEN_5036;
                                                            end
                                                        end else begin
                                                            toRegsPort_r_dst <= _GEN_5036;
                                                        end
                                                    end else begin
                                                        toRegsPort_r_dst <= _GEN_5036;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1550) begin
                                                                            if (io_fromMemoryPort_sync) begin
                                                                                toRegsPort_r_dst <= _GEN_352;
                                                                            end else begin
                                                                                toRegsPort_r_dst <= _GEN_5036;
                                                                            end
                                                                        end else begin
                                                                            toRegsPort_r_dst <= _GEN_5036;
                                                                        end
                                                                    end else begin
                                                                        toRegsPort_r_dst <= _GEN_5036;
                                                                    end
                                                                end else begin
                                                                    toRegsPort_r_dst <= _GEN_5036;
                                                                end
                                                            end else begin
                                                                toRegsPort_r_dst <= _GEN_5036;
                                                            end
                                                        end else begin
                                                            toRegsPort_r_dst <= _GEN_5036;
                                                        end
                                                    end else begin
                                                        toRegsPort_r_dst <= _GEN_5036;
                                                    end
                                                end else begin
                                                    toRegsPort_r_dst <= _GEN_5036;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1550) begin
                                                                        if (io_fromMemoryPort_sync) begin
                                                                            toRegsPort_r_dst <= _GEN_352;
                                                                        end else begin
                                                                            toRegsPort_r_dst <= _GEN_5036;
                                                                        end
                                                                    end else begin
                                                                        toRegsPort_r_dst <= _GEN_5036;
                                                                    end
                                                                end else begin
                                                                    toRegsPort_r_dst <= _GEN_5036;
                                                                end
                                                            end else begin
                                                                toRegsPort_r_dst <= _GEN_5036;
                                                            end
                                                        end else begin
                                                            toRegsPort_r_dst <= _GEN_5036;
                                                        end
                                                    end else begin
                                                        toRegsPort_r_dst <= _GEN_5036;
                                                    end
                                                end else begin
                                                    toRegsPort_r_dst <= _GEN_5036;
                                                end
                                            end else begin
                                                toRegsPort_r_dst <= _GEN_5036;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1550) begin
                                                                    if (io_fromMemoryPort_sync) begin
                                                                        toRegsPort_r_dst <= _GEN_352;
                                                                    end else begin
                                                                        toRegsPort_r_dst <= _GEN_5036;
                                                                    end
                                                                end else begin
                                                                    toRegsPort_r_dst <= _GEN_5036;
                                                                end
                                                            end else begin
                                                                toRegsPort_r_dst <= _GEN_5036;
                                                            end
                                                        end else begin
                                                            toRegsPort_r_dst <= _GEN_5036;
                                                        end
                                                    end else begin
                                                        toRegsPort_r_dst <= _GEN_5036;
                                                    end
                                                end else begin
                                                    toRegsPort_r_dst <= _GEN_5036;
                                                end
                                            end else begin
                                                toRegsPort_r_dst <= _GEN_5036;
                                            end
                                        end else begin
                                            toRegsPort_r_dst <= _GEN_5036;
                                        end
                                    end
                                end else begin
                                    toRegsPort_r_dst <= _GEN_5444;
                                end
                            end else begin
                                toRegsPort_r_dst <= _GEN_5444;
                            end
                        end else begin
                            toRegsPort_r_dst <= _GEN_5444;
                        end
                    end else begin
                        toRegsPort_r_dst <= _GEN_5444;
                    end
                end else begin
                    toRegsPort_r_dst <= _GEN_5444;
                end
            end else begin
                toRegsPort_r_dst <= _GEN_5444;
            end
        end
        toRegsPort_r_dstData <= _GEN_6224[31:0];
        memoryAccess_signal_r_addrIn <= _GEN_6209[31:0];
        if (reset) begin
            memoryAccess_signal_r_dataIn <= 32'h0;
        end else begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    memoryAccess_signal_r_dataIn <= 32'h0;
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1552) begin
                                                                                if (_T_1793) begin
                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                        memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                    end else begin
                                                                                        if (_T_85) begin
                                                                                            if (_T_337) begin
                                                                                                if (_T_580) begin
                                                                                                    if (_T_823) begin
                                                                                                        if (_T_1066) begin
                                                                                                            if (_T_1309) begin
                                                                                                                if (_T_1550) begin
                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                        memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                    end else begin
                                                                                                                        if (_T_85) begin
                                                                                                                            if (_T_337) begin
                                                                                                                                if (_T_580) begin
                                                                                                                                    if (_T_823) begin
                                                                                                                                        if (_T_1066) begin
                                                                                                                                            if (_T_1307) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_85) begin
                                                                                                                                                        if (_T_337) begin
                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                    if (_T_1064) begin
                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                            memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                        if (_T_821) begin
                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                if (_T_8209) begin
                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_8217) begin
                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_01;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_8229) begin
                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_02;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_8246) begin
                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_03;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_8268) begin
                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_04;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_8295) begin
                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_05;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_8327) begin
                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_06;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_8364) begin
                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_07;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                if (_T_8406) begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_08;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    if (_T_8453) begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_09;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        if (_T_8505) begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_10;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            if (_T_8562) begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_11;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                if (_T_8624) begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_12;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    if (_T_8691) begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_13;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_8763) begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_14;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_8840) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_15;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_8922) begin
                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_16;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_9009) begin
                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_17;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_9101) begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_18;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_9198) begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_19;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_9300) begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_20;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_9407) begin
                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_21;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_9519) begin
                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_22;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_9636) begin
                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_23;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_9758) begin
                                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_24;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                    if (_T_9885) begin
                                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_25;
                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                        if (_T_10017) begin
                                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_26;
                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                            if (_T_10154) begin
                                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_27;
                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                if (_T_10296) begin
                                                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_28;
                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                    if (_T_10443) begin
                                                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_29;
                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                        if (_T_10595) begin
                                                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_30;
                                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_31;
                                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                                                        if (_T_578) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                                    if (_T_335) begin
                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                                                                        if (_T_823) begin
                                                                                                                                                                                                                                            if (_T_1066) begin
                                                                                                                                                                                                                                                if (_T_1309) begin
                                                                                                                                                                                                                                                    if (_T_1552) begin
                                                                                                                                                                                                                                                        if (_T_1795) begin
                                                                                                                                                                                                                                                            if (_T_2038) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_81) begin
                                                                                                                                                                                                                                                                        if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                            if (_T_66) begin
                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_62) begin
                                                                                                                                                                                                                                                                                        if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                            if (_T_47) begin
                                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_47) begin
                                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_39;
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_39;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_62) begin
                                                                                                                                                                                                                                                                                if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_39;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_39;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_81) begin
                                                                                                                                                                                                                                                                    if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_65;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_65;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_66) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_65;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_65;
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_81) begin
                                                                                                                                                                                                                                                                if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_93;
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_93;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_81) begin
                                                                                                                                                                                                                                                            if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_93;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_93;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                                                                                    if (_T_1066) begin
                                                                                                                                                                                                                                        if (_T_1309) begin
                                                                                                                                                                                                                                            if (_T_1552) begin
                                                                                                                                                                                                                                                if (_T_1795) begin
                                                                                                                                                                                                                                                    if (_T_2038) begin
                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                if (_T_335) begin
                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_121;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_331;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_331;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_331;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_331;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_331;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                        if (_T_335) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_331;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_331;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_331;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                    if (_T_578) begin
                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_658;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_658;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_658;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_658;
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                if (_T_578) begin
                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_658;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_658;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_658;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_658;
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                            if (_T_578) begin
                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_658;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_658;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_658;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_658;
                                                                                                                                                                                    end
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                            end
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                    if (_T_821) begin
                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                            if (_T_8209) begin
                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_8217) begin
                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_01;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_8229) begin
                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_02;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_8246) begin
                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_03;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_8268) begin
                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_04;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_8295) begin
                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_05;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_8327) begin
                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_06;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_8364) begin
                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_07;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_8406) begin
                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_08;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                if (_T_8453) begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_09;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    if (_T_8505) begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_10;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        if (_T_8562) begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_11;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            if (_T_8624) begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_12;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                if (_T_8691) begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_13;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    if (_T_8763) begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_14;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_8840) begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_15;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_8922) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_16;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_9009) begin
                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_17;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_9101) begin
                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_18;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_9198) begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_19;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_9300) begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_20;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_9407) begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_21;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_9519) begin
                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_22;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_9636) begin
                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_23;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_9758) begin
                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_24;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_9885) begin
                                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_25;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                    if (_T_10017) begin
                                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_26;
                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                        if (_T_10154) begin
                                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_27;
                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                            if (_T_10296) begin
                                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_28;
                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                if (_T_10443) begin
                                                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_29;
                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                    if (_T_10595) begin
                                                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_30;
                                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_31;
                                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                        end
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                if (_T_821) begin
                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                        if (_T_8209) begin
                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_8217) begin
                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_01;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_8229) begin
                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_02;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_8246) begin
                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_03;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_8268) begin
                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_04;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_8295) begin
                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_05;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_8327) begin
                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_06;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_8364) begin
                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_07;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_8406) begin
                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_08;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_8453) begin
                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_09;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                if (_T_8505) begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_10;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    if (_T_8562) begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_11;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        if (_T_8624) begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_12;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            if (_T_8691) begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_13;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                if (_T_8763) begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_14;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    if (_T_8840) begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_15;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_8922) begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_16;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_9009) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_17;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_9101) begin
                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_18;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_9198) begin
                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_19;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_9300) begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_20;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_9407) begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_21;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_9519) begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_22;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_9636) begin
                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_23;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_9758) begin
                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_24;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_9885) begin
                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_25;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_10017) begin
                                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_26;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                    if (_T_10154) begin
                                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_27;
                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                        if (_T_10296) begin
                                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_28;
                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                            if (_T_10443) begin
                                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_29;
                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                if (_T_10595) begin
                                                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_30;
                                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_31;
                                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                    end
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                        if (_T_580) begin
                                                                                                                                                                            if (_T_821) begin
                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                    if (_T_8209) begin
                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_8217) begin
                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_01;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_8229) begin
                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_02;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_8246) begin
                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_03;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_8268) begin
                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_04;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_8295) begin
                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_05;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_8327) begin
                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_06;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_8364) begin
                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_07;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_8406) begin
                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_08;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_8453) begin
                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_09;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_8505) begin
                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_10;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                if (_T_8562) begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_11;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    if (_T_8624) begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_12;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        if (_T_8691) begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_13;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            if (_T_8763) begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_14;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                if (_T_8840) begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_15;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    if (_T_8922) begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_16;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_9009) begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_17;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_9101) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_18;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_9198) begin
                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_19;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_9300) begin
                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_20;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_9407) begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_21;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_9519) begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_22;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_9636) begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_23;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_9758) begin
                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_24;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_9885) begin
                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_25;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_10017) begin
                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_26;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_10154) begin
                                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_27;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                    if (_T_10296) begin
                                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_28;
                                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                                        if (_T_10443) begin
                                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_29;
                                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                                            if (_T_10595) begin
                                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_30;
                                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_dataIn <= io_fromRegsPort_reg_file_31;
                                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4153;
                                                                                                                                                                end
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_85) begin
                                                                                                                                                    if (_T_337) begin
                                                                                                                                                        if (_T_580) begin
                                                                                                                                                            if (_T_823) begin
                                                                                                                                                                if (_T_1064) begin
                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                        memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_85) begin
                                                                                                                                                if (_T_337) begin
                                                                                                                                                    if (_T_580) begin
                                                                                                                                                        if (_T_823) begin
                                                                                                                                                            if (_T_1064) begin
                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                    memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_337) begin
                                                                                                                                                if (_T_580) begin
                                                                                                                                                    if (_T_823) begin
                                                                                                                                                        if (_T_1064) begin
                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                                            end else begin
                                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4524;
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                        end
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    if (_T_85) begin
                                                                                                                        if (_T_337) begin
                                                                                                                            if (_T_580) begin
                                                                                                                                if (_T_823) begin
                                                                                                                                    if (_T_1066) begin
                                                                                                                                        if (_T_1307) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                            end else begin
                                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                    end
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1066) begin
                                                                                                                                    if (_T_1307) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                        end else begin
                                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1066) begin
                                                                                                                                if (_T_1307) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                                    end else begin
                                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_4838;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                    end
                                                                                                end else begin
                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                end
                                                                                            end else begin
                                                                                                memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                            end
                                                                                        end else begin
                                                                                            memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                        end
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1309) begin
                                                                                                            if (_T_1550) begin
                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                    memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                                end else begin
                                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                    end
                                                                                                end else begin
                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                end
                                                                                            end else begin
                                                                                                memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                            end
                                                                                        end else begin
                                                                                            memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                        end
                                                                                    end else begin
                                                                                        memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1309) begin
                                                                                                        if (_T_1550) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                            end else begin
                                                                                                                memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                    end
                                                                                                end else begin
                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                end
                                                                                            end else begin
                                                                                                memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                            end
                                                                                        end else begin
                                                                                            memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                        end
                                                                                    end else begin
                                                                                        memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                    end
                                                                                end else begin
                                                                                    memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1309) begin
                                                                                                    if (_T_1550) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                                        end else begin
                                                                                                            memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                    end
                                                                                                end else begin
                                                                                                    memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                                end
                                                                                            end else begin
                                                                                                memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                            end
                                                                                        end else begin
                                                                                            memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                        end
                                                                                    end else begin
                                                                                        memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                    end
                                                                                end else begin
                                                                                    memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                                end
                                                                            end else begin
                                                                                memoryAccess_signal_r_dataIn <= _GEN_5026;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                    end
                                                                end else begin
                                                                    memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                end
                                                            end else begin
                                                                memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                            end
                                                        end else begin
                                                            memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                        end
                                                    end else begin
                                                        memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1552) begin
                                                                            if (_T_1793) begin
                                                                                if (io_fromMemoryPort_sync) begin
                                                                                    memoryAccess_signal_r_dataIn <= 32'h0;
                                                                                end else begin
                                                                                    memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                                end
                                                                            end else begin
                                                                                memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                            end
                                                                        end else begin
                                                                            memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                        end
                                                                    end else begin
                                                                        memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                    end
                                                                end else begin
                                                                    memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                end
                                                            end else begin
                                                                memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                            end
                                                        end else begin
                                                            memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                        end
                                                    end else begin
                                                        memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                    end
                                                end else begin
                                                    memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1552) begin
                                                                        if (_T_1793) begin
                                                                            if (io_fromMemoryPort_sync) begin
                                                                                memoryAccess_signal_r_dataIn <= 32'h0;
                                                                            end else begin
                                                                                memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                            end
                                                                        end else begin
                                                                            memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                        end
                                                                    end else begin
                                                                        memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                    end
                                                                end else begin
                                                                    memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                end
                                                            end else begin
                                                                memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                            end
                                                        end else begin
                                                            memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                        end
                                                    end else begin
                                                        memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                    end
                                                end else begin
                                                    memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                end
                                            end else begin
                                                memoryAccess_signal_r_dataIn <= _GEN_5434;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1552) begin
                                                                    if (_T_1793) begin
                                                                        if (io_fromMemoryPort_sync) begin
                                                                            memoryAccess_signal_r_dataIn <= 32'h0;
                                                                        end else begin
                                                                            memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                        end
                                                                    end else begin
                                                                        memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                    end
                                                                end else begin
                                                                    memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                                end
                                                            end else begin
                                                                memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                            end
                                                        end else begin
                                                            memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                        end
                                                    end else begin
                                                        memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                    end
                                                end else begin
                                                    memoryAccess_signal_r_dataIn <= _GEN_5434;
                                                end
                                            end else begin
                                                memoryAccess_signal_r_dataIn <= _GEN_5434;
                                            end
                                        end else begin
                                            memoryAccess_signal_r_dataIn <= _GEN_5434;
                                        end
                                    end
                                end else begin
                                    memoryAccess_signal_r_dataIn <= _GEN_5836;
                                end
                            end else begin
                                memoryAccess_signal_r_dataIn <= _GEN_5836;
                            end
                        end else begin
                            memoryAccess_signal_r_dataIn <= _GEN_5836;
                        end
                    end else begin
                        memoryAccess_signal_r_dataIn <= _GEN_5836;
                    end
                end else begin
                    memoryAccess_signal_r_dataIn <= _GEN_5836;
                end
            end else begin
                memoryAccess_signal_r_dataIn <= _GEN_5836;
            end
        end
        if (reset) begin
            memoryAccess_signal_r_mask <= 32'h1;
        end else begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    memoryAccess_signal_r_mask <= 32'h1;
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1552) begin
                                                                                if (_T_1793) begin
                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                        if (_T_228862) begin
                                                                                            memoryAccess_signal_r_mask <= 32'h3;
                                                                                        end else begin
                                                                                            if (_T_228877) begin
                                                                                                memoryAccess_signal_r_mask <= 32'h2;
                                                                                            end else begin
                                                                                                if (_T_228892) begin
                                                                                                    memoryAccess_signal_r_mask <= 32'h1;
                                                                                                end else begin
                                                                                                    if (_T_228911) begin
                                                                                                        memoryAccess_signal_r_mask <= 32'h5;
                                                                                                    end else begin
                                                                                                        if (_T_228934) begin
                                                                                                            memoryAccess_signal_r_mask <= 32'h4;
                                                                                                        end else begin
                                                                                                            memoryAccess_signal_r_mask <= 32'h0;
                                                                                                        end
                                                                                                    end
                                                                                                end
                                                                                            end
                                                                                        end
                                                                                    end else begin
                                                                                        if (_T_85) begin
                                                                                            if (_T_337) begin
                                                                                                if (_T_580) begin
                                                                                                    if (_T_823) begin
                                                                                                        if (_T_1066) begin
                                                                                                            if (_T_1309) begin
                                                                                                                if (_T_1550) begin
                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                        memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                    end else begin
                                                                                                                        if (_T_85) begin
                                                                                                                            if (_T_337) begin
                                                                                                                                if (_T_580) begin
                                                                                                                                    if (_T_823) begin
                                                                                                                                        if (_T_1066) begin
                                                                                                                                            if (_T_1307) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_85) begin
                                                                                                                                                        if (_T_337) begin
                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                    if (_T_1064) begin
                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                            memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                        end else begin
                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                        if (_T_821) begin
                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                if (_T_228862) begin
                                                                                                                                                                                                    memoryAccess_signal_r_mask <= 32'h3;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_228877) begin
                                                                                                                                                                                                        memoryAccess_signal_r_mask <= 32'h2;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_228892) begin
                                                                                                                                                                                                            memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_228911) begin
                                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h5;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_228934) begin
                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= 32'h4;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= 32'h0;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                                                        if (_T_578) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                                    if (_T_335) begin
                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                                                                        if (_T_823) begin
                                                                                                                                                                                                                                            if (_T_1066) begin
                                                                                                                                                                                                                                                if (_T_1309) begin
                                                                                                                                                                                                                                                    if (_T_1552) begin
                                                                                                                                                                                                                                                        if (_T_1795) begin
                                                                                                                                                                                                                                                            if (_T_2038) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_81) begin
                                                                                                                                                                                                                                                                        if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                            if (_T_66) begin
                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_62) begin
                                                                                                                                                                                                                                                                                        if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                            if (_T_47) begin
                                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_47) begin
                                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_40;
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_40;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_62) begin
                                                                                                                                                                                                                                                                                if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_40;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_40;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_81) begin
                                                                                                                                                                                                                                                                    if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_66;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_66;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_66) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_66;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_66;
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_81) begin
                                                                                                                                                                                                                                                                if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_94;
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_94;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_81) begin
                                                                                                                                                                                                                                                            if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_94;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_94;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                                                                                    if (_T_1066) begin
                                                                                                                                                                                                                                        if (_T_1309) begin
                                                                                                                                                                                                                                            if (_T_1552) begin
                                                                                                                                                                                                                                                if (_T_1795) begin
                                                                                                                                                                                                                                                    if (_T_2038) begin
                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                if (_T_335) begin
                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                        memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_122;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_332;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_332;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_332;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_332;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_332;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                        if (_T_335) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_332;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_332;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_332;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                    if (_T_578) begin
                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                            memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_659;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_659;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_659;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_659;
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                if (_T_578) begin
                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                        memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_659;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_659;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_659;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_659;
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                            if (_T_578) begin
                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                    memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_659;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_659;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_659;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_659;
                                                                                                                                                                                    end
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                            end
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                    if (_T_821) begin
                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                            if (_T_228862) begin
                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h3;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_228877) begin
                                                                                                                                                                                                    memoryAccess_signal_r_mask <= 32'h2;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_228892) begin
                                                                                                                                                                                                        memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_228911) begin
                                                                                                                                                                                                            memoryAccess_signal_r_mask <= 32'h5;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_228934) begin
                                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h4;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h0;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                        end
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                if (_T_821) begin
                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                        if (_T_228862) begin
                                                                                                                                                                                            memoryAccess_signal_r_mask <= 32'h3;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_228877) begin
                                                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h2;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_228892) begin
                                                                                                                                                                                                    memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_228911) begin
                                                                                                                                                                                                        memoryAccess_signal_r_mask <= 32'h5;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_228934) begin
                                                                                                                                                                                                            memoryAccess_signal_r_mask <= 32'h4;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            memoryAccess_signal_r_mask <= 32'h0;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                    end
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                        if (_T_580) begin
                                                                                                                                                                            if (_T_821) begin
                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4325;
                                                                                                                                                                                end else begin
                                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4154;
                                                                                                                                                                end
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_85) begin
                                                                                                                                                    if (_T_337) begin
                                                                                                                                                        if (_T_580) begin
                                                                                                                                                            if (_T_823) begin
                                                                                                                                                                if (_T_1064) begin
                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                        memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                    end else begin
                                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_85) begin
                                                                                                                                                if (_T_337) begin
                                                                                                                                                    if (_T_580) begin
                                                                                                                                                        if (_T_823) begin
                                                                                                                                                            if (_T_1064) begin
                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                    memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                                end else begin
                                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_337) begin
                                                                                                                                                if (_T_580) begin
                                                                                                                                                    if (_T_823) begin
                                                                                                                                                        if (_T_1064) begin
                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                                            end else begin
                                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4525;
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                        end
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    if (_T_85) begin
                                                                                                                        if (_T_337) begin
                                                                                                                            if (_T_580) begin
                                                                                                                                if (_T_823) begin
                                                                                                                                    if (_T_1066) begin
                                                                                                                                        if (_T_1307) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                            end else begin
                                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                    end
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1066) begin
                                                                                                                                    if (_T_1307) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                        end else begin
                                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1066) begin
                                                                                                                                if (_T_1307) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                                    end else begin
                                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                memoryAccess_signal_r_mask <= _GEN_4839;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                    end
                                                                                                end else begin
                                                                                                    memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                end
                                                                                            end else begin
                                                                                                memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                            end
                                                                                        end else begin
                                                                                            memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                        end
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1309) begin
                                                                                                            if (_T_1550) begin
                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                    memoryAccess_signal_r_mask <= 32'h1;
                                                                                                                end else begin
                                                                                                                    memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                    end
                                                                                                end else begin
                                                                                                    memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                end
                                                                                            end else begin
                                                                                                memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                            end
                                                                                        end else begin
                                                                                            memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                        end
                                                                                    end else begin
                                                                                        memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1309) begin
                                                                                                        if (_T_1550) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                memoryAccess_signal_r_mask <= 32'h1;
                                                                                                            end else begin
                                                                                                                memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                    end
                                                                                                end else begin
                                                                                                    memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                end
                                                                                            end else begin
                                                                                                memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                            end
                                                                                        end else begin
                                                                                            memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                        end
                                                                                    end else begin
                                                                                        memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                    end
                                                                                end else begin
                                                                                    memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1309) begin
                                                                                                    if (_T_1550) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            memoryAccess_signal_r_mask <= 32'h1;
                                                                                                        end else begin
                                                                                                            memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                    end
                                                                                                end else begin
                                                                                                    memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                                end
                                                                                            end else begin
                                                                                                memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                            end
                                                                                        end else begin
                                                                                            memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                        end
                                                                                    end else begin
                                                                                        memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                    end
                                                                                end else begin
                                                                                    memoryAccess_signal_r_mask <= _GEN_5027;
                                                                                end
                                                                            end else begin
                                                                                memoryAccess_signal_r_mask <= _GEN_5027;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        memoryAccess_signal_r_mask <= _GEN_5435;
                                                                    end
                                                                end else begin
                                                                    memoryAccess_signal_r_mask <= _GEN_5435;
                                                                end
                                                            end else begin
                                                                memoryAccess_signal_r_mask <= _GEN_5435;
                                                            end
                                                        end else begin
                                                            memoryAccess_signal_r_mask <= _GEN_5435;
                                                        end
                                                    end else begin
                                                        memoryAccess_signal_r_mask <= _GEN_5435;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1552) begin
                                                                            if (_T_1793) begin
                                                                                if (io_fromMemoryPort_sync) begin
                                                                                    memoryAccess_signal_r_mask <= _GEN_4325;
                                                                                end else begin
                                                                                    memoryAccess_signal_r_mask <= _GEN_5435;
                                                                                end
                                                                            end else begin
                                                                                memoryAccess_signal_r_mask <= _GEN_5435;
                                                                            end
                                                                        end else begin
                                                                            memoryAccess_signal_r_mask <= _GEN_5435;
                                                                        end
                                                                    end else begin
                                                                        memoryAccess_signal_r_mask <= _GEN_5435;
                                                                    end
                                                                end else begin
                                                                    memoryAccess_signal_r_mask <= _GEN_5435;
                                                                end
                                                            end else begin
                                                                memoryAccess_signal_r_mask <= _GEN_5435;
                                                            end
                                                        end else begin
                                                            memoryAccess_signal_r_mask <= _GEN_5435;
                                                        end
                                                    end else begin
                                                        memoryAccess_signal_r_mask <= _GEN_5435;
                                                    end
                                                end else begin
                                                    memoryAccess_signal_r_mask <= _GEN_5435;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1552) begin
                                                                        if (_T_1793) begin
                                                                            if (io_fromMemoryPort_sync) begin
                                                                                memoryAccess_signal_r_mask <= _GEN_4325;
                                                                            end else begin
                                                                                memoryAccess_signal_r_mask <= _GEN_5435;
                                                                            end
                                                                        end else begin
                                                                            memoryAccess_signal_r_mask <= _GEN_5435;
                                                                        end
                                                                    end else begin
                                                                        memoryAccess_signal_r_mask <= _GEN_5435;
                                                                    end
                                                                end else begin
                                                                    memoryAccess_signal_r_mask <= _GEN_5435;
                                                                end
                                                            end else begin
                                                                memoryAccess_signal_r_mask <= _GEN_5435;
                                                            end
                                                        end else begin
                                                            memoryAccess_signal_r_mask <= _GEN_5435;
                                                        end
                                                    end else begin
                                                        memoryAccess_signal_r_mask <= _GEN_5435;
                                                    end
                                                end else begin
                                                    memoryAccess_signal_r_mask <= _GEN_5435;
                                                end
                                            end else begin
                                                memoryAccess_signal_r_mask <= _GEN_5435;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1552) begin
                                                                    if (_T_1793) begin
                                                                        if (io_fromMemoryPort_sync) begin
                                                                            memoryAccess_signal_r_mask <= _GEN_4325;
                                                                        end else begin
                                                                            memoryAccess_signal_r_mask <= _GEN_5435;
                                                                        end
                                                                    end else begin
                                                                        memoryAccess_signal_r_mask <= _GEN_5435;
                                                                    end
                                                                end else begin
                                                                    memoryAccess_signal_r_mask <= _GEN_5435;
                                                                end
                                                            end else begin
                                                                memoryAccess_signal_r_mask <= _GEN_5435;
                                                            end
                                                        end else begin
                                                            memoryAccess_signal_r_mask <= _GEN_5435;
                                                        end
                                                    end else begin
                                                        memoryAccess_signal_r_mask <= _GEN_5435;
                                                    end
                                                end else begin
                                                    memoryAccess_signal_r_mask <= _GEN_5435;
                                                end
                                            end else begin
                                                memoryAccess_signal_r_mask <= _GEN_5435;
                                            end
                                        end else begin
                                            memoryAccess_signal_r_mask <= _GEN_5435;
                                        end
                                    end
                                end else begin
                                    memoryAccess_signal_r_mask <= _GEN_5837;
                                end
                            end else begin
                                memoryAccess_signal_r_mask <= _GEN_5837;
                            end
                        end else begin
                            memoryAccess_signal_r_mask <= _GEN_5837;
                        end
                    end else begin
                        memoryAccess_signal_r_mask <= _GEN_5837;
                    end
                end else begin
                    memoryAccess_signal_r_mask <= _GEN_5837;
                end
            end else begin
                memoryAccess_signal_r_mask <= _GEN_5837;
            end
        end
        if (reset) begin
            memoryAccess_signal_r_req <= 32'h1;
        end else begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    memoryAccess_signal_r_req <= 32'h1;
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1552) begin
                                                                                if (_T_1793) begin
                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                        memoryAccess_signal_r_req <= 32'h1;
                                                                                    end else begin
                                                                                        if (_T_85) begin
                                                                                            if (_T_337) begin
                                                                                                if (_T_580) begin
                                                                                                    if (_T_823) begin
                                                                                                        if (_T_1066) begin
                                                                                                            if (_T_1309) begin
                                                                                                                if (_T_1550) begin
                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                        memoryAccess_signal_r_req <= 32'h1;
                                                                                                                    end else begin
                                                                                                                        if (_T_85) begin
                                                                                                                            if (_T_337) begin
                                                                                                                                if (_T_580) begin
                                                                                                                                    if (_T_823) begin
                                                                                                                                        if (_T_1066) begin
                                                                                                                                            if (_T_1307) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_85) begin
                                                                                                                                                        if (_T_337) begin
                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                    if (_T_1064) begin
                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                            memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                        end else begin
                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                        if (_T_821) begin
                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                memoryAccess_signal_r_req <= 32'h2;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                                                        if (_T_578) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                                    if (_T_335) begin
                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                            memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                                                                        if (_T_823) begin
                                                                                                                                                                                                                                            if (_T_1066) begin
                                                                                                                                                                                                                                                if (_T_1309) begin
                                                                                                                                                                                                                                                    if (_T_1552) begin
                                                                                                                                                                                                                                                        if (_T_1795) begin
                                                                                                                                                                                                                                                            if (_T_2038) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_81) begin
                                                                                                                                                                                                                                                                        if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                            if (_T_66) begin
                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_62) begin
                                                                                                                                                                                                                                                                                        if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                            if (_T_47) begin
                                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_47) begin
                                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_41;
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_41;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_62) begin
                                                                                                                                                                                                                                                                                if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_41;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_41;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_81) begin
                                                                                                                                                                                                                                                                    if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_67;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_67;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_66) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_67;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_67;
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_81) begin
                                                                                                                                                                                                                                                                if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_95;
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_95;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_81) begin
                                                                                                                                                                                                                                                            if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_95;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_95;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                                                                                    if (_T_1066) begin
                                                                                                                                                                                                                                        if (_T_1309) begin
                                                                                                                                                                                                                                            if (_T_1552) begin
                                                                                                                                                                                                                                                if (_T_1795) begin
                                                                                                                                                                                                                                                    if (_T_2038) begin
                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                if (_T_335) begin
                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                        memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_123;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_333;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_333;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                    memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_333;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_333;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_333;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                        if (_T_335) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_333;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_333;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_333;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                    if (_T_578) begin
                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                            memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_660;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_660;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_660;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_660;
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                if (_T_578) begin
                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                        memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_660;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_660;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_660;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_660;
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                            if (_T_578) begin
                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                    memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_660;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_660;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_660;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_660;
                                                                                                                                                                                    end
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                            end
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                    if (_T_821) begin
                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                            memoryAccess_signal_r_req <= 32'h2;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                        end
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                if (_T_821) begin
                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                        memoryAccess_signal_r_req <= 32'h2;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                    end
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                        if (_T_580) begin
                                                                                                                                                                            if (_T_821) begin
                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                    memoryAccess_signal_r_req <= 32'h2;
                                                                                                                                                                                end else begin
                                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4155;
                                                                                                                                                                end
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_85) begin
                                                                                                                                                    if (_T_337) begin
                                                                                                                                                        if (_T_580) begin
                                                                                                                                                            if (_T_823) begin
                                                                                                                                                                if (_T_1064) begin
                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                        memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                    end else begin
                                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_85) begin
                                                                                                                                                if (_T_337) begin
                                                                                                                                                    if (_T_580) begin
                                                                                                                                                        if (_T_823) begin
                                                                                                                                                            if (_T_1064) begin
                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                    memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                                end else begin
                                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_337) begin
                                                                                                                                                if (_T_580) begin
                                                                                                                                                    if (_T_823) begin
                                                                                                                                                        if (_T_1064) begin
                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                                            end else begin
                                                                                                                                                                memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            memoryAccess_signal_r_req <= _GEN_4526;
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                        end
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    if (_T_85) begin
                                                                                                                        if (_T_337) begin
                                                                                                                            if (_T_580) begin
                                                                                                                                if (_T_823) begin
                                                                                                                                    if (_T_1066) begin
                                                                                                                                        if (_T_1307) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                            end else begin
                                                                                                                                                memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                    end
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1066) begin
                                                                                                                                    if (_T_1307) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                        end else begin
                                                                                                                                            memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1066) begin
                                                                                                                                if (_T_1307) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        memoryAccess_signal_r_req <= 32'h1;
                                                                                                                                    end else begin
                                                                                                                                        memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                memoryAccess_signal_r_req <= _GEN_4840;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                    end
                                                                                                end else begin
                                                                                                    memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                end
                                                                                            end else begin
                                                                                                memoryAccess_signal_r_req <= _GEN_5028;
                                                                                            end
                                                                                        end else begin
                                                                                            memoryAccess_signal_r_req <= _GEN_5028;
                                                                                        end
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1309) begin
                                                                                                            if (_T_1550) begin
                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                    memoryAccess_signal_r_req <= 32'h1;
                                                                                                                end else begin
                                                                                                                    memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                    end
                                                                                                end else begin
                                                                                                    memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                end
                                                                                            end else begin
                                                                                                memoryAccess_signal_r_req <= _GEN_5028;
                                                                                            end
                                                                                        end else begin
                                                                                            memoryAccess_signal_r_req <= _GEN_5028;
                                                                                        end
                                                                                    end else begin
                                                                                        memoryAccess_signal_r_req <= _GEN_5028;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1309) begin
                                                                                                        if (_T_1550) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                memoryAccess_signal_r_req <= 32'h1;
                                                                                                            end else begin
                                                                                                                memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                    end
                                                                                                end else begin
                                                                                                    memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                end
                                                                                            end else begin
                                                                                                memoryAccess_signal_r_req <= _GEN_5028;
                                                                                            end
                                                                                        end else begin
                                                                                            memoryAccess_signal_r_req <= _GEN_5028;
                                                                                        end
                                                                                    end else begin
                                                                                        memoryAccess_signal_r_req <= _GEN_5028;
                                                                                    end
                                                                                end else begin
                                                                                    memoryAccess_signal_r_req <= _GEN_5028;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1309) begin
                                                                                                    if (_T_1550) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            memoryAccess_signal_r_req <= 32'h1;
                                                                                                        end else begin
                                                                                                            memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                    end
                                                                                                end else begin
                                                                                                    memoryAccess_signal_r_req <= _GEN_5028;
                                                                                                end
                                                                                            end else begin
                                                                                                memoryAccess_signal_r_req <= _GEN_5028;
                                                                                            end
                                                                                        end else begin
                                                                                            memoryAccess_signal_r_req <= _GEN_5028;
                                                                                        end
                                                                                    end else begin
                                                                                        memoryAccess_signal_r_req <= _GEN_5028;
                                                                                    end
                                                                                end else begin
                                                                                    memoryAccess_signal_r_req <= _GEN_5028;
                                                                                end
                                                                            end else begin
                                                                                memoryAccess_signal_r_req <= _GEN_5028;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        memoryAccess_signal_r_req <= _GEN_5436;
                                                                    end
                                                                end else begin
                                                                    memoryAccess_signal_r_req <= _GEN_5436;
                                                                end
                                                            end else begin
                                                                memoryAccess_signal_r_req <= _GEN_5436;
                                                            end
                                                        end else begin
                                                            memoryAccess_signal_r_req <= _GEN_5436;
                                                        end
                                                    end else begin
                                                        memoryAccess_signal_r_req <= _GEN_5436;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1552) begin
                                                                            if (_T_1793) begin
                                                                                if (io_fromMemoryPort_sync) begin
                                                                                    memoryAccess_signal_r_req <= 32'h1;
                                                                                end else begin
                                                                                    memoryAccess_signal_r_req <= _GEN_5436;
                                                                                end
                                                                            end else begin
                                                                                memoryAccess_signal_r_req <= _GEN_5436;
                                                                            end
                                                                        end else begin
                                                                            memoryAccess_signal_r_req <= _GEN_5436;
                                                                        end
                                                                    end else begin
                                                                        memoryAccess_signal_r_req <= _GEN_5436;
                                                                    end
                                                                end else begin
                                                                    memoryAccess_signal_r_req <= _GEN_5436;
                                                                end
                                                            end else begin
                                                                memoryAccess_signal_r_req <= _GEN_5436;
                                                            end
                                                        end else begin
                                                            memoryAccess_signal_r_req <= _GEN_5436;
                                                        end
                                                    end else begin
                                                        memoryAccess_signal_r_req <= _GEN_5436;
                                                    end
                                                end else begin
                                                    memoryAccess_signal_r_req <= _GEN_5436;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1552) begin
                                                                        if (_T_1793) begin
                                                                            if (io_fromMemoryPort_sync) begin
                                                                                memoryAccess_signal_r_req <= 32'h1;
                                                                            end else begin
                                                                                memoryAccess_signal_r_req <= _GEN_5436;
                                                                            end
                                                                        end else begin
                                                                            memoryAccess_signal_r_req <= _GEN_5436;
                                                                        end
                                                                    end else begin
                                                                        memoryAccess_signal_r_req <= _GEN_5436;
                                                                    end
                                                                end else begin
                                                                    memoryAccess_signal_r_req <= _GEN_5436;
                                                                end
                                                            end else begin
                                                                memoryAccess_signal_r_req <= _GEN_5436;
                                                            end
                                                        end else begin
                                                            memoryAccess_signal_r_req <= _GEN_5436;
                                                        end
                                                    end else begin
                                                        memoryAccess_signal_r_req <= _GEN_5436;
                                                    end
                                                end else begin
                                                    memoryAccess_signal_r_req <= _GEN_5436;
                                                end
                                            end else begin
                                                memoryAccess_signal_r_req <= _GEN_5436;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1552) begin
                                                                    if (_T_1793) begin
                                                                        if (io_fromMemoryPort_sync) begin
                                                                            memoryAccess_signal_r_req <= 32'h1;
                                                                        end else begin
                                                                            memoryAccess_signal_r_req <= _GEN_5436;
                                                                        end
                                                                    end else begin
                                                                        memoryAccess_signal_r_req <= _GEN_5436;
                                                                    end
                                                                end else begin
                                                                    memoryAccess_signal_r_req <= _GEN_5436;
                                                                end
                                                            end else begin
                                                                memoryAccess_signal_r_req <= _GEN_5436;
                                                            end
                                                        end else begin
                                                            memoryAccess_signal_r_req <= _GEN_5436;
                                                        end
                                                    end else begin
                                                        memoryAccess_signal_r_req <= _GEN_5436;
                                                    end
                                                end else begin
                                                    memoryAccess_signal_r_req <= _GEN_5436;
                                                end
                                            end else begin
                                                memoryAccess_signal_r_req <= _GEN_5436;
                                            end
                                        end else begin
                                            memoryAccess_signal_r_req <= _GEN_5436;
                                        end
                                    end
                                end else begin
                                    memoryAccess_signal_r_req <= _GEN_5838;
                                end
                            end else begin
                                memoryAccess_signal_r_req <= _GEN_5838;
                            end
                        end else begin
                            memoryAccess_signal_r_req <= _GEN_5838;
                        end
                    end else begin
                        memoryAccess_signal_r_req <= _GEN_5838;
                    end
                end else begin
                    memoryAccess_signal_r_req <= _GEN_5838;
                end
            end else begin
                memoryAccess_signal_r_req <= _GEN_5838;
            end
        end
        if (reset) begin
            pcReg_signal_r <= 32'h0;
        end else begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    pcReg_signal_r <= _T_223493;
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1552) begin
                                                                                if (_T_1793) begin
                                                                                    if (!(io_fromMemoryPort_sync)) begin
                                                                                        if (_T_85) begin
                                                                                            if (_T_337) begin
                                                                                                if (_T_580) begin
                                                                                                    if (_T_823) begin
                                                                                                        if (_T_1066) begin
                                                                                                            if (_T_1309) begin
                                                                                                                if (_T_1550) begin
                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                        pcReg_signal_r <= _T_50;
                                                                                                                    end else begin
                                                                                                                        if (_T_85) begin
                                                                                                                            if (_T_337) begin
                                                                                                                                if (_T_580) begin
                                                                                                                                    if (_T_823) begin
                                                                                                                                        if (_T_1066) begin
                                                                                                                                            if (_T_1307) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    pcReg_signal_r <= _T_31602;
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_85) begin
                                                                                                                                                        if (_T_337) begin
                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                    if (_T_1064) begin
                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                            pcReg_signal_r <= _T_50;
                                                                                                                                                                        end else begin
                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                        if (_T_821) begin
                                                                                                                                                                                            if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                                                        if (_T_578) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                if (_T_31160) begin
                                                                                                                                                                                                                    pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_36881) begin
                                                                                                                                                                                                                        pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_45243) begin
                                                                                                                                                                                                                            pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_56246) begin
                                                                                                                                                                                                                                pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                if (_T_69890) begin
                                                                                                                                                                                                                                    pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    if (_T_86175) begin
                                                                                                                                                                                                                                        pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        pcReg_signal_r <= _T_86620;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                                    if (_T_335) begin
                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                            pcReg_signal_r <= _T_50;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                                                                        if (_T_823) begin
                                                                                                                                                                                                                                            if (_T_1066) begin
                                                                                                                                                                                                                                                if (_T_1309) begin
                                                                                                                                                                                                                                                    if (_T_1552) begin
                                                                                                                                                                                                                                                        if (_T_1795) begin
                                                                                                                                                                                                                                                            if (_T_2038) begin
                                                                                                                                                                                                                                                                if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                    if (_T_81) begin
                                                                                                                                                                                                                                                                        if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                            if (_T_66) begin
                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    pcReg_signal_r <= _T_50;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_62) begin
                                                                                                                                                                                                                                                                                        if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                            if (_T_47) begin
                                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                    pcReg_signal_r <= _T_50;
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                pcReg_signal_r <= _T_50;
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                pcReg_signal_r <= _T_50;
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_47) begin
                                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                            pcReg_signal_r <= _T_50;
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                pcReg_signal_r <= _T_50;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                        pcReg_signal_r <= _GEN_42;
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_42;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_62) begin
                                                                                                                                                                                                                                                                                if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_42;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_42;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_81) begin
                                                                                                                                                                                                                                                                    if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                pcReg_signal_r <= _T_50;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_68;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_68;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_66) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            pcReg_signal_r <= _T_50;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_68;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        pcReg_signal_r <= _GEN_68;
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_81) begin
                                                                                                                                                                                                                                                                if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_96;
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_96;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_81) begin
                                                                                                                                                                                                                                                            if (!(io_toMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_96;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_96;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                                                                                    if (_T_1066) begin
                                                                                                                                                                                                                                        if (_T_1309) begin
                                                                                                                                                                                                                                            if (_T_1552) begin
                                                                                                                                                                                                                                                if (_T_1795) begin
                                                                                                                                                                                                                                                    if (_T_2038) begin
                                                                                                                                                                                                                                                        if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                if (_T_335) begin
                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                        pcReg_signal_r <= _T_50;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            pcReg_signal_r <= _GEN_124;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_334;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                pcReg_signal_r <= _GEN_334;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                    pcReg_signal_r <= _T_50;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    pcReg_signal_r <= _GEN_334;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                pcReg_signal_r <= _GEN_334;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            pcReg_signal_r <= _GEN_334;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                        if (_T_335) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                pcReg_signal_r <= _T_50;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                pcReg_signal_r <= _GEN_334;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            pcReg_signal_r <= _GEN_334;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        pcReg_signal_r <= _GEN_334;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                    if (_T_578) begin
                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                            if (_T_31160) begin
                                                                                                                                                                                                                pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_36881) begin
                                                                                                                                                                                                                    pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_45243) begin
                                                                                                                                                                                                                        pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_56246) begin
                                                                                                                                                                                                                            pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_69890) begin
                                                                                                                                                                                                                                pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                if (_T_86175) begin
                                                                                                                                                                                                                                    pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    pcReg_signal_r <= _T_86620;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            pcReg_signal_r <= _GEN_661;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        pcReg_signal_r <= _GEN_661;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    pcReg_signal_r <= _GEN_661;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                pcReg_signal_r <= _GEN_661;
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                if (_T_578) begin
                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                        if (_T_31160) begin
                                                                                                                                                                                                            pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_36881) begin
                                                                                                                                                                                                                pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_45243) begin
                                                                                                                                                                                                                    pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_56246) begin
                                                                                                                                                                                                                        pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_69890) begin
                                                                                                                                                                                                                            pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_86175) begin
                                                                                                                                                                                                                                pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                pcReg_signal_r <= _T_86620;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        pcReg_signal_r <= _GEN_661;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    pcReg_signal_r <= _GEN_661;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                pcReg_signal_r <= _GEN_661;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            pcReg_signal_r <= _GEN_661;
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                            if (_T_578) begin
                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                    if (_T_31160) begin
                                                                                                                                                                                                        pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_36881) begin
                                                                                                                                                                                                            pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_45243) begin
                                                                                                                                                                                                                pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_56246) begin
                                                                                                                                                                                                                    pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_69890) begin
                                                                                                                                                                                                                        pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_86175) begin
                                                                                                                                                                                                                            pcReg_signal_r <= _T_31602;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            pcReg_signal_r <= _T_86620;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    pcReg_signal_r <= _GEN_661;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                pcReg_signal_r <= _GEN_661;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            pcReg_signal_r <= _GEN_661;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        pcReg_signal_r <= _GEN_661;
                                                                                                                                                                                    end
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                            end
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                    if (_T_821) begin
                                                                                                                                                                                        if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                            pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                        end
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                if (_T_821) begin
                                                                                                                                                                                    if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                        pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                    end
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                        if (_T_580) begin
                                                                                                                                                                            if (_T_821) begin
                                                                                                                                                                                if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                    pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    pcReg_signal_r <= _GEN_4156;
                                                                                                                                                                end
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            pcReg_signal_r <= _GEN_4527;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        pcReg_signal_r <= _GEN_4527;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_85) begin
                                                                                                                                                    if (_T_337) begin
                                                                                                                                                        if (_T_580) begin
                                                                                                                                                            if (_T_823) begin
                                                                                                                                                                if (_T_1064) begin
                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                        pcReg_signal_r <= _T_50;
                                                                                                                                                                    end else begin
                                                                                                                                                                        pcReg_signal_r <= _GEN_4527;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    pcReg_signal_r <= _GEN_4527;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                pcReg_signal_r <= _GEN_4527;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            pcReg_signal_r <= _GEN_4527;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        pcReg_signal_r <= _GEN_4527;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    pcReg_signal_r <= _GEN_4527;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_85) begin
                                                                                                                                                if (_T_337) begin
                                                                                                                                                    if (_T_580) begin
                                                                                                                                                        if (_T_823) begin
                                                                                                                                                            if (_T_1064) begin
                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                    pcReg_signal_r <= _T_50;
                                                                                                                                                                end else begin
                                                                                                                                                                    pcReg_signal_r <= _GEN_4527;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                pcReg_signal_r <= _GEN_4527;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            pcReg_signal_r <= _GEN_4527;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        pcReg_signal_r <= _GEN_4527;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    pcReg_signal_r <= _GEN_4527;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                pcReg_signal_r <= _GEN_4527;
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_337) begin
                                                                                                                                                if (_T_580) begin
                                                                                                                                                    if (_T_823) begin
                                                                                                                                                        if (_T_1064) begin
                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                pcReg_signal_r <= _T_50;
                                                                                                                                                            end else begin
                                                                                                                                                                pcReg_signal_r <= _GEN_4527;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            pcReg_signal_r <= _GEN_4527;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        pcReg_signal_r <= _GEN_4527;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    pcReg_signal_r <= _GEN_4527;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                pcReg_signal_r <= _GEN_4527;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            pcReg_signal_r <= _GEN_4527;
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    pcReg_signal_r <= _GEN_4841;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                pcReg_signal_r <= _GEN_4841;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            pcReg_signal_r <= _GEN_4841;
                                                                                                                        end
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    if (_T_85) begin
                                                                                                                        if (_T_337) begin
                                                                                                                            if (_T_580) begin
                                                                                                                                if (_T_823) begin
                                                                                                                                    if (_T_1066) begin
                                                                                                                                        if (_T_1307) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                pcReg_signal_r <= _T_31602;
                                                                                                                                            end else begin
                                                                                                                                                pcReg_signal_r <= _GEN_4841;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            pcReg_signal_r <= _GEN_4841;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        pcReg_signal_r <= _GEN_4841;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    pcReg_signal_r <= _GEN_4841;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                pcReg_signal_r <= _GEN_4841;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            pcReg_signal_r <= _GEN_4841;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        pcReg_signal_r <= _GEN_4841;
                                                                                                                    end
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1066) begin
                                                                                                                                    if (_T_1307) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            pcReg_signal_r <= _T_31602;
                                                                                                                                        end else begin
                                                                                                                                            pcReg_signal_r <= _GEN_4841;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        pcReg_signal_r <= _GEN_4841;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    pcReg_signal_r <= _GEN_4841;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                pcReg_signal_r <= _GEN_4841;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            pcReg_signal_r <= _GEN_4841;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        pcReg_signal_r <= _GEN_4841;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    pcReg_signal_r <= _GEN_4841;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1066) begin
                                                                                                                                if (_T_1307) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        pcReg_signal_r <= _T_31602;
                                                                                                                                    end else begin
                                                                                                                                        pcReg_signal_r <= _GEN_4841;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    pcReg_signal_r <= _GEN_4841;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                pcReg_signal_r <= _GEN_4841;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            pcReg_signal_r <= _GEN_4841;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        pcReg_signal_r <= _GEN_4841;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    pcReg_signal_r <= _GEN_4841;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                pcReg_signal_r <= _GEN_4841;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        pcReg_signal_r <= _GEN_5029;
                                                                                                    end
                                                                                                end else begin
                                                                                                    pcReg_signal_r <= _GEN_5029;
                                                                                                end
                                                                                            end else begin
                                                                                                pcReg_signal_r <= _GEN_5029;
                                                                                            end
                                                                                        end else begin
                                                                                            pcReg_signal_r <= _GEN_5029;
                                                                                        end
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1309) begin
                                                                                                            if (_T_1550) begin
                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                    pcReg_signal_r <= _T_50;
                                                                                                                end else begin
                                                                                                                    pcReg_signal_r <= _GEN_5029;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                pcReg_signal_r <= _GEN_5029;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            pcReg_signal_r <= _GEN_5029;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        pcReg_signal_r <= _GEN_5029;
                                                                                                    end
                                                                                                end else begin
                                                                                                    pcReg_signal_r <= _GEN_5029;
                                                                                                end
                                                                                            end else begin
                                                                                                pcReg_signal_r <= _GEN_5029;
                                                                                            end
                                                                                        end else begin
                                                                                            pcReg_signal_r <= _GEN_5029;
                                                                                        end
                                                                                    end else begin
                                                                                        pcReg_signal_r <= _GEN_5029;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1309) begin
                                                                                                        if (_T_1550) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                pcReg_signal_r <= _T_50;
                                                                                                            end else begin
                                                                                                                pcReg_signal_r <= _GEN_5029;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            pcReg_signal_r <= _GEN_5029;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        pcReg_signal_r <= _GEN_5029;
                                                                                                    end
                                                                                                end else begin
                                                                                                    pcReg_signal_r <= _GEN_5029;
                                                                                                end
                                                                                            end else begin
                                                                                                pcReg_signal_r <= _GEN_5029;
                                                                                            end
                                                                                        end else begin
                                                                                            pcReg_signal_r <= _GEN_5029;
                                                                                        end
                                                                                    end else begin
                                                                                        pcReg_signal_r <= _GEN_5029;
                                                                                    end
                                                                                end else begin
                                                                                    pcReg_signal_r <= _GEN_5029;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1309) begin
                                                                                                    if (_T_1550) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            pcReg_signal_r <= _T_50;
                                                                                                        end else begin
                                                                                                            pcReg_signal_r <= _GEN_5029;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        pcReg_signal_r <= _GEN_5029;
                                                                                                    end
                                                                                                end else begin
                                                                                                    pcReg_signal_r <= _GEN_5029;
                                                                                                end
                                                                                            end else begin
                                                                                                pcReg_signal_r <= _GEN_5029;
                                                                                            end
                                                                                        end else begin
                                                                                            pcReg_signal_r <= _GEN_5029;
                                                                                        end
                                                                                    end else begin
                                                                                        pcReg_signal_r <= _GEN_5029;
                                                                                    end
                                                                                end else begin
                                                                                    pcReg_signal_r <= _GEN_5029;
                                                                                end
                                                                            end else begin
                                                                                pcReg_signal_r <= _GEN_5029;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        pcReg_signal_r <= _GEN_5437;
                                                                    end
                                                                end else begin
                                                                    pcReg_signal_r <= _GEN_5437;
                                                                end
                                                            end else begin
                                                                pcReg_signal_r <= _GEN_5437;
                                                            end
                                                        end else begin
                                                            pcReg_signal_r <= _GEN_5437;
                                                        end
                                                    end else begin
                                                        pcReg_signal_r <= _GEN_5437;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1552) begin
                                                                            if (_T_1793) begin
                                                                                if (!(io_fromMemoryPort_sync)) begin
                                                                                    pcReg_signal_r <= _GEN_5437;
                                                                                end
                                                                            end else begin
                                                                                pcReg_signal_r <= _GEN_5437;
                                                                            end
                                                                        end else begin
                                                                            pcReg_signal_r <= _GEN_5437;
                                                                        end
                                                                    end else begin
                                                                        pcReg_signal_r <= _GEN_5437;
                                                                    end
                                                                end else begin
                                                                    pcReg_signal_r <= _GEN_5437;
                                                                end
                                                            end else begin
                                                                pcReg_signal_r <= _GEN_5437;
                                                            end
                                                        end else begin
                                                            pcReg_signal_r <= _GEN_5437;
                                                        end
                                                    end else begin
                                                        pcReg_signal_r <= _GEN_5437;
                                                    end
                                                end else begin
                                                    pcReg_signal_r <= _GEN_5437;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1552) begin
                                                                        if (_T_1793) begin
                                                                            if (!(io_fromMemoryPort_sync)) begin
                                                                                pcReg_signal_r <= _GEN_5437;
                                                                            end
                                                                        end else begin
                                                                            pcReg_signal_r <= _GEN_5437;
                                                                        end
                                                                    end else begin
                                                                        pcReg_signal_r <= _GEN_5437;
                                                                    end
                                                                end else begin
                                                                    pcReg_signal_r <= _GEN_5437;
                                                                end
                                                            end else begin
                                                                pcReg_signal_r <= _GEN_5437;
                                                            end
                                                        end else begin
                                                            pcReg_signal_r <= _GEN_5437;
                                                        end
                                                    end else begin
                                                        pcReg_signal_r <= _GEN_5437;
                                                    end
                                                end else begin
                                                    pcReg_signal_r <= _GEN_5437;
                                                end
                                            end else begin
                                                pcReg_signal_r <= _GEN_5437;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1552) begin
                                                                    if (_T_1793) begin
                                                                        if (!(io_fromMemoryPort_sync)) begin
                                                                            pcReg_signal_r <= _GEN_5437;
                                                                        end
                                                                    end else begin
                                                                        pcReg_signal_r <= _GEN_5437;
                                                                    end
                                                                end else begin
                                                                    pcReg_signal_r <= _GEN_5437;
                                                                end
                                                            end else begin
                                                                pcReg_signal_r <= _GEN_5437;
                                                            end
                                                        end else begin
                                                            pcReg_signal_r <= _GEN_5437;
                                                        end
                                                    end else begin
                                                        pcReg_signal_r <= _GEN_5437;
                                                    end
                                                end else begin
                                                    pcReg_signal_r <= _GEN_5437;
                                                end
                                            end else begin
                                                pcReg_signal_r <= _GEN_5437;
                                            end
                                        end else begin
                                            pcReg_signal_r <= _GEN_5437;
                                        end
                                    end
                                end else begin
                                    pcReg_signal_r <= _GEN_5839;
                                end
                            end else begin
                                pcReg_signal_r <= _GEN_5839;
                            end
                        end else begin
                            pcReg_signal_r <= _GEN_5839;
                        end
                    end else begin
                        pcReg_signal_r <= _GEN_5839;
                    end
                end else begin
                    pcReg_signal_r <= _GEN_5839;
                end
            end else begin
                pcReg_signal_r <= _GEN_5839;
            end
        end
        if (reset) begin
            regfileWrite_signal_r_dst <= 32'h0;
        end else begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    if (_T_2328) begin
                                                        regfileWrite_signal_r_dst <= _T_2333;
                                                    end else begin
                                                        regfileWrite_signal_r_dst <= 32'h0;
                                                    end
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1552) begin
                                                                                if (_T_1793) begin
                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                        if (_T_2328) begin
                                                                                            regfileWrite_signal_r_dst <= _T_2333;
                                                                                        end else begin
                                                                                            regfileWrite_signal_r_dst <= 32'h0;
                                                                                        end
                                                                                    end else begin
                                                                                        if (_T_85) begin
                                                                                            if (_T_337) begin
                                                                                                if (_T_580) begin
                                                                                                    if (_T_823) begin
                                                                                                        if (_T_1066) begin
                                                                                                            if (_T_1309) begin
                                                                                                                if (_T_1550) begin
                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                        if (_T_2328) begin
                                                                                                                            regfileWrite_signal_r_dst <= _T_2333;
                                                                                                                        end else begin
                                                                                                                            regfileWrite_signal_r_dst <= 32'h0;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        if (_T_85) begin
                                                                                                                            if (_T_337) begin
                                                                                                                                if (_T_580) begin
                                                                                                                                    if (_T_823) begin
                                                                                                                                        if (_T_1066) begin
                                                                                                                                            if (_T_1307) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    if (_T_2328) begin
                                                                                                                                                        regfileWrite_signal_r_dst <= _T_2333;
                                                                                                                                                    end else begin
                                                                                                                                                        regfileWrite_signal_r_dst <= 32'h0;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_85) begin
                                                                                                                                                        if (_T_337) begin
                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                    if (_T_1064) begin
                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                                                                                        end else begin
                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                        if (_T_821) begin
                                                                                                                                                                                            if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                                                        if (_T_578) begin
                                                                                                                                                                                                            if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                                    if (_T_335) begin
                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                if (_T_335) begin
                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                        if (_T_335) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                    if (_T_578) begin
                                                                                                                                                                                                        if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_662;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_662;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_662;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_662;
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                if (_T_578) begin
                                                                                                                                                                                                    if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_662;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_662;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_662;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_662;
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                            if (_T_578) begin
                                                                                                                                                                                                if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_662;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_662;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_662;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_662;
                                                                                                                                                                                    end
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                            end
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                    if (_T_821) begin
                                                                                                                                                                                        if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                        end
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                if (_T_821) begin
                                                                                                                                                                                    if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                    end
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                        if (_T_580) begin
                                                                                                                                                                            if (_T_821) begin
                                                                                                                                                                                if (!(io_fromMemoryPort_sync)) begin
                                                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4157;
                                                                                                                                                                end
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_85) begin
                                                                                                                                                    if (_T_337) begin
                                                                                                                                                        if (_T_580) begin
                                                                                                                                                            if (_T_823) begin
                                                                                                                                                                if (_T_1064) begin
                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                                                                                    end else begin
                                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_85) begin
                                                                                                                                                if (_T_337) begin
                                                                                                                                                    if (_T_580) begin
                                                                                                                                                        if (_T_823) begin
                                                                                                                                                            if (_T_1064) begin
                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                                                                                end else begin
                                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_337) begin
                                                                                                                                                if (_T_580) begin
                                                                                                                                                    if (_T_823) begin
                                                                                                                                                        if (_T_1064) begin
                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                                                                            end else begin
                                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4528;
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                        end
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    if (_T_85) begin
                                                                                                                        if (_T_337) begin
                                                                                                                            if (_T_580) begin
                                                                                                                                if (_T_823) begin
                                                                                                                                    if (_T_1066) begin
                                                                                                                                        if (_T_1307) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                                                            end else begin
                                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                    end
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1066) begin
                                                                                                                                    if (_T_1307) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                                                        end else begin
                                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1066) begin
                                                                                                                                if (_T_1307) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                                                    end else begin
                                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                regfileWrite_signal_r_dst <= _GEN_4842;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                    end
                                                                                                end else begin
                                                                                                    regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                end
                                                                                            end else begin
                                                                                                regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                            end
                                                                                        end else begin
                                                                                            regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                        end
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1309) begin
                                                                                                            if (_T_1550) begin
                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                    regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                                end else begin
                                                                                                                    regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                    end
                                                                                                end else begin
                                                                                                    regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                end
                                                                                            end else begin
                                                                                                regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                            end
                                                                                        end else begin
                                                                                            regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                        end
                                                                                    end else begin
                                                                                        regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1309) begin
                                                                                                        if (_T_1550) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                            end else begin
                                                                                                                regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                    end
                                                                                                end else begin
                                                                                                    regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                end
                                                                                            end else begin
                                                                                                regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                            end
                                                                                        end else begin
                                                                                            regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                        end
                                                                                    end else begin
                                                                                        regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                    end
                                                                                end else begin
                                                                                    regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1309) begin
                                                                                                    if (_T_1550) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            regfileWrite_signal_r_dst <= _GEN_352;
                                                                                                        end else begin
                                                                                                            regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                    end
                                                                                                end else begin
                                                                                                    regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                                end
                                                                                            end else begin
                                                                                                regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                            end
                                                                                        end else begin
                                                                                            regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                        end
                                                                                    end else begin
                                                                                        regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                    end
                                                                                end else begin
                                                                                    regfileWrite_signal_r_dst <= _GEN_5030;
                                                                                end
                                                                            end else begin
                                                                                regfileWrite_signal_r_dst <= _GEN_5030;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        regfileWrite_signal_r_dst <= _GEN_5438;
                                                                    end
                                                                end else begin
                                                                    regfileWrite_signal_r_dst <= _GEN_5438;
                                                                end
                                                            end else begin
                                                                regfileWrite_signal_r_dst <= _GEN_5438;
                                                            end
                                                        end else begin
                                                            regfileWrite_signal_r_dst <= _GEN_5438;
                                                        end
                                                    end else begin
                                                        regfileWrite_signal_r_dst <= _GEN_5438;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1552) begin
                                                                            if (_T_1793) begin
                                                                                if (io_fromMemoryPort_sync) begin
                                                                                    regfileWrite_signal_r_dst <= _GEN_352;
                                                                                end else begin
                                                                                    regfileWrite_signal_r_dst <= _GEN_5438;
                                                                                end
                                                                            end else begin
                                                                                regfileWrite_signal_r_dst <= _GEN_5438;
                                                                            end
                                                                        end else begin
                                                                            regfileWrite_signal_r_dst <= _GEN_5438;
                                                                        end
                                                                    end else begin
                                                                        regfileWrite_signal_r_dst <= _GEN_5438;
                                                                    end
                                                                end else begin
                                                                    regfileWrite_signal_r_dst <= _GEN_5438;
                                                                end
                                                            end else begin
                                                                regfileWrite_signal_r_dst <= _GEN_5438;
                                                            end
                                                        end else begin
                                                            regfileWrite_signal_r_dst <= _GEN_5438;
                                                        end
                                                    end else begin
                                                        regfileWrite_signal_r_dst <= _GEN_5438;
                                                    end
                                                end else begin
                                                    regfileWrite_signal_r_dst <= _GEN_5438;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1552) begin
                                                                        if (_T_1793) begin
                                                                            if (io_fromMemoryPort_sync) begin
                                                                                regfileWrite_signal_r_dst <= _GEN_352;
                                                                            end else begin
                                                                                regfileWrite_signal_r_dst <= _GEN_5438;
                                                                            end
                                                                        end else begin
                                                                            regfileWrite_signal_r_dst <= _GEN_5438;
                                                                        end
                                                                    end else begin
                                                                        regfileWrite_signal_r_dst <= _GEN_5438;
                                                                    end
                                                                end else begin
                                                                    regfileWrite_signal_r_dst <= _GEN_5438;
                                                                end
                                                            end else begin
                                                                regfileWrite_signal_r_dst <= _GEN_5438;
                                                            end
                                                        end else begin
                                                            regfileWrite_signal_r_dst <= _GEN_5438;
                                                        end
                                                    end else begin
                                                        regfileWrite_signal_r_dst <= _GEN_5438;
                                                    end
                                                end else begin
                                                    regfileWrite_signal_r_dst <= _GEN_5438;
                                                end
                                            end else begin
                                                regfileWrite_signal_r_dst <= _GEN_5438;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1552) begin
                                                                    if (_T_1793) begin
                                                                        if (io_fromMemoryPort_sync) begin
                                                                            regfileWrite_signal_r_dst <= _GEN_352;
                                                                        end else begin
                                                                            regfileWrite_signal_r_dst <= _GEN_5438;
                                                                        end
                                                                    end else begin
                                                                        regfileWrite_signal_r_dst <= _GEN_5438;
                                                                    end
                                                                end else begin
                                                                    regfileWrite_signal_r_dst <= _GEN_5438;
                                                                end
                                                            end else begin
                                                                regfileWrite_signal_r_dst <= _GEN_5438;
                                                            end
                                                        end else begin
                                                            regfileWrite_signal_r_dst <= _GEN_5438;
                                                        end
                                                    end else begin
                                                        regfileWrite_signal_r_dst <= _GEN_5438;
                                                    end
                                                end else begin
                                                    regfileWrite_signal_r_dst <= _GEN_5438;
                                                end
                                            end else begin
                                                regfileWrite_signal_r_dst <= _GEN_5438;
                                            end
                                        end else begin
                                            regfileWrite_signal_r_dst <= _GEN_5438;
                                        end
                                    end
                                end else begin
                                    regfileWrite_signal_r_dst <= _GEN_5840;
                                end
                            end else begin
                                regfileWrite_signal_r_dst <= _GEN_5840;
                            end
                        end else begin
                            regfileWrite_signal_r_dst <= _GEN_5840;
                        end
                    end else begin
                        regfileWrite_signal_r_dst <= _GEN_5840;
                    end
                end else begin
                    regfileWrite_signal_r_dst <= _GEN_5840;
                end
            end else begin
                regfileWrite_signal_r_dst <= _GEN_5840;
            end
        end
        regfileWrite_signal_r_dstData <= _GEN_6215[31:0];
        if (reset) begin
            state_r <= 3'h4;
        end else begin
            if (_T_85) begin
                if (_T_337) begin
                    if (_T_580) begin
                        if (_T_823) begin
                            if (_T_1066) begin
                                if (_T_1309) begin
                                    if (_T_1552) begin
                                        if (_T_1795) begin
                                            if (_T_2036) begin
                                                if (io_fromMemoryPort_sync) begin
                                                    state_r <= 3'h4;
                                                end else begin
                                                    if (_T_85) begin
                                                        if (_T_337) begin
                                                            if (_T_580) begin
                                                                if (_T_823) begin
                                                                    if (_T_1066) begin
                                                                        if (_T_1309) begin
                                                                            if (_T_1552) begin
                                                                                if (_T_1793) begin
                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                        state_r <= 3'h2;
                                                                                    end else begin
                                                                                        if (_T_85) begin
                                                                                            if (_T_337) begin
                                                                                                if (_T_580) begin
                                                                                                    if (_T_823) begin
                                                                                                        if (_T_1066) begin
                                                                                                            if (_T_1309) begin
                                                                                                                if (_T_1550) begin
                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                        state_r <= 3'h4;
                                                                                                                    end else begin
                                                                                                                        if (_T_85) begin
                                                                                                                            if (_T_337) begin
                                                                                                                                if (_T_580) begin
                                                                                                                                    if (_T_823) begin
                                                                                                                                        if (_T_1066) begin
                                                                                                                                            if (_T_1307) begin
                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                    state_r <= 3'h4;
                                                                                                                                                end else begin
                                                                                                                                                    if (_T_85) begin
                                                                                                                                                        if (_T_337) begin
                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                    if (_T_1064) begin
                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                            state_r <= 3'h4;
                                                                                                                                                                        end else begin
                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                        if (_T_821) begin
                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                state_r <= 3'h0;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                                                        if (_T_578) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                state_r <= 3'h4;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                                                                    if (_T_335) begin
                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                            state_r <= 3'h4;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                                                    if (_T_580) begin
                                                                                                                                                                                                                                        if (_T_823) begin
                                                                                                                                                                                                                                            if (_T_1066) begin
                                                                                                                                                                                                                                                if (_T_1309) begin
                                                                                                                                                                                                                                                    if (_T_1552) begin
                                                                                                                                                                                                                                                        if (_T_1795) begin
                                                                                                                                                                                                                                                            if (_T_2038) begin
                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    state_r <= 3'h4;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_81) begin
                                                                                                                                                                                                                                                                        if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            state_r <= 3'h5;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_66) begin
                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    state_r <= 3'h4;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_62) begin
                                                                                                                                                                                                                                                                                        if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                            state_r <= 3'h3;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_47) begin
                                                                                                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                    state_r <= 3'h4;
                                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                                    if (_T_43) begin
                                                                                                                                                                                                                                                                                                        if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                            state_r <= 3'h1;
                                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_43) begin
                                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                        state_r <= 3'h1;
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                state_r <= 3'h4;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                if (_T_43) begin
                                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                        state_r <= 3'h1;
                                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            if (_T_43) begin
                                                                                                                                                                                                                                                                                                if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                    state_r <= 3'h1;
                                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                        state_r <= 3'h3;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        if (_T_47) begin
                                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                                state_r <= 3'h4;
                                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                                state_r <= _GEN_11;
                                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            state_r <= _GEN_11;
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    if (_T_47) begin
                                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                            state_r <= 3'h4;
                                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                                            state_r <= _GEN_11;
                                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        state_r <= _GEN_11;
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                state_r <= 3'h4;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                if (_T_62) begin
                                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                        state_r <= 3'h3;
                                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                                        state_r <= _GEN_37;
                                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    state_r <= _GEN_37;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            if (_T_62) begin
                                                                                                                                                                                                                                                                                if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                    state_r <= 3'h3;
                                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                                    state_r <= _GEN_37;
                                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                state_r <= _GEN_37;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                if (_T_81) begin
                                                                                                                                                                                                                                                                    if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                        state_r <= 3'h5;
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        if (_T_66) begin
                                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                                state_r <= 3'h4;
                                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                                state_r <= _GEN_63;
                                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            state_r <= _GEN_63;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    if (_T_66) begin
                                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                            state_r <= 3'h4;
                                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                                            state_r <= _GEN_63;
                                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                                        state_r <= _GEN_63;
                                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            if (_T_81) begin
                                                                                                                                                                                                                                                                if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                    state_r <= 3'h5;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                    state_r <= _GEN_91;
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                state_r <= _GEN_91;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        if (_T_81) begin
                                                                                                                                                                                                                                                            if (io_toMemoryPort_sync) begin
                                                                                                                                                                                                                                                                state_r <= 3'h5;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                state_r <= _GEN_91;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            state_r <= _GEN_91;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    state_r <= _GEN_119;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                state_r <= _GEN_119;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            state_r <= _GEN_119;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        state_r <= _GEN_119;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    state_r <= _GEN_119;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                state_r <= _GEN_119;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                state_r <= 3'h4;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                state_r <= _GEN_119;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            state_r <= _GEN_119;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        state_r <= _GEN_119;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    state_r <= _GEN_119;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                state_r <= _GEN_119;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            state_r <= _GEN_119;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        state_r <= _GEN_119;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    state_r <= _GEN_119;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                state_r <= _GEN_119;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            state_r <= _GEN_119;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                                                                if (_T_823) begin
                                                                                                                                                                                                                                    if (_T_1066) begin
                                                                                                                                                                                                                                        if (_T_1309) begin
                                                                                                                                                                                                                                            if (_T_1552) begin
                                                                                                                                                                                                                                                if (_T_1795) begin
                                                                                                                                                                                                                                                    if (_T_2038) begin
                                                                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                            state_r <= 3'h4;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            state_r <= _GEN_119;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        state_r <= _GEN_119;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    state_r <= _GEN_119;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                state_r <= _GEN_119;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            state_r <= _GEN_119;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        state_r <= _GEN_119;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    state_r <= _GEN_119;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                state_r <= _GEN_119;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            state_r <= _GEN_119;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        state_r <= _GEN_119;
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                                if (_T_335) begin
                                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                        state_r <= 3'h4;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                                                                    if (_T_823) begin
                                                                                                                                                                                                                                        if (_T_1066) begin
                                                                                                                                                                                                                                            if (_T_1309) begin
                                                                                                                                                                                                                                                if (_T_1552) begin
                                                                                                                                                                                                                                                    if (_T_1795) begin
                                                                                                                                                                                                                                                        if (_T_2038) begin
                                                                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                                                                state_r <= 3'h4;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                                state_r <= _GEN_119;
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                            state_r <= _GEN_119;
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                        state_r <= _GEN_119;
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                    state_r <= _GEN_119;
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                state_r <= _GEN_119;
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                            state_r <= _GEN_119;
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                        state_r <= _GEN_119;
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                    state_r <= _GEN_119;
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                state_r <= _GEN_119;
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                            state_r <= _GEN_119;
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    state_r <= _GEN_329;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                state_r <= _GEN_329;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                                            if (_T_335) begin
                                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                    state_r <= 3'h4;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                    state_r <= _GEN_329;
                                                                                                                                                                                                                end
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                state_r <= _GEN_329;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            state_r <= _GEN_329;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                                        if (_T_335) begin
                                                                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                                state_r <= 3'h4;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                state_r <= _GEN_329;
                                                                                                                                                                                                            end
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            state_r <= _GEN_329;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        state_r <= _GEN_329;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            if (_T_85) begin
                                                                                                                                                                                                if (_T_337) begin
                                                                                                                                                                                                    if (_T_578) begin
                                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                            state_r <= 3'h4;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                            state_r <= _GEN_656;
                                                                                                                                                                                                        end
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        state_r <= _GEN_656;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    state_r <= _GEN_656;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                state_r <= _GEN_656;
                                                                                                                                                                                            end
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                                if (_T_578) begin
                                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                        state_r <= 3'h4;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                        state_r <= _GEN_656;
                                                                                                                                                                                                    end
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    state_r <= _GEN_656;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                state_r <= _GEN_656;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            state_r <= _GEN_656;
                                                                                                                                                                                        end
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                                            if (_T_578) begin
                                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                                    state_r <= 3'h4;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                    state_r <= _GEN_656;
                                                                                                                                                                                                end
                                                                                                                                                                                            end else begin
                                                                                                                                                                                                state_r <= _GEN_656;
                                                                                                                                                                                            end
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            state_r <= _GEN_656;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        state_r <= _GEN_656;
                                                                                                                                                                                    end
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                state_r <= _GEN_4151;
                                                                                                                                                                            end
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        if (_T_85) begin
                                                                                                                                                                            if (_T_337) begin
                                                                                                                                                                                if (_T_580) begin
                                                                                                                                                                                    if (_T_821) begin
                                                                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                            state_r <= 3'h0;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                            state_r <= _GEN_4151;
                                                                                                                                                                                        end
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        state_r <= _GEN_4151;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    state_r <= _GEN_4151;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                state_r <= _GEN_4151;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            state_r <= _GEN_4151;
                                                                                                                                                                        end
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    if (_T_85) begin
                                                                                                                                                                        if (_T_337) begin
                                                                                                                                                                            if (_T_580) begin
                                                                                                                                                                                if (_T_821) begin
                                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                        state_r <= 3'h0;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                        state_r <= _GEN_4151;
                                                                                                                                                                                    end
                                                                                                                                                                                end else begin
                                                                                                                                                                                    state_r <= _GEN_4151;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                state_r <= _GEN_4151;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            state_r <= _GEN_4151;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        state_r <= _GEN_4151;
                                                                                                                                                                    end
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                if (_T_85) begin
                                                                                                                                                                    if (_T_337) begin
                                                                                                                                                                        if (_T_580) begin
                                                                                                                                                                            if (_T_821) begin
                                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                                    state_r <= 3'h0;
                                                                                                                                                                                end else begin
                                                                                                                                                                                    state_r <= _GEN_4151;
                                                                                                                                                                                end
                                                                                                                                                                            end else begin
                                                                                                                                                                                state_r <= _GEN_4151;
                                                                                                                                                                            end
                                                                                                                                                                        end else begin
                                                                                                                                                                            state_r <= _GEN_4151;
                                                                                                                                                                        end
                                                                                                                                                                    end else begin
                                                                                                                                                                        state_r <= _GEN_4151;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    state_r <= _GEN_4151;
                                                                                                                                                                end
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            state_r <= _GEN_4522;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        state_r <= _GEN_4522;
                                                                                                                                                    end
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                if (_T_85) begin
                                                                                                                                                    if (_T_337) begin
                                                                                                                                                        if (_T_580) begin
                                                                                                                                                            if (_T_823) begin
                                                                                                                                                                if (_T_1064) begin
                                                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                                                        state_r <= 3'h4;
                                                                                                                                                                    end else begin
                                                                                                                                                                        state_r <= _GEN_4522;
                                                                                                                                                                    end
                                                                                                                                                                end else begin
                                                                                                                                                                    state_r <= _GEN_4522;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                state_r <= _GEN_4522;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            state_r <= _GEN_4522;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        state_r <= _GEN_4522;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    state_r <= _GEN_4522;
                                                                                                                                                end
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            if (_T_85) begin
                                                                                                                                                if (_T_337) begin
                                                                                                                                                    if (_T_580) begin
                                                                                                                                                        if (_T_823) begin
                                                                                                                                                            if (_T_1064) begin
                                                                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                                                                    state_r <= 3'h4;
                                                                                                                                                                end else begin
                                                                                                                                                                    state_r <= _GEN_4522;
                                                                                                                                                                end
                                                                                                                                                            end else begin
                                                                                                                                                                state_r <= _GEN_4522;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            state_r <= _GEN_4522;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        state_r <= _GEN_4522;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    state_r <= _GEN_4522;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                state_r <= _GEN_4522;
                                                                                                                                            end
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        if (_T_85) begin
                                                                                                                                            if (_T_337) begin
                                                                                                                                                if (_T_580) begin
                                                                                                                                                    if (_T_823) begin
                                                                                                                                                        if (_T_1064) begin
                                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                                state_r <= 3'h4;
                                                                                                                                                            end else begin
                                                                                                                                                                state_r <= _GEN_4522;
                                                                                                                                                            end
                                                                                                                                                        end else begin
                                                                                                                                                            state_r <= _GEN_4522;
                                                                                                                                                        end
                                                                                                                                                    end else begin
                                                                                                                                                        state_r <= _GEN_4522;
                                                                                                                                                    end
                                                                                                                                                end else begin
                                                                                                                                                    state_r <= _GEN_4522;
                                                                                                                                                end
                                                                                                                                            end else begin
                                                                                                                                                state_r <= _GEN_4522;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            state_r <= _GEN_4522;
                                                                                                                                        end
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    state_r <= _GEN_4836;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                state_r <= _GEN_4836;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            state_r <= _GEN_4836;
                                                                                                                        end
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    if (_T_85) begin
                                                                                                                        if (_T_337) begin
                                                                                                                            if (_T_580) begin
                                                                                                                                if (_T_823) begin
                                                                                                                                    if (_T_1066) begin
                                                                                                                                        if (_T_1307) begin
                                                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                                                state_r <= 3'h4;
                                                                                                                                            end else begin
                                                                                                                                                state_r <= _GEN_4836;
                                                                                                                                            end
                                                                                                                                        end else begin
                                                                                                                                            state_r <= _GEN_4836;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        state_r <= _GEN_4836;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    state_r <= _GEN_4836;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                state_r <= _GEN_4836;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            state_r <= _GEN_4836;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        state_r <= _GEN_4836;
                                                                                                                    end
                                                                                                                end
                                                                                                            end else begin
                                                                                                                if (_T_85) begin
                                                                                                                    if (_T_337) begin
                                                                                                                        if (_T_580) begin
                                                                                                                            if (_T_823) begin
                                                                                                                                if (_T_1066) begin
                                                                                                                                    if (_T_1307) begin
                                                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                                                            state_r <= 3'h4;
                                                                                                                                        end else begin
                                                                                                                                            state_r <= _GEN_4836;
                                                                                                                                        end
                                                                                                                                    end else begin
                                                                                                                                        state_r <= _GEN_4836;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    state_r <= _GEN_4836;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                state_r <= _GEN_4836;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            state_r <= _GEN_4836;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        state_r <= _GEN_4836;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    state_r <= _GEN_4836;
                                                                                                                end
                                                                                                            end
                                                                                                        end else begin
                                                                                                            if (_T_85) begin
                                                                                                                if (_T_337) begin
                                                                                                                    if (_T_580) begin
                                                                                                                        if (_T_823) begin
                                                                                                                            if (_T_1066) begin
                                                                                                                                if (_T_1307) begin
                                                                                                                                    if (io_fromMemoryPort_sync) begin
                                                                                                                                        state_r <= 3'h4;
                                                                                                                                    end else begin
                                                                                                                                        state_r <= _GEN_4836;
                                                                                                                                    end
                                                                                                                                end else begin
                                                                                                                                    state_r <= _GEN_4836;
                                                                                                                                end
                                                                                                                            end else begin
                                                                                                                                state_r <= _GEN_4836;
                                                                                                                            end
                                                                                                                        end else begin
                                                                                                                            state_r <= _GEN_4836;
                                                                                                                        end
                                                                                                                    end else begin
                                                                                                                        state_r <= _GEN_4836;
                                                                                                                    end
                                                                                                                end else begin
                                                                                                                    state_r <= _GEN_4836;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                state_r <= _GEN_4836;
                                                                                                            end
                                                                                                        end
                                                                                                    end else begin
                                                                                                        state_r <= _GEN_5024;
                                                                                                    end
                                                                                                end else begin
                                                                                                    state_r <= _GEN_5024;
                                                                                                end
                                                                                            end else begin
                                                                                                state_r <= _GEN_5024;
                                                                                            end
                                                                                        end else begin
                                                                                            state_r <= _GEN_5024;
                                                                                        end
                                                                                    end
                                                                                end else begin
                                                                                    if (_T_85) begin
                                                                                        if (_T_337) begin
                                                                                            if (_T_580) begin
                                                                                                if (_T_823) begin
                                                                                                    if (_T_1066) begin
                                                                                                        if (_T_1309) begin
                                                                                                            if (_T_1550) begin
                                                                                                                if (io_fromMemoryPort_sync) begin
                                                                                                                    state_r <= 3'h4;
                                                                                                                end else begin
                                                                                                                    state_r <= _GEN_5024;
                                                                                                                end
                                                                                                            end else begin
                                                                                                                state_r <= _GEN_5024;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            state_r <= _GEN_5024;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        state_r <= _GEN_5024;
                                                                                                    end
                                                                                                end else begin
                                                                                                    state_r <= _GEN_5024;
                                                                                                end
                                                                                            end else begin
                                                                                                state_r <= _GEN_5024;
                                                                                            end
                                                                                        end else begin
                                                                                            state_r <= _GEN_5024;
                                                                                        end
                                                                                    end else begin
                                                                                        state_r <= _GEN_5024;
                                                                                    end
                                                                                end
                                                                            end else begin
                                                                                if (_T_85) begin
                                                                                    if (_T_337) begin
                                                                                        if (_T_580) begin
                                                                                            if (_T_823) begin
                                                                                                if (_T_1066) begin
                                                                                                    if (_T_1309) begin
                                                                                                        if (_T_1550) begin
                                                                                                            if (io_fromMemoryPort_sync) begin
                                                                                                                state_r <= 3'h4;
                                                                                                            end else begin
                                                                                                                state_r <= _GEN_5024;
                                                                                                            end
                                                                                                        end else begin
                                                                                                            state_r <= _GEN_5024;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        state_r <= _GEN_5024;
                                                                                                    end
                                                                                                end else begin
                                                                                                    state_r <= _GEN_5024;
                                                                                                end
                                                                                            end else begin
                                                                                                state_r <= _GEN_5024;
                                                                                            end
                                                                                        end else begin
                                                                                            state_r <= _GEN_5024;
                                                                                        end
                                                                                    end else begin
                                                                                        state_r <= _GEN_5024;
                                                                                    end
                                                                                end else begin
                                                                                    state_r <= _GEN_5024;
                                                                                end
                                                                            end
                                                                        end else begin
                                                                            if (_T_85) begin
                                                                                if (_T_337) begin
                                                                                    if (_T_580) begin
                                                                                        if (_T_823) begin
                                                                                            if (_T_1066) begin
                                                                                                if (_T_1309) begin
                                                                                                    if (_T_1550) begin
                                                                                                        if (io_fromMemoryPort_sync) begin
                                                                                                            state_r <= 3'h4;
                                                                                                        end else begin
                                                                                                            state_r <= _GEN_5024;
                                                                                                        end
                                                                                                    end else begin
                                                                                                        state_r <= _GEN_5024;
                                                                                                    end
                                                                                                end else begin
                                                                                                    state_r <= _GEN_5024;
                                                                                                end
                                                                                            end else begin
                                                                                                state_r <= _GEN_5024;
                                                                                            end
                                                                                        end else begin
                                                                                            state_r <= _GEN_5024;
                                                                                        end
                                                                                    end else begin
                                                                                        state_r <= _GEN_5024;
                                                                                    end
                                                                                end else begin
                                                                                    state_r <= _GEN_5024;
                                                                                end
                                                                            end else begin
                                                                                state_r <= _GEN_5024;
                                                                            end
                                                                        end
                                                                    end else begin
                                                                        state_r <= _GEN_5432;
                                                                    end
                                                                end else begin
                                                                    state_r <= _GEN_5432;
                                                                end
                                                            end else begin
                                                                state_r <= _GEN_5432;
                                                            end
                                                        end else begin
                                                            state_r <= _GEN_5432;
                                                        end
                                                    end else begin
                                                        state_r <= _GEN_5432;
                                                    end
                                                end
                                            end else begin
                                                if (_T_85) begin
                                                    if (_T_337) begin
                                                        if (_T_580) begin
                                                            if (_T_823) begin
                                                                if (_T_1066) begin
                                                                    if (_T_1309) begin
                                                                        if (_T_1552) begin
                                                                            if (_T_1793) begin
                                                                                if (io_fromMemoryPort_sync) begin
                                                                                    state_r <= 3'h2;
                                                                                end else begin
                                                                                    state_r <= _GEN_5432;
                                                                                end
                                                                            end else begin
                                                                                state_r <= _GEN_5432;
                                                                            end
                                                                        end else begin
                                                                            state_r <= _GEN_5432;
                                                                        end
                                                                    end else begin
                                                                        state_r <= _GEN_5432;
                                                                    end
                                                                end else begin
                                                                    state_r <= _GEN_5432;
                                                                end
                                                            end else begin
                                                                state_r <= _GEN_5432;
                                                            end
                                                        end else begin
                                                            state_r <= _GEN_5432;
                                                        end
                                                    end else begin
                                                        state_r <= _GEN_5432;
                                                    end
                                                end else begin
                                                    state_r <= _GEN_5432;
                                                end
                                            end
                                        end else begin
                                            if (_T_85) begin
                                                if (_T_337) begin
                                                    if (_T_580) begin
                                                        if (_T_823) begin
                                                            if (_T_1066) begin
                                                                if (_T_1309) begin
                                                                    if (_T_1552) begin
                                                                        if (_T_1793) begin
                                                                            if (io_fromMemoryPort_sync) begin
                                                                                state_r <= 3'h2;
                                                                            end else begin
                                                                                state_r <= _GEN_5432;
                                                                            end
                                                                        end else begin
                                                                            state_r <= _GEN_5432;
                                                                        end
                                                                    end else begin
                                                                        state_r <= _GEN_5432;
                                                                    end
                                                                end else begin
                                                                    state_r <= _GEN_5432;
                                                                end
                                                            end else begin
                                                                state_r <= _GEN_5432;
                                                            end
                                                        end else begin
                                                            state_r <= _GEN_5432;
                                                        end
                                                    end else begin
                                                        state_r <= _GEN_5432;
                                                    end
                                                end else begin
                                                    state_r <= _GEN_5432;
                                                end
                                            end else begin
                                                state_r <= _GEN_5432;
                                            end
                                        end
                                    end else begin
                                        if (_T_85) begin
                                            if (_T_337) begin
                                                if (_T_580) begin
                                                    if (_T_823) begin
                                                        if (_T_1066) begin
                                                            if (_T_1309) begin
                                                                if (_T_1552) begin
                                                                    if (_T_1793) begin
                                                                        if (io_fromMemoryPort_sync) begin
                                                                            state_r <= 3'h2;
                                                                        end else begin
                                                                            state_r <= _GEN_5432;
                                                                        end
                                                                    end else begin
                                                                        state_r <= _GEN_5432;
                                                                    end
                                                                end else begin
                                                                    state_r <= _GEN_5432;
                                                                end
                                                            end else begin
                                                                state_r <= _GEN_5432;
                                                            end
                                                        end else begin
                                                            state_r <= _GEN_5432;
                                                        end
                                                    end else begin
                                                        state_r <= _GEN_5432;
                                                    end
                                                end else begin
                                                    state_r <= _GEN_5432;
                                                end
                                            end else begin
                                                state_r <= _GEN_5432;
                                            end
                                        end else begin
                                            state_r <= _GEN_5432;
                                        end
                                    end
                                end else begin
                                    state_r <= _GEN_5834;
                                end
                            end else begin
                                state_r <= _GEN_5834;
                            end
                        end else begin
                            state_r <= _GEN_5834;
                        end
                    end else begin
                        state_r <= _GEN_5834;
                    end
                end else begin
                    state_r <= _GEN_5834;
                end
            end else begin
                state_r <= _GEN_5834;
            end
        end
    end
endmodule
