library ieee;
use IEEE.numeric_std.all;

package TestBasic6_types is
end package TestBasic6_types;