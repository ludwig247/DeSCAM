library ieee;
use IEEE.numeric_std.all;

package TestBasic14_types is
type TestBasic14_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic14_types;
