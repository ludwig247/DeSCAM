library ieee;
use IEEE.numeric_std.all;
use work.SCAM_Model_types.all;

package TestMasterSlave5_types is
type Sections is (SECTION_A, SECTION_B);
end package TestMasterSlave5_types;