package testbasic9_types;

endpackage