library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave1_types is
type TestMasterSlave1_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave1_types;
