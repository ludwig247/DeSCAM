library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestArray2_types is
end package TestArray2_types;