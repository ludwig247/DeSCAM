library ieee;
use IEEE.numeric_std.all;

package TestBasic3_types is
end package TestBasic3_types;