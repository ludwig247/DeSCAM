package testarray3_types;

	import scam_model_types::*;
endpackage