package testbasic0_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic0_SECTIONS;

endpackage
