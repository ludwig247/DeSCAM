package testbasic6_types;

	import scam_model_types::*;
endpackage