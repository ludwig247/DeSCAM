package testmasterslave3_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave3_SECTIONS;

endpackage
