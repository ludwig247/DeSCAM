package testbasic4_types;

	typedef enum logic {
		run
	} TestBasic4_SECTIONS;

endpackage
