package testmasterslave10_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave10_SECTIONS;

endpackage
