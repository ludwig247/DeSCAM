library ieee;
use IEEE.numeric_std.all;
use work.SCAM_Model_types.all;

package TestBasic7_types is
end package TestBasic7_types;