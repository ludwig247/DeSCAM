package testbasic6_types;

	typedef enum logic {
		run
	} TestBasic6_SECTIONS;

endpackage
