-- External data type definition package
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package SCAM_Model_types is
	type ME_MaskType is (MT_B, MT_BU, MT_H, MT_HU, MT_W, MT_X);
	type ME_AccessType is (ME_RD, ME_WR, ME_X);
	type CUtoME_IF is record
		addrIn: unsigned(31 downto 0);
		dataIn: unsigned(31 downto 0);
		mask: ME_MaskType;
		req: ME_AccessType;
	end record;
	type AccessType_Reg is (REG_RD, REG_WR);
	type CtlToRegs_IF is record
		dst: unsigned(31 downto 0);
		dst_data: unsigned(31 downto 0);
		req: AccessType_Reg;
		src1: unsigned(31 downto 0);
		src2: unsigned(31 downto 0);
	end record;
	type EncType is (B, Error_Type, I, J, R, S, U);
	type InstrType is (And_Instr, Or_Instr, Unknown, Xor_Instr, add, addI, andI, auipc, beq, bge, bgeu, blt, bltu, bne, jal, jalr, lb, lbu, lh, lhu, lui, lw, orI, sb, sh, sllI, sll_Instr, slt, sltI, sltIu, sltu, sraI, sra_Instr, srlI, srl_Instr, sub, sw, xorI);
	type DecodedInstr is record
		encType: EncType;
		imm: unsigned(31 downto 0);
		instrType: InstrType;
		rd_addr: unsigned(31 downto 0);
		rs1_addr: unsigned(31 downto 0);
		rs2_addr: unsigned(31 downto 0);
	end record;
	type MEtoCU_IF is record
		loadedData: unsigned(31 downto 0);
	end record;
	type RegsToCtl_IF is record
		contents1: unsigned(31 downto 0);
		contents2: unsigned(31 downto 0);
	end record;
end package SCAM_Model_types;



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.SCAM_Model_types.all;

entity ISA is
port(	
	CtlToDec_port_sig: out unsigned(31 downto 0);
	CtlToDec_port_notify: out boolean;
	CtlToMem_port_sig: out CUtoME_IF;
	CtlToMem_port_sync: in boolean;
	CtlToMem_port_notify: out boolean;
	CtlToRegs_port_sig: out CtlToRegs_IF;
	CtlToRegs_port_notify: out boolean;
	DecToCtl_port_sig: in DecodedInstr;
	MemToCtl_port_sig: in MEtoCU_IF;
	MemToCtl_port_sync: in boolean;
	MemToCtl_port_notify: out boolean;
	RegsToCtl_port_sig: in RegsToCtl_IF;
	dummy_port_sig: in boolean;
	clk: in std_logic;
	rst: in std_logic
);
end ISA;

architecture ISA_arch of ISA is
	-- Define internal data types
	type ISA_operation_t is (op_wait_fetch_4, op_fetch_4_write_97, op_wait_fetch_5, op_fetch_5_read_98, op_fetch_5_read_99, op_fetch_5_read_100, op_fetch_5_read_101, op_fetch_5_read_102, op_fetch_5_read_103, op_fetch_5_read_104, op_fetch_5_read_105, op_fetch_5_read_106, op_fetch_5_read_107, op_fetch_5_read_108, op_fetch_5_read_109, op_fetch_5_read_110, op_fetch_5_read_111, op_fetch_5_read_112, op_fetch_5_read_113, op_fetch_5_read_114, op_fetch_5_read_115, op_fetch_5_read_116, op_fetch_5_read_117, op_fetch_5_read_118, op_fetch_5_read_119, op_fetch_5_read_120, op_fetch_5_read_121, op_fetch_5_read_122, op_fetch_5_read_123, op_fetch_5_read_124, op_fetch_5_read_125, op_fetch_5_read_126, op_fetch_5_read_127, op_fetch_5_read_128, op_fetch_5_read_129, op_fetch_5_read_130, op_fetch_5_read_131, op_fetch_5_read_132, op_fetch_5_read_133, op_fetch_5_read_134, op_fetch_5_read_135, op_fetch_5_read_136, op_fetch_5_read_137, op_fetch_5_read_138, op_fetch_5_read_139, op_fetch_5_read_140, op_fetch_5_read_141, op_fetch_5_read_142, op_fetch_5_read_143, op_fetch_5_read_144, op_fetch_5_read_145, op_fetch_5_read_146, op_fetch_5_read_147, op_fetch_5_read_148, op_fetch_5_read_149, op_fetch_5_read_150, op_fetch_5_read_151, op_fetch_5_read_152, op_fetch_5_read_153, op_fetch_5_read_154, op_fetch_5_read_155, op_fetch_5_read_156, op_fetch_5_read_157, op_fetch_5_read_158, op_fetch_5_read_159, op_fetch_5_read_160, op_fetch_5_read_161, op_fetch_5_read_162, op_fetch_5_read_163, op_fetch_5_read_164, op_fetch_5_read_165, op_fetch_5_read_166, op_fetch_5_read_167, op_fetch_5_read_168, op_fetch_5_read_169, op_fetch_5_read_170, op_fetch_5_read_171, op_fetch_5_read_172, op_fetch_5_read_173, op_fetch_5_read_174, op_fetch_5_read_175, op_fetch_5_read_176, op_fetch_5_read_177, op_fetch_5_read_178, op_fetch_5_read_179, op_fetch_5_read_180, op_fetch_5_read_181, op_fetch_5_read_182, op_fetch_5_read_183, op_fetch_5_read_184, op_fetch_5_read_185, op_fetch_5_read_186, op_fetch_5_read_187, op_fetch_5_read_188, op_fetch_5_read_189, op_fetch_5_read_190, op_fetch_5_read_191, op_fetch_5_read_192, op_fetch_5_read_193, op_fetch_5_read_194, op_fetch_5_read_195, op_fetch_5_read_196, op_fetch_5_read_197, op_fetch_5_read_198, op_fetch_5_read_199, op_fetch_5_read_200, op_fetch_5_read_201, op_fetch_5_read_202, op_fetch_5_read_203, op_fetch_5_read_204, op_fetch_5_read_205, op_fetch_5_read_206, op_fetch_5_read_207, op_fetch_5_read_208, op_fetch_5_read_209, op_fetch_5_read_210, op_fetch_5_read_211, op_fetch_5_read_212, op_fetch_5_read_213, op_fetch_5_read_214, op_fetch_5_read_215, op_fetch_5_read_216, op_fetch_5_read_217, op_fetch_5_read_218, op_fetch_5_read_219, op_fetch_5_read_220, op_fetch_5_read_221, op_fetch_5_read_222, op_fetch_5_read_223, op_fetch_5_read_224, op_fetch_5_read_225, op_fetch_5_read_226, op_fetch_5_read_227, op_fetch_5_read_228, op_fetch_5_read_229, op_fetch_5_read_230, op_fetch_5_read_231, op_fetch_5_read_232, op_fetch_5_read_233, op_fetch_5_read_234, op_fetch_5_read_235, op_fetch_5_read_236, op_fetch_5_read_237, op_fetch_5_read_238, op_fetch_5_read_239, op_fetch_5_read_240, op_fetch_5_read_241, op_fetch_5_read_242, op_fetch_5_read_243, op_fetch_5_read_244, op_fetch_5_read_245, op_fetch_5_read_246, op_fetch_5_read_247, op_fetch_5_read_248, op_fetch_5_read_249, op_fetch_5_read_250, op_fetch_5_read_251, op_fetch_5_read_252, op_fetch_5_read_253, op_fetch_5_read_254, op_fetch_5_read_255, op_fetch_5_read_256, op_fetch_5_read_257, op_fetch_5_read_258, op_fetch_5_read_259, op_fetch_5_read_260, op_fetch_5_read_261, op_fetch_5_read_262, op_fetch_5_read_263, op_fetch_5_read_264, op_fetch_5_read_265, op_fetch_5_read_266, op_fetch_5_read_267, op_fetch_5_read_268, op_fetch_5_read_269, op_fetch_5_read_270, op_fetch_5_read_271, op_fetch_5_read_272, op_fetch_5_read_273, op_fetch_5_read_274, op_fetch_5_read_275, op_fetch_5_read_276, op_fetch_5_read_277, op_fetch_5_read_278, op_fetch_5_read_279, op_fetch_5_read_280, op_fetch_5_read_281, op_fetch_5_read_282, op_fetch_5_read_283, op_fetch_5_read_284, op_fetch_5_read_285, op_fetch_5_read_286, op_fetch_5_read_287, op_fetch_5_read_288, op_fetch_5_read_289, op_fetch_5_read_290, op_fetch_5_read_291, op_fetch_5_read_292, op_fetch_5_read_293, op_fetch_5_read_294, op_fetch_5_read_295, op_fetch_5_read_296, op_fetch_5_read_297, op_fetch_5_read_298, op_fetch_5_read_299, op_fetch_5_read_300, op_fetch_5_read_301, op_fetch_5_read_302, op_fetch_5_read_303, op_fetch_5_read_304, op_fetch_5_read_305, op_fetch_5_read_306, op_fetch_5_read_307, op_fetch_5_read_308, op_fetch_5_read_309, op_fetch_5_read_310, op_fetch_5_read_311, op_fetch_5_read_312, op_fetch_5_read_313, op_fetch_5_read_314, op_fetch_5_read_315, op_fetch_5_read_316, op_fetch_5_read_317, op_fetch_5_read_318, op_fetch_5_read_319, op_fetch_5_read_320, op_fetch_5_read_321, op_fetch_5_read_322, op_fetch_5_read_323, op_fetch_5_read_324, op_fetch_5_read_325, op_fetch_5_read_326, op_fetch_5_read_327, op_fetch_5_read_328, op_fetch_5_read_329, op_fetch_5_read_330, op_fetch_5_read_331, op_fetch_5_read_332, op_fetch_5_read_333, op_fetch_5_read_334, op_fetch_5_read_335, op_fetch_5_read_336, op_fetch_5_read_337, op_fetch_5_read_338, op_fetch_5_read_339, op_fetch_5_read_340, op_fetch_5_read_341, op_fetch_5_read_342, op_fetch_5_read_343, op_fetch_5_read_344, op_fetch_5_read_345, op_fetch_5_read_346, op_fetch_5_read_347, op_fetch_5_read_348, op_fetch_5_read_349, op_fetch_5_read_350, op_fetch_5_read_351, op_fetch_5_read_352, op_fetch_5_read_353, op_fetch_5_read_354, op_fetch_5_read_355, op_fetch_5_read_356, op_fetch_5_read_357, op_fetch_5_read_358, op_fetch_5_read_359, op_fetch_5_read_360, op_fetch_5_read_361, op_fetch_5_read_362, op_fetch_5_read_363, op_fetch_5_read_364, op_fetch_5_read_365, op_fetch_5_read_366, op_fetch_5_read_367, op_fetch_5_read_368, op_fetch_5_read_369, op_fetch_5_read_370, op_fetch_5_read_371, op_fetch_5_read_372, op_fetch_5_read_373, op_fetch_5_read_374, op_fetch_5_read_375, op_fetch_5_read_376, op_fetch_5_read_377, op_fetch_5_read_378, op_fetch_5_read_379, op_fetch_5_read_380, op_fetch_5_read_381, op_fetch_5_read_382, op_fetch_5_read_383, op_fetch_5_read_384, op_fetch_5_read_385, op_fetch_5_read_386, op_fetch_5_read_387, op_fetch_5_read_388, op_fetch_5_read_389, op_fetch_5_read_390, op_fetch_5_read_391, op_fetch_5_read_392, op_fetch_5_read_393, op_fetch_5_read_394, op_fetch_5_read_395, op_fetch_5_read_396, op_fetch_5_read_397, op_fetch_5_read_398, op_fetch_5_read_399, op_fetch_5_read_400, op_fetch_5_read_401, op_fetch_5_read_402, op_fetch_5_read_403, op_fetch_5_read_404, op_fetch_5_read_405, op_fetch_5_read_406, op_fetch_5_read_407, op_fetch_5_read_408, op_fetch_5_read_409, op_fetch_5_read_410, op_fetch_5_read_411, op_fetch_5_read_412, op_fetch_5_read_413, op_fetch_5_read_414, op_fetch_5_read_415, op_fetch_5_read_416, op_fetch_5_read_417, op_fetch_5_read_418, op_fetch_5_read_419, op_fetch_5_read_420, op_fetch_5_read_421, op_fetch_5_read_422, op_fetch_5_read_423, op_fetch_5_read_424, op_fetch_5_read_425, op_fetch_5_read_426, op_fetch_5_read_427, op_fetch_5_read_428, op_fetch_5_read_429, op_fetch_5_read_430, op_fetch_5_read_431, op_fetch_5_read_432, op_fetch_5_read_433, op_fetch_5_read_434, op_fetch_5_read_435, op_fetch_5_read_436, op_fetch_5_read_437, op_fetch_5_read_438, op_fetch_5_read_439, op_fetch_5_read_440, op_fetch_5_read_441, op_fetch_5_read_442, op_fetch_5_read_443, op_fetch_5_read_444, op_fetch_5_read_445, op_fetch_5_read_446, op_fetch_5_read_447, op_fetch_5_read_448, op_fetch_5_read_449, op_fetch_5_read_450, op_fetch_5_read_451, op_fetch_5_read_452, op_fetch_5_read_453, op_fetch_5_read_454, op_fetch_5_read_455, op_fetch_5_read_456, op_fetch_5_read_457, op_fetch_5_read_458, op_fetch_5_read_459, op_fetch_5_read_460, op_fetch_5_read_461, op_fetch_5_read_462, op_fetch_5_read_463, op_fetch_5_read_464, op_fetch_5_read_465, op_fetch_5_read_466, op_fetch_5_read_467, op_fetch_5_read_468, op_fetch_5_read_469, op_fetch_5_read_470, op_fetch_5_read_471, op_fetch_5_read_472, op_fetch_5_read_473, op_fetch_5_read_474, op_fetch_5_read_475, op_fetch_5_read_476, op_fetch_5_read_477, op_fetch_5_read_478, op_fetch_5_read_479, op_fetch_5_read_480, op_fetch_5_read_481, op_fetch_5_read_482, op_fetch_5_read_483, op_fetch_5_read_484, op_fetch_5_read_485, op_fetch_5_read_486, op_fetch_5_read_487, op_fetch_5_read_488, op_fetch_5_read_489, op_fetch_5_read_490, op_fetch_5_read_491, op_fetch_5_read_492, op_fetch_5_read_493, op_fetch_5_read_494, op_fetch_5_read_495, op_fetch_5_read_496, op_fetch_5_read_497, op_fetch_5_read_498, op_fetch_5_read_499, op_fetch_5_read_500, op_fetch_5_read_501, op_fetch_5_read_502, op_fetch_5_read_503, op_fetch_5_read_504, op_fetch_5_read_505, op_fetch_5_read_506, op_fetch_5_read_507, op_fetch_5_read_508, op_fetch_5_read_509, op_fetch_5_read_510, op_fetch_5_read_511, op_fetch_5_read_512, op_fetch_5_read_513, op_fetch_5_read_514, op_fetch_5_read_515, op_fetch_5_read_516, op_fetch_5_read_517, op_fetch_5_read_518, op_fetch_5_read_519, op_fetch_5_read_520, op_fetch_5_read_521, op_fetch_5_read_522, op_fetch_5_read_523, op_fetch_5_read_524, op_fetch_5_read_525, op_fetch_5_read_526, op_fetch_5_read_527, op_fetch_5_read_528, op_fetch_5_read_529, op_fetch_5_read_530, op_fetch_5_read_531, op_fetch_5_read_532, op_fetch_5_read_533, op_fetch_5_read_534, op_fetch_5_read_535, op_fetch_5_read_536, op_fetch_5_read_537, op_fetch_5_read_538, op_fetch_5_read_539, op_fetch_5_read_540, op_fetch_5_read_541, op_fetch_5_read_542, op_fetch_5_read_543, op_fetch_5_read_544, op_fetch_5_read_545, op_fetch_5_read_546, op_fetch_5_read_547, op_fetch_5_read_548, op_fetch_5_read_549, op_fetch_5_read_550, op_fetch_5_read_551, op_fetch_5_read_552, op_fetch_5_read_553, op_fetch_5_read_554, op_fetch_5_read_555, op_fetch_5_read_556, op_fetch_5_read_557, op_fetch_5_read_558, op_fetch_5_read_559, op_fetch_5_read_560, op_fetch_5_read_561, op_fetch_5_read_562, op_fetch_5_read_563, op_fetch_5_read_564, op_fetch_5_read_565, op_fetch_5_read_566, op_fetch_5_read_567, op_fetch_5_read_568, op_fetch_5_read_569, op_fetch_5_read_570, op_fetch_5_read_571, op_fetch_5_read_572, op_fetch_5_read_573, op_fetch_5_read_574, op_fetch_5_read_575, op_fetch_5_read_576, op_fetch_5_read_577, op_fetch_5_read_578, op_fetch_5_read_579, op_fetch_5_read_580, op_fetch_5_read_581, op_fetch_5_read_582, op_fetch_5_read_583, op_fetch_5_read_584, op_fetch_5_read_585, op_fetch_5_read_586, op_fetch_5_read_587, op_fetch_5_read_588, op_fetch_5_read_589, op_fetch_5_read_590, op_fetch_5_read_591, op_fetch_5_read_592, op_fetch_5_read_593, op_fetch_5_read_594, op_fetch_5_read_595, op_fetch_5_read_596, op_fetch_5_read_597, op_fetch_5_read_598, op_fetch_5_read_599, op_fetch_5_read_600, op_fetch_5_read_601, op_fetch_5_read_602, op_fetch_5_read_603, op_fetch_5_read_604, op_fetch_5_read_605, op_fetch_5_read_606, op_fetch_5_read_607, op_fetch_5_read_608, op_fetch_5_read_609, op_fetch_5_read_610, op_fetch_5_read_611, op_fetch_5_read_612, op_fetch_5_read_613, op_fetch_5_read_614, op_fetch_5_read_615, op_fetch_5_read_616, op_fetch_5_read_617, op_fetch_5_read_618, op_fetch_5_read_619, op_fetch_5_read_620, op_fetch_5_read_621, op_fetch_5_read_622, op_fetch_5_read_623, op_fetch_5_read_624, op_fetch_5_read_625, op_fetch_5_read_626, op_fetch_5_read_627, op_fetch_5_read_628, op_fetch_5_read_629, op_fetch_5_read_630, op_fetch_5_read_631, op_fetch_5_read_632, op_fetch_5_read_633, op_fetch_5_read_634, op_fetch_5_read_635, op_fetch_5_read_636, op_fetch_5_read_637, op_fetch_5_read_638, op_fetch_5_read_639, op_fetch_5_read_640, op_fetch_5_read_641, op_fetch_5_read_642, op_fetch_5_read_643, op_fetch_5_read_644, op_fetch_5_read_645, op_fetch_5_read_646, op_fetch_5_read_647, op_fetch_5_read_648, op_fetch_5_read_649, op_fetch_5_read_650, op_fetch_5_read_651, op_fetch_5_read_652, op_fetch_5_read_653, op_fetch_5_read_654, op_fetch_5_read_655, op_fetch_5_read_656, op_fetch_5_read_657, op_fetch_5_read_658, op_fetch_5_read_659, op_fetch_5_read_660, op_fetch_5_read_661, op_fetch_5_read_662, op_fetch_5_read_663, op_fetch_5_read_664, op_fetch_5_read_665, op_fetch_5_read_666, op_fetch_5_read_667, op_fetch_5_read_668, op_fetch_5_read_669, op_fetch_5_read_670, op_fetch_5_read_671, op_fetch_5_read_672, op_fetch_5_read_673, op_fetch_5_read_674, op_fetch_5_read_675, op_fetch_5_read_676, op_fetch_5_read_677, op_fetch_5_read_678, op_fetch_5_read_679, op_fetch_5_read_680, op_fetch_5_read_681, op_fetch_5_read_682, op_fetch_5_read_683, op_fetch_5_read_684, op_fetch_5_read_685, op_fetch_5_read_686, op_fetch_5_read_687, op_fetch_5_read_688, op_fetch_5_read_689, op_fetch_5_read_690, op_fetch_5_read_691, op_fetch_5_read_692, op_fetch_5_read_693, op_fetch_5_read_694, op_fetch_5_read_695, op_fetch_5_read_696, op_fetch_5_read_697, op_fetch_5_read_698, op_fetch_5_read_699, op_fetch_5_read_700, op_fetch_5_read_701, op_fetch_5_read_702, op_fetch_5_read_703, op_fetch_5_read_704, op_fetch_5_read_705, op_fetch_5_read_706, op_fetch_5_read_707, op_fetch_5_read_708, op_fetch_5_read_709, op_fetch_5_read_710, op_fetch_5_read_711, op_fetch_5_read_712, op_fetch_5_read_713, op_fetch_5_read_714, op_fetch_5_read_715, op_fetch_5_read_716, op_fetch_5_read_717, op_fetch_5_read_718, op_fetch_5_read_719, op_fetch_5_read_720, op_fetch_5_read_721, op_fetch_5_read_722, op_fetch_5_read_723, op_fetch_5_read_724, op_fetch_5_read_725, op_fetch_5_read_726, op_fetch_5_read_727, op_fetch_5_read_728, op_fetch_5_read_729, op_fetch_5_read_730, op_fetch_5_read_731, op_fetch_5_read_732, op_fetch_5_read_733, op_fetch_5_read_734, op_fetch_5_read_735, op_fetch_5_read_736, op_fetch_5_read_737, op_fetch_5_read_738, op_fetch_5_read_739, op_fetch_5_read_740, op_fetch_5_read_741, op_fetch_5_read_742, op_fetch_5_read_743, op_fetch_5_read_744, op_fetch_5_read_745, op_fetch_5_read_746, op_fetch_5_read_747, op_fetch_5_read_748, op_fetch_5_read_749, op_fetch_5_read_750, op_fetch_5_read_751, op_fetch_5_read_752, op_fetch_5_read_753, op_fetch_5_read_754, op_fetch_5_read_755, op_fetch_5_read_756, op_fetch_5_read_757, op_fetch_5_read_758, op_fetch_5_read_759, op_fetch_5_read_760, op_fetch_5_read_761, op_fetch_5_read_762, op_fetch_5_read_763, op_fetch_5_read_764, op_fetch_5_read_765, op_fetch_5_read_766, op_fetch_5_read_767, op_fetch_5_read_768, op_fetch_5_read_769, op_fetch_5_read_770, op_fetch_5_read_771, op_fetch_5_read_772, op_fetch_5_read_773, op_fetch_5_read_774, op_fetch_5_read_775, op_fetch_5_read_776, op_fetch_5_read_777, op_fetch_5_read_778, op_fetch_5_read_779, op_fetch_5_read_780, op_fetch_5_read_781, op_fetch_5_read_782, op_fetch_5_read_783, op_fetch_5_read_784, op_fetch_5_read_785, op_fetch_5_read_786, op_fetch_5_read_787, op_fetch_5_read_788, op_fetch_5_read_789, op_fetch_5_read_790, op_fetch_5_read_791, op_fetch_5_read_792, op_fetch_5_read_793, op_fetch_5_read_794, op_fetch_5_read_795, op_fetch_5_read_796, op_fetch_5_read_797, op_fetch_5_read_798, op_fetch_5_read_799, op_fetch_5_read_800, op_fetch_5_read_801, op_fetch_5_read_802, op_fetch_5_read_803, op_fetch_5_read_804, op_fetch_5_read_805, op_fetch_5_read_806, op_fetch_5_read_807, op_fetch_5_read_808, op_fetch_5_read_809, op_fetch_5_read_810, op_fetch_5_read_811, op_fetch_5_read_812, op_fetch_5_read_813, op_fetch_5_read_814, op_fetch_5_read_815, op_fetch_5_read_816, op_fetch_5_read_817, op_fetch_5_read_818, op_fetch_5_read_819, op_fetch_5_read_820, op_fetch_5_read_821, op_fetch_5_read_822, op_fetch_5_read_823, op_fetch_5_read_824, op_fetch_5_read_825, op_fetch_5_read_826, op_fetch_5_read_827, op_fetch_5_read_828, op_fetch_5_read_829, op_fetch_5_read_830, op_fetch_5_read_831, op_fetch_5_read_832, op_fetch_5_read_833, op_fetch_5_read_834, op_fetch_5_read_835, op_fetch_5_read_836, op_fetch_5_read_837, op_fetch_5_read_838, op_fetch_5_read_839, op_fetch_5_read_840, op_fetch_5_read_841, op_fetch_5_read_842, op_fetch_5_read_843, op_fetch_5_read_844, op_fetch_5_read_845, op_fetch_5_read_846, op_fetch_5_read_847, op_fetch_5_read_848, op_fetch_5_read_849, op_fetch_5_read_850, op_fetch_5_read_851, op_fetch_5_read_852, op_fetch_5_read_853, op_fetch_5_read_854, op_fetch_5_read_855, op_fetch_5_read_856, op_fetch_5_read_857, op_fetch_5_read_858, op_fetch_5_read_859, op_fetch_5_read_860, op_fetch_5_read_861, op_fetch_5_read_862, op_fetch_5_read_863, op_fetch_5_read_864, op_fetch_5_read_865, op_fetch_5_read_866, op_fetch_5_read_867, op_fetch_5_read_868, op_fetch_5_read_869, op_fetch_5_read_870, op_fetch_5_read_871, op_fetch_5_read_872, op_fetch_5_read_873, op_fetch_5_read_874, op_fetch_5_read_875, op_fetch_5_read_876, op_fetch_5_read_877, op_fetch_5_read_878, op_fetch_5_read_879, op_fetch_5_read_880, op_fetch_5_read_881, op_fetch_5_read_882, op_fetch_5_read_883, op_fetch_5_read_884, op_fetch_5_read_885, op_fetch_5_read_886, op_fetch_5_read_887, op_fetch_5_read_888, op_fetch_5_read_889, op_fetch_5_read_890, op_fetch_5_read_891, op_fetch_5_read_892, op_fetch_5_read_893, op_fetch_5_read_894, op_fetch_5_read_895, op_fetch_5_read_896, op_fetch_5_read_897, op_fetch_5_read_898, op_fetch_5_read_899, op_fetch_5_read_900, op_fetch_5_read_901, op_fetch_5_read_902, op_fetch_5_read_903, op_fetch_5_read_904, op_fetch_5_read_905, op_fetch_5_read_906, op_fetch_5_read_907, op_fetch_5_read_908, op_fetch_5_read_909, op_fetch_5_read_910, op_fetch_5_read_911, op_fetch_5_read_912, op_fetch_5_read_913, op_fetch_5_read_914, op_fetch_5_read_915, op_fetch_5_read_916, op_fetch_5_read_917, op_fetch_5_read_918, op_fetch_5_read_919, op_fetch_5_read_920, op_fetch_5_read_921, op_fetch_5_read_922, op_fetch_5_read_923, op_fetch_5_read_924, op_fetch_5_read_925, op_fetch_5_read_926, op_fetch_5_read_927, op_fetch_5_read_928, op_fetch_5_read_929, op_fetch_5_read_930, op_fetch_5_read_931, op_fetch_5_read_932, op_fetch_5_read_933, op_fetch_5_read_934, op_fetch_5_read_935, op_fetch_5_read_936, op_fetch_5_read_937, op_fetch_5_read_938, op_fetch_5_read_939, op_fetch_5_read_940, op_fetch_5_read_941, op_fetch_5_read_942, op_fetch_5_read_943, op_fetch_5_read_944, op_fetch_5_read_945, op_fetch_5_read_946, op_fetch_5_read_947, op_fetch_5_read_948, op_fetch_5_read_949, op_fetch_5_read_950, op_fetch_5_read_951, op_fetch_5_read_952, op_fetch_5_read_953, op_fetch_5_read_954, op_fetch_5_read_955, op_fetch_5_read_956, op_fetch_5_read_957, op_fetch_5_read_958, op_fetch_5_read_959, op_fetch_5_read_960, op_fetch_5_read_961, op_fetch_5_read_962, op_fetch_5_read_963, op_fetch_5_read_964, op_fetch_5_read_965, op_fetch_5_read_966, op_fetch_5_read_967, op_fetch_5_read_968, op_fetch_5_read_969, op_fetch_5_read_970, op_fetch_5_read_971, op_fetch_5_read_972, op_fetch_5_read_973, op_fetch_5_read_974, op_fetch_5_read_975, op_fetch_5_read_976, op_fetch_5_read_977, op_fetch_5_read_978, op_fetch_5_read_979, op_fetch_5_read_980, op_fetch_5_read_981, op_fetch_5_read_982, op_fetch_5_read_983, op_fetch_5_read_984, op_fetch_5_read_985, op_fetch_5_read_986, op_fetch_5_read_987, op_fetch_5_read_988, op_executeALU_2_read_0, op_readRegisterFile_8_write_1004, op_readRegisterFile_8_write_1005, op_readRegisterFile_8_write_1006, op_readRegisterFile_8_write_1007, op_readRegisterFile_8_write_1008, op_readRegisterFile_8_write_1009, op_readRegisterFile_8_write_1010, op_readRegisterFile_8_write_1011, op_readRegisterFile_8_write_1012, op_readRegisterFile_8_write_1013, op_readRegisterFile_8_write_1014, op_readRegisterFile_8_write_1015, op_readRegisterFile_8_write_1016, op_readRegisterFile_8_write_1017, op_readRegisterFile_8_write_1018, op_readRegisterFile_8_write_1019, op_readRegisterFile_8_write_1020, op_readRegisterFile_8_write_1021, op_readRegisterFile_8_write_1022, op_readRegisterFile_8_write_1023, op_readRegisterFile_8_write_1024, op_readRegisterFile_8_write_1025, op_readRegisterFile_8_write_1026, op_readRegisterFile_8_write_1027, op_readRegisterFile_8_write_1028, op_readRegisterFile_8_write_1029, op_readRegisterFile_8_write_1030, op_readRegisterFile_8_write_1031, op_readRegisterFile_8_write_1032, op_readRegisterFile_8_write_1033, op_readRegisterFile_8_write_1034, op_readRegisterFile_8_write_1035, op_readRegisterFile_8_write_1036, op_readRegisterFile_8_write_1037, op_readRegisterFile_8_write_1038, op_readRegisterFile_8_write_1039, op_readRegisterFile_8_write_1040, op_readRegisterFile_8_write_1041, op_readRegisterFile_8_write_1042, op_readRegisterFile_8_write_1043, op_readRegisterFile_8_write_1044, op_readRegisterFile_8_write_1045, op_readRegisterFile_8_write_1046, op_readRegisterFile_8_write_1047, op_readRegisterFile_8_write_1048, op_readRegisterFile_8_write_1049, op_readRegisterFile_8_write_1050, op_readRegisterFile_8_write_1051, op_readRegisterFile_8_write_1052, op_readRegisterFile_8_write_1053, op_readRegisterFile_8_write_1054, op_readRegisterFile_8_write_1055, op_readRegisterFile_8_write_1056, op_readRegisterFile_8_write_1057, op_readRegisterFile_8_write_1058, op_readRegisterFile_8_write_1059, op_readRegisterFile_8_write_1060, op_readRegisterFile_8_write_1061, op_readRegisterFile_8_write_1062, op_readRegisterFile_8_write_1063, op_readRegisterFile_8_write_1064, op_readRegisterFile_8_write_1065, op_readRegisterFile_8_write_1066, op_readRegisterFile_8_write_1067, op_readRegisterFile_8_write_1068, op_readRegisterFile_8_write_1069, op_readRegisterFile_8_write_1070, op_readRegisterFile_8_write_1071, op_readRegisterFile_8_write_1072, op_readRegisterFile_8_write_1073, op_readRegisterFile_8_write_1074, op_readRegisterFile_8_write_1075, op_readRegisterFile_8_write_1076, op_readRegisterFile_8_write_1077, op_readRegisterFile_8_write_1078, op_readRegisterFile_8_write_1079, op_readRegisterFile_8_write_1080, op_readRegisterFile_8_write_1081, op_readRegisterFile_8_write_1082, op_readRegisterFile_8_write_1083, op_readRegisterFile_8_write_1084, op_readRegisterFile_8_write_1085, op_readRegisterFile_8_write_1086, op_readRegisterFile_8_write_1087, op_readRegisterFile_8_write_1088, op_readRegisterFile_8_write_1089, op_readRegisterFile_8_write_1090, op_readRegisterFile_8_write_1091, op_readRegisterFile_8_write_1092, op_readRegisterFile_8_write_1093, op_readRegisterFile_8_write_1094, op_readRegisterFile_8_write_1095, op_readRegisterFile_8_write_1096, op_readRegisterFile_8_write_1097, op_readRegisterFile_8_write_1098, op_readRegisterFile_8_write_1099, op_readRegisterFile_8_write_1100, op_readRegisterFile_8_write_1101, op_readRegisterFile_8_write_1102, op_readRegisterFile_8_write_1103, op_readRegisterFile_8_write_1104, op_readRegisterFile_8_write_1105, op_readRegisterFile_8_write_1106, op_readRegisterFile_8_write_1107, op_readRegisterFile_8_write_1108, op_readRegisterFile_8_write_1109, op_readRegisterFile_8_write_1110, op_readRegisterFile_8_write_1111, op_readRegisterFile_8_write_1112, op_readRegisterFile_8_write_1113, op_readRegisterFile_8_write_1114, op_readRegisterFile_8_write_1115, op_readRegisterFile_8_write_1116, op_readRegisterFile_8_write_1117, op_readRegisterFile_8_write_1118, op_readRegisterFile_8_write_1119, op_readRegisterFile_8_write_1120, op_readRegisterFile_8_write_1121, op_readRegisterFile_8_write_1122, op_readRegisterFile_8_write_1123, op_readRegisterFile_8_write_1124, op_readRegisterFile_8_write_1125, op_readRegisterFile_8_write_1126, op_readRegisterFile_8_write_1127, op_readRegisterFile_8_write_1128, op_readRegisterFile_8_write_1129, op_readRegisterFile_8_write_1130, op_readRegisterFile_8_write_1131, op_readRegisterFile_8_write_1132, op_readRegisterFile_8_write_1133, op_readRegisterFile_8_write_1134, op_readRegisterFile_8_write_1135, op_readRegisterFile_8_write_1136, op_readRegisterFile_8_write_1137, op_readRegisterFile_8_write_1138, op_readRegisterFile_8_write_1139, op_readRegisterFile_8_write_1140, op_readRegisterFile_8_write_1141, op_readRegisterFile_8_write_1142, op_readRegisterFile_8_write_1143, op_readRegisterFile_8_write_1144, op_readRegisterFile_8_write_1145, op_readRegisterFile_8_write_1146, op_readRegisterFile_8_write_1147, op_readRegisterFile_8_write_1148, op_readRegisterFile_8_write_1149, op_readRegisterFile_8_write_1150, op_readRegisterFile_8_write_1151, op_readRegisterFile_8_write_1152, op_readRegisterFile_8_write_1153, op_readRegisterFile_8_write_1154, op_readRegisterFile_8_write_1155, op_readRegisterFile_8_write_1156, op_readRegisterFile_8_write_1157, op_readRegisterFile_8_write_1158, op_readRegisterFile_8_write_1159, op_readRegisterFile_8_write_1160, op_readRegisterFile_8_write_1161, op_readRegisterFile_8_write_1162, op_readRegisterFile_8_write_1163, op_readRegisterFile_8_write_1164, op_readRegisterFile_8_write_1165, op_readRegisterFile_8_write_1166, op_readRegisterFile_8_write_1167, op_readRegisterFile_8_write_1168, op_readRegisterFile_8_write_1169, op_readRegisterFile_8_write_1170, op_readRegisterFile_8_write_1171, op_readRegisterFile_8_write_1172, op_readRegisterFile_8_write_1173, op_readRegisterFile_8_write_1174, op_readRegisterFile_8_write_1175, op_readRegisterFile_8_write_1176, op_readRegisterFile_8_write_1177, op_readRegisterFile_8_write_1178, op_readRegisterFile_8_write_1179, op_readRegisterFile_8_write_1180, op_readRegisterFile_8_write_1181, op_readRegisterFile_8_write_1182, op_readRegisterFile_8_write_1183, op_readRegisterFile_8_write_1184, op_readRegisterFile_8_write_1185, op_readRegisterFile_8_write_1186, op_readRegisterFile_8_write_1187, op_readRegisterFile_8_write_1188, op_readRegisterFile_8_write_1189, op_readRegisterFile_8_write_1190, op_readRegisterFile_8_write_1191, op_readRegisterFile_8_write_1192, op_readRegisterFile_8_write_1193, op_readRegisterFile_8_write_1194, op_readRegisterFile_8_write_1195, op_readRegisterFile_8_write_1196, op_readRegisterFile_8_write_1197, op_readRegisterFile_8_write_1198, op_readRegisterFile_8_write_1199, op_readRegisterFile_8_write_1200, op_readRegisterFile_8_write_1201, op_readRegisterFile_8_write_1202, op_readRegisterFile_8_write_1203, op_readRegisterFile_8_write_1204, op_readRegisterFile_8_write_1205, op_readRegisterFile_8_write_1206, op_readRegisterFile_8_write_1207, op_readRegisterFile_8_write_1208, op_readRegisterFile_8_write_1209, op_readRegisterFile_8_write_1210, op_readRegisterFile_8_write_1211, op_readRegisterFile_8_write_1212, op_readRegisterFile_8_write_1213, op_readRegisterFile_8_write_1214, op_readRegisterFile_8_write_1215, op_executeALU_3_read_1, op_executeALU_3_read_2, op_executeALU_3_read_3, op_executeALU_3_read_4, op_executeALU_3_read_5, op_executeALU_3_read_6, op_executeALU_3_read_7, op_executeALU_3_read_8, op_executeALU_3_read_9, op_executeALU_3_read_10, op_executeALU_3_read_11, op_executeALU_3_read_12, op_executeALU_3_read_13, op_executeALU_3_read_14, op_executeALU_3_read_15, op_executeALU_3_read_16, op_executeALU_3_read_17, op_executeALU_3_read_18, op_executeALU_3_read_19, op_executeALU_3_read_20, op_executeALU_3_read_21, op_executeALU_3_read_22, op_executeALU_3_read_23, op_executeALU_3_read_24, op_executeALU_3_read_25, op_executeALU_3_read_26, op_executeALU_3_read_27, op_executeALU_3_read_28, op_executeALU_3_read_29, op_executeALU_3_read_30, op_executeALU_3_read_31, op_executeALU_3_read_32, op_executeALU_3_read_33, op_executeALU_3_read_34, op_executeALU_3_read_35, op_executeALU_3_read_36, op_executeALU_3_read_37, op_executeALU_3_read_38, op_executeALU_3_read_39, op_executeALU_3_read_40, op_executeALU_3_read_41, op_executeALU_3_read_42, op_executeALU_3_read_43, op_executeALU_3_read_44, op_executeALU_3_read_45, op_executeALU_3_read_46, op_executeALU_3_read_47, op_executeALU_3_read_48, op_executeALU_3_read_49, op_executeALU_3_read_50, op_executeALU_3_read_51, op_executeALU_3_read_52, op_executeALU_3_read_53, op_executeALU_3_read_54, op_executeALU_3_read_55, op_executeALU_3_read_56, op_executeALU_3_read_57, op_executeALU_3_read_58, op_executeALU_3_read_59, op_executeALU_3_read_60, op_executeALU_3_read_61, op_executeALU_3_read_62, op_executeALU_3_read_63, op_executeALU_3_read_64, op_executeALU_3_read_65, op_executeALU_3_read_66, op_executeALU_3_read_67, op_executeALU_3_read_68, op_executeALU_3_read_69, op_executeALU_3_read_70, op_executeALU_3_read_71, op_executeALU_3_read_72, op_executeALU_3_read_73, op_executeALU_3_read_74, op_executeALU_3_read_75, op_executeALU_3_read_76, op_executeALU_3_read_77, op_executeALU_3_read_78, op_executeALU_3_read_79, op_executeALU_3_read_80, op_executeALU_3_read_81, op_executeALU_3_read_82, op_executeALU_3_read_83, op_executeALU_3_read_84, op_executeALU_3_read_85, op_executeALU_3_read_86, op_executeALU_3_read_87, op_executeALU_3_read_88, op_executeALU_3_read_89, op_executeALU_3_read_90, op_executeALU_3_read_91, op_executeALU_3_read_92, op_executeALU_3_read_93, op_executeALU_3_read_94, op_executeALU_3_read_95, op_executeALU_3_read_96, op_memoryOperation_6_write_989, op_memoryOperation_6_write_990, op_memoryOperation_6_write_991, op_memoryOperation_6_write_992, op_wait_memoryOperation_6, op_memoryOperation_6_write_993, op_memoryOperation_6_write_994, op_memoryOperation_6_write_995, op_memoryOperation_6_write_996, op_writeBack_10_write_1216, op_memoryOperation_7_read_997, op_memoryOperation_7_read_998, op_memoryOperation_7_read_999, op_memoryOperation_7_read_1000, op_wait_memoryOperation_7, op_memoryOperation_7_read_1001, op_memoryOperation_7_read_1002, op_memoryOperation_7_read_1003);
	type ISA_state_t is (st_executeALU_2, st_executeALU_3, st_fetch_4, st_fetch_5, st_memoryOperation_6, st_memoryOperation_7, st_readRegisterFile_8, st_writeBack_10);
	type ALUtoCtl_IF is record
		ALU_result: unsigned(31 downto 0);
	end record;
	type ALU_function is (ALU_ADD, ALU_AND, ALU_COPY1, ALU_OR, ALU_SLL, ALU_SLT, ALU_SLTU, ALU_SRA, ALU_SRL, ALU_SUB, ALU_X, ALU_XOR);
	type ALUopType is (OP_IMM, OP_PC, OP_REG, OP_X);
	type CtlToALU_IF is record
		alu_fun: ALU_function;
		imm: unsigned(31 downto 0);
		op1_sel: ALUopType;
		op2_sel: ALUopType;
		pc_reg: unsigned(31 downto 0);
		reg1_contents: unsigned(31 downto 0);
		reg2_contents: unsigned(31 downto 0);
	end record;
	type WBselType is (WB_ALU, WB_MEM, WB_PC4, WB_X);

	-- Declare signals
	signal active_state: ISA_state_t;
	signal active_operation: ISA_operation_t;
	signal ALUtoCtl_data: ALUtoCtl_IF;
	signal CtlToALU_data: CtlToALU_IF;
	signal CtlToRegs_data: CtlToRegs_IF;
	signal RegsToCtl_data: RegsToCtl_IF;
	signal br_en: boolean;
	signal decodedInstr: DecodedInstr;
	signal fromMemoryData: MEtoCU_IF;
	signal mem_en: boolean;
	signal memoryAccess: CUtoME_IF;
	signal pc_next: unsigned(31 downto 0);
	signal pc_reg: unsigned(31 downto 0);
	signal reg_rd_en: boolean;
	signal wb_en: boolean;
	signal wb_sel: WBselType;

	-- Declare state signals that are used by ITL properties for OneSpin
	signal executeALU_2: boolean;
	signal executeALU_3: boolean;
	signal fetch_4: boolean;
	signal fetch_5: boolean;
	signal memoryOperation_6: boolean;
	signal memoryOperation_7: boolean;
	signal readRegisterFile_8: boolean;
	signal writeBack_10: boolean;


begin
	-- Combinational logic that selects current operation
	process (active_state, CtlToMem_port_sync, MemToCtl_port_sync, DecToCtl_port_sig.instrType, DecToCtl_port_sig.imm, RegsToCtl_port_sig.contents2, RegsToCtl_port_sig.contents1, DecToCtl_port_sig.encType, memoryAccess.req, pc_reg, ALUtoCtl_data.ALU_result, mem_en, CtlToALU_data.alu_fun, wb_sel, CtlToALU_data.op1_sel, CtlToALU_data.op2_sel, decodedInstr.instrType, decodedInstr.rd_addr, decodedInstr.imm, br_en, RegsToCtl_data.contents2, reg_rd_en, wb_en, RegsToCtl_data.contents1)
	begin
	active_operation <= op_wait_fetch_4;
		case active_state is
		when st_executeALU_2 =>
			if (true) then 
				active_operation <= op_executeALU_2_read_0;
			end if;
		when st_executeALU_3 =>
			if (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_1;
			elsif (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_2;
			elsif (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4)) then 
				active_operation <= op_executeALU_3_read_3;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_4;
			elsif (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_5;
			elsif (br_en and (decodedInstr.instrType = beq) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_6;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_7;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4)) then 
				active_operation <= op_executeALU_3_read_8;
			elsif (br_en and (decodedInstr.instrType = beq) and not(mem_en) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_9;
			elsif (br_en and (decodedInstr.instrType = beq) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_10;
			elsif (br_en and (decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000") and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_11;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_12;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_13;
			elsif (br_en and (decodedInstr.instrType = beq) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_14;
			elsif (br_en and (decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000") and not(mem_en) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_15;
			elsif (br_en and (decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000") and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4)) then 
				active_operation <= op_executeALU_3_read_16;
			elsif (br_en and (decodedInstr.instrType = blt) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_17;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_18;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4)) then 
				active_operation <= op_executeALU_3_read_19;
			elsif (br_en and (decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000") and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_20;
			elsif (br_en and (decodedInstr.instrType = blt) and not(mem_en) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_21;
			elsif (br_en and (decodedInstr.instrType = blt) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_22;
			elsif (br_en and (decodedInstr.instrType = bge) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_23;
			elsif (br_en and not((decodedInstr.instrType = beq) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = blt) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bge) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bltu) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bgeu) and (ALUtoCtl_data.ALU_result = x"00000000")) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_24;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_25;
			elsif (br_en and (decodedInstr.instrType = blt) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_26;
			elsif (br_en and (decodedInstr.instrType = bge) and not(mem_en) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_27;
			elsif (br_en and (decodedInstr.instrType = bge) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_28;
			elsif (br_en and (decodedInstr.instrType = bltu) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_29;
			elsif (br_en and not((decodedInstr.instrType = beq) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = blt) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bge) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bltu) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bgeu) and (ALUtoCtl_data.ALU_result = x"00000000")) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_30;
			elsif (br_en and not((decodedInstr.instrType = beq) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = blt) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bge) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bltu) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bgeu) and (ALUtoCtl_data.ALU_result = x"00000000")) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4)) then 
				active_operation <= op_executeALU_3_read_31;
			elsif (br_en and (decodedInstr.instrType = bge) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_32;
			elsif (br_en and (decodedInstr.instrType = bltu) and not(mem_en) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_33;
			elsif (br_en and (decodedInstr.instrType = bltu) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_34;
			elsif (br_en and (decodedInstr.instrType = bgeu) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_35;
			elsif (br_en and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_36;
			elsif (br_en and not((decodedInstr.instrType = beq) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = blt) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bge) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bltu) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bgeu) and (ALUtoCtl_data.ALU_result = x"00000000")) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_37;
			elsif (br_en and (decodedInstr.instrType = bltu) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_38;
			elsif (br_en and (decodedInstr.instrType = bgeu) and not(mem_en) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_39;
			elsif (br_en and (decodedInstr.instrType = bgeu) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_40;
			elsif (br_en and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_41;
			elsif (br_en and (decodedInstr.instrType = jal) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4)) then 
				active_operation <= op_executeALU_3_read_42;
			elsif (br_en and (decodedInstr.instrType = bgeu) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_43;
			elsif (br_en and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_44;
			elsif (br_en and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_45;
			elsif (br_en and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_46;
			elsif (br_en and (decodedInstr.instrType = jalr) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4)) then 
				active_operation <= op_executeALU_3_read_47;
			elsif (br_en and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_48;
			elsif (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and mem_en) then 
				active_operation <= op_executeALU_3_read_49;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and mem_en) then 
				active_operation <= op_executeALU_3_read_50;
			elsif (br_en and (decodedInstr.instrType = beq) and mem_en and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_51;
			elsif (br_en and (decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000") and mem_en) then 
				active_operation <= op_executeALU_3_read_52;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and mem_en) then 
				active_operation <= op_executeALU_3_read_53;
			elsif (br_en and (decodedInstr.instrType = blt) and mem_en and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_54;
			elsif (br_en and (decodedInstr.instrType = bge) and mem_en and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_55;
			elsif (br_en and not((decodedInstr.instrType = beq) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = blt) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bge) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bltu) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bgeu) and (ALUtoCtl_data.ALU_result = x"00000000")) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and mem_en) then 
				active_operation <= op_executeALU_3_read_56;
			elsif (br_en and (decodedInstr.instrType = bltu) and mem_en and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_57;
			elsif (br_en and (decodedInstr.instrType = bgeu) and mem_en and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_58;
			elsif (br_en and (decodedInstr.instrType = jal) and mem_en) then 
				active_operation <= op_executeALU_3_read_59;
			elsif (br_en and (decodedInstr.instrType = jalr) and mem_en) then 
				active_operation <= op_executeALU_3_read_60;
			elsif (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_61;
			elsif (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_62;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_63;
			elsif (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_64;
			elsif (br_en and (decodedInstr.instrType = beq) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_65;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_66;
			elsif (br_en and (decodedInstr.instrType = beq) and not(mem_en) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_67;
			elsif (br_en and (decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000") and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_68;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_69;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_70;
			elsif (br_en and (decodedInstr.instrType = beq) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_71;
			elsif (br_en and (decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000") and not(mem_en) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_72;
			elsif (br_en and (decodedInstr.instrType = blt) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_73;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_74;
			elsif (br_en and (decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000") and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_75;
			elsif (br_en and (decodedInstr.instrType = blt) and not(mem_en) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_76;
			elsif (br_en and (decodedInstr.instrType = bge) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_77;
			elsif (br_en and not((decodedInstr.instrType = beq) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = blt) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bge) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bltu) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bgeu) and (ALUtoCtl_data.ALU_result = x"00000000")) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_78;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_79;
			elsif (br_en and (decodedInstr.instrType = blt) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_80;
			elsif (br_en and (decodedInstr.instrType = bge) and not(mem_en) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_81;
			elsif (br_en and (decodedInstr.instrType = bltu) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_82;
			elsif (br_en and not((decodedInstr.instrType = beq) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = blt) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bge) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bltu) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bgeu) and (ALUtoCtl_data.ALU_result = x"00000000")) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_83;
			elsif (br_en and (decodedInstr.instrType = bge) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_84;
			elsif (br_en and (decodedInstr.instrType = bltu) and not(mem_en) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_85;
			elsif (br_en and (decodedInstr.instrType = bgeu) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_86;
			elsif (br_en and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_87;
			elsif (br_en and not((decodedInstr.instrType = beq) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = blt) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bge) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bltu) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bgeu) and (ALUtoCtl_data.ALU_result = x"00000000")) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_88;
			elsif (br_en and (decodedInstr.instrType = bltu) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_89;
			elsif (br_en and (decodedInstr.instrType = bgeu) and not(mem_en) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_90;
			elsif (br_en and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_91;
			elsif (br_en and (decodedInstr.instrType = bgeu) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000") and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_92;
			elsif (br_en and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_93;
			elsif (br_en and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_94;
			elsif (br_en and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_95;
			elsif (br_en and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_96;
			end if;
		when st_fetch_4 =>
			if (not(CtlToMem_port_sync)) then 
				active_operation <= op_wait_fetch_4;
			elsif (CtlToMem_port_sync) then 
				active_operation <= op_fetch_4_write_97;
			end if;
		when st_fetch_5 =>
			if (not(MemToCtl_port_sync)) then 
				active_operation <= op_wait_fetch_5;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_98;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_99;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_100;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_101;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_102;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_103;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_104;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_105;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_106;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_107;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_108;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_109;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_110;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_111;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_112;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_113;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_114;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_115;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_116;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_117;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_118;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_119;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_120;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_121;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_122;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_123;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_124;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_125;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_126;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_127;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_128;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_129;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_130;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_131;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_132;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_133;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_134;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_135;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_136;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_137;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_138;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_139;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_140;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_141;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_142;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_143;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_144;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_145;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_146;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_147;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_148;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_149;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_150;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_151;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_152;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_153;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_154;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_155;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_156;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_157;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_158;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_159;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_160;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_161;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_162;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_163;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_164;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_165;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_166;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_167;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_168;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_169;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_170;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_171;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_172;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_173;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_174;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_175;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_176;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_177;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_178;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_179;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_180;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_181;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_182;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_183;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_184;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_185;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_186;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_187;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_188;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_189;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_190;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_191;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_192;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_193;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_194;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_195;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_196;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_197;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_198;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_199;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_200;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_201;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_202;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_203;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_204;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_205;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_206;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_207;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_208;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_209;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_210;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_211;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_212;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_213;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_214;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_215;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_216;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_217;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_218;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_219;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_220;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_221;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_222;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_223;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_224;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_225;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_226;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_227;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_228;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_229;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_230;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_231;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_232;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_233;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_234;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_235;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_236;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_237;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_238;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_239;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_240;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_241;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_242;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_243;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_244;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_245;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_246;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_247;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_248;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_249;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_250;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_251;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_252;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_253;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_254;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_255;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_256;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_257;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_258;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_259;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_260;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_261;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_262;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_263;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_264;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_265;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_266;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_267;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_268;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_269;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_270;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_271;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_272;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_273;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_274;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_275;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_276;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_277;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_278;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_279;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_280;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_281;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_282;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_283;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_284;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_285;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_286;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_287;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_288;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_289;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_290;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_291;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_292;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_293;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_294;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_295;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_296;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_297;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_298;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_299;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_300;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_301;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_302;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_303;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_304;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_305;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_306;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_307;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_308;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_309;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_310;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_311;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_312;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_313;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_314;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_315;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_316;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_317;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_318;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_319;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_320;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_321;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_322;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_323;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_324;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_325;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_326;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_327;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_328;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_329;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_330;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_331;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_332;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_333;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_334;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_335;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_336;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_337;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_338;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_339;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_340;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_341;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_342;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_343;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_344;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_345;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_346;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_347;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_348;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_349;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_350;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_351;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_352;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_353;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_354;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_355;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_356;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_357;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_358;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_359;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_360;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_361;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_362;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_363;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_364;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_365;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_366;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_367;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_368;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_369;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_370;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_371;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_372;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_373;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_374;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_375;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_376;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_377;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_378;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_379;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_380;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_381;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_382;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_383;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_384;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_385;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_386;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_387;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_388;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_389;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_390;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_391;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_392;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_393;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_394;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_395;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_396;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_397;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_398;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_399;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_400;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_401;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_402;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_403;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_404;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_405;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_406;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_407;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_408;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_409;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_410;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_411;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_412;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_413;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_414;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_415;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_416;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_417;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_418;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_419;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_420;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_421;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_422;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_423;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_424;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_425;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_426;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_427;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_428;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_429;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_430;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_431;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_432;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_433;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_434;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_435;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_436;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_437;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_438;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_439;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_440;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_441;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_442;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_443;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_444;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_445;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_446;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_447;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_448;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_449;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_450;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_451;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_452;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_453;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_454;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_455;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_456;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_457;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_458;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_459;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_460;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_461;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_462;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_463;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_464;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_465;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_466;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_467;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_468;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_469;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_470;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_471;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_472;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_473;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_474;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_475;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_476;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_477;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_478;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_479;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_480;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_481;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_482;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_483;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_484;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_485;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_486;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_487;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_488;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_489;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_490;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_491;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_492;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_493;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_494;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_495;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_496;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_497;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_498;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_499;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_500;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_501;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_502;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_503;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_504;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_505;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_506;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_507;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_508;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_509;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_510;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_511;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_512;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_513;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_514;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_515;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_516;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_517;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_518;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_519;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_520;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_521;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_522;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_523;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_524;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_525;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_526;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_527;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_528;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_529;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_530;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_531;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_532;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_533;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_534;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_535;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_536;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_537;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_538;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_539;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_540;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_541;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_542;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_543;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_544;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_545;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_546;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_547;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_548;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_549;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_550;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_551;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_552;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_553;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_554;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_555;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_556;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_557;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_558;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_559;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_560;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_561;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_562;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_563;
			elsif ((DecToCtl_port_sig.encType = J) and (DecToCtl_port_sig.instrType = jal) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_564;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_565;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_566;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_567;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_568;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_569;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_570;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_571;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_572;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_573;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_574;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_575;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_576;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_577;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_578;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_579;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_580;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_581;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_582;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_583;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_584;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_585;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_586;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_587;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_588;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_589;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_590;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_591;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_592;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_593;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_594;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_595;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_596;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_597;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_598;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_599;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_600;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_601;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_602;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_603;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_604;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_605;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_606;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_607;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_608;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_609;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_610;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_611;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_612;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_613;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_614;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_615;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_616;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_617;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_618;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_619;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_620;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_621;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_622;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_623;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_624;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_625;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_626;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_627;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_628;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_629;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_630;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_631;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_632;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_633;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_634;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_635;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_636;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_637;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_638;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_639;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_640;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_641;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_642;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_643;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_644;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_645;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_646;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_647;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_648;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_649;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_650;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_651;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_652;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_653;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_654;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_655;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_656;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_657;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_658;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_659;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_660;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_661;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_662;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_663;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_664;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_665;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_666;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_667;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_668;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_669;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_670;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_671;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_672;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_673;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_674;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_675;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_676;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_677;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_678;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_679;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_680;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_681;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_682;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_683;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_684;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_685;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_686;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_687;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_688;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_689;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_690;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_691;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_692;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_693;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_694;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_695;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_696;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_697;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_698;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_699;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_700;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_701;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_702;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_703;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_704;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_705;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_706;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_707;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_708;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_709;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_710;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_711;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_712;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_713;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_714;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_715;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_716;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_717;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_718;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_719;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_720;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_721;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_722;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_723;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_724;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_725;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_726;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_727;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_728;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_729;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_730;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_731;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_732;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_733;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_734;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_735;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_736;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_737;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_738;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_739;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_740;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_741;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_742;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_743;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_744;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_745;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_746;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_747;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_748;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_749;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_750;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_751;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_752;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_753;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_754;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_755;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_756;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_757;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_758;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_759;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_760;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_761;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_762;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_763;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_764;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_765;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_766;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_767;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_768;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_769;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_770;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_771;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_772;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_773;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_774;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_775;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_776;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_777;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_778;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_779;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_780;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_781;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_782;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_783;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_784;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_785;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_786;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_787;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_788;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_789;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_790;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_791;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_792;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_793;
			elsif ((DecToCtl_port_sig.encType = U) and (DecToCtl_port_sig.instrType = auipc) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_794;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_795;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_796;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_797;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_798;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_799;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_800;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_801;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_802;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_803;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_804;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_805;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_806;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_807;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_808;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_809;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_810;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_811;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_812;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_813;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_814;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_815;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_816;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_817;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_818;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_819;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_820;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_821;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_822;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_823;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_824;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_825;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_826;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_827;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_828;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_829;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_830;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_831;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_832;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_833;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_834;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_835;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_836;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_837;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_838;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_839;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_840;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_841;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_842;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_843;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_844;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_845;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_846;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_847;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_848;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_849;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_850;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_851;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_852;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_853;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_854;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_855;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_856;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_857;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_858;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_859;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_860;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_861;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_862;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_863;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_864;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_865;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_866;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_867;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_868;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_869;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_870;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_871;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_872;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_873;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_874;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_875;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_876;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_877;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_878;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_879;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_880;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_881;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_882;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_883;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_884;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_885;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg <= DecToCtl_port_sig.imm) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_886;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_887;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_888;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_889;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_890;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_891;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm <= pc_reg) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_892;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_893;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_894;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_895;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_896;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_897;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_898;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_899;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_900;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_901;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_902;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_903;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_904;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_905;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_906;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_907;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_908;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_909;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_910;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_911;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_912;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_913;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_914;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_915;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_916;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_917;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_918;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_919;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_920;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_921;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_922;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_923;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_924;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_925;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_926;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_927;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_928;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_929;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_930;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_931;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_932;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_933;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_934;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_935;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_936;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_937;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_938;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_939;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_940;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_941;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_942;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_943;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_944;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_945;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_946;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_947;
			elsif ((DecToCtl_port_sig.encType = U) and (DecToCtl_port_sig.instrType = lui) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_948;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and reg_rd_en and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_949;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and reg_rd_en and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_950;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and reg_rd_en and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_951;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = addI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_952;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = add) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_953;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = sltI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_954;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = jalr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_955;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = sub) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_956;
			elsif ((DecToCtl_port_sig.encType = B) and (DecToCtl_port_sig.instrType = beq) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_957;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = sltIu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_958;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = sll_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_959;
			elsif ((DecToCtl_port_sig.encType = B) and (DecToCtl_port_sig.instrType = bne) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_960;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = xorI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_961;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = lb) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_962;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = slt) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_963;
			elsif ((DecToCtl_port_sig.encType = B) and (DecToCtl_port_sig.instrType = blt) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_964;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = orI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_965;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = lh) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_966;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = sltu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_967;
			elsif ((DecToCtl_port_sig.encType = B) and (DecToCtl_port_sig.instrType = bge) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_968;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = andI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_969;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = lw) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_970;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = Xor_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_971;
			elsif ((DecToCtl_port_sig.encType = B) and (DecToCtl_port_sig.instrType = bltu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_972;
			elsif ((DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.instrType = beq) and not(DecToCtl_port_sig.instrType = bne) and not(DecToCtl_port_sig.instrType = blt) and not(DecToCtl_port_sig.instrType = bge) and not(DecToCtl_port_sig.instrType = bltu) and not(DecToCtl_port_sig.instrType = bgeu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_973;
			elsif ((DecToCtl_port_sig.encType = S) and (DecToCtl_port_sig.instrType = sb) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_974;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = sllI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_975;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = lbu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_976;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = srl_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_977;
			elsif ((DecToCtl_port_sig.encType = B) and (DecToCtl_port_sig.instrType = bgeu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_978;
			elsif ((DecToCtl_port_sig.encType = S) and (DecToCtl_port_sig.instrType = sh) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_979;
			elsif ((DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.instrType = sb) and not(DecToCtl_port_sig.instrType = sh) and not(DecToCtl_port_sig.instrType = sw) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_980;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = srlI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_981;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = lhu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_982;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = sra_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_983;
			elsif ((DecToCtl_port_sig.encType = S) and (DecToCtl_port_sig.instrType = sw) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_984;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = sraI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_985;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = Or_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_986;
			elsif ((DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.instrType = add) and not(DecToCtl_port_sig.instrType = sub) and not(DecToCtl_port_sig.instrType = sll_Instr) and not(DecToCtl_port_sig.instrType = slt) and not(DecToCtl_port_sig.instrType = sltu) and not(DecToCtl_port_sig.instrType = Xor_Instr) and not(DecToCtl_port_sig.instrType = srl_Instr) and not(DecToCtl_port_sig.instrType = sra_Instr) and not(DecToCtl_port_sig.instrType = Or_Instr) and not(DecToCtl_port_sig.instrType = And_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_987;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = And_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_988;
			end if;
		when st_memoryOperation_6 =>
			if (not(memoryAccess.req = ME_RD) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and CtlToMem_port_sync) then 
				active_operation <= op_memoryOperation_6_write_989;
			elsif (not(memoryAccess.req = ME_RD) and (wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and CtlToMem_port_sync) then 
				active_operation <= op_memoryOperation_6_write_990;
			elsif (not(memoryAccess.req = ME_RD) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and CtlToMem_port_sync) then 
				active_operation <= op_memoryOperation_6_write_991;
			elsif (not(memoryAccess.req = ME_RD) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and CtlToMem_port_sync) then 
				active_operation <= op_memoryOperation_6_write_992;
			elsif (not(CtlToMem_port_sync)) then 
				active_operation <= op_wait_memoryOperation_6;
			elsif ((memoryAccess.req = ME_RD) and CtlToMem_port_sync) then 
				active_operation <= op_memoryOperation_6_write_993;
			elsif (not(memoryAccess.req = ME_RD) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000") and CtlToMem_port_sync) then 
				active_operation <= op_memoryOperation_6_write_994;
			elsif (not(memoryAccess.req = ME_RD) and (wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000") and CtlToMem_port_sync) then 
				active_operation <= op_memoryOperation_6_write_995;
			elsif (not(memoryAccess.req = ME_RD) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000") and CtlToMem_port_sync) then 
				active_operation <= op_memoryOperation_6_write_996;
			end if;
		when st_memoryOperation_7 =>
			if ((wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and MemToCtl_port_sync) then 
				active_operation <= op_memoryOperation_7_read_997;
			elsif ((wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and MemToCtl_port_sync) then 
				active_operation <= op_memoryOperation_7_read_998;
			elsif (not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and MemToCtl_port_sync) then 
				active_operation <= op_memoryOperation_7_read_999;
			elsif ((wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and MemToCtl_port_sync) then 
				active_operation <= op_memoryOperation_7_read_1000;
			elsif (not(MemToCtl_port_sync)) then 
				active_operation <= op_wait_memoryOperation_7;
			elsif ((wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_memoryOperation_7_read_1001;
			elsif ((wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_memoryOperation_7_read_1002;
			elsif ((wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_memoryOperation_7_read_1003;
			end if;
		when st_readRegisterFile_8 =>
			if ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1004;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1005;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1006;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1007;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1008;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1009;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1010;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1011;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1012;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1013;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1014;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1015;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1016;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1017;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1018;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1019;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1020;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1021;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1022;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1023;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1024;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1025;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1026;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1027;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1028;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1029;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1030;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1031;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1032;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1033;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1034;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1035;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1036;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1037;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1038;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1039;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1040;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1041;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1042;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1043;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1044;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1045;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1046;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1047;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1048;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1049;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1050;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1051;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1052;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1053;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1054;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1055;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1056;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1057;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1058;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1059;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1060;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1061;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1062;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1063;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1064;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1065;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1066;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1067;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1068;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1069;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1070;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1071;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1072;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1073;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1074;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_port_sig.contents2 <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1075;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_port_sig.contents2 <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1076;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1077;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1078;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1079;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1080;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1081;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1082;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1083;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1084;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1085;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1086;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1087;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1088;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1089;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_port_sig.contents2 <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1090;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_port_sig.contents2 <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1091;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1092;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(decodedInstr.imm <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1093;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (decodedInstr.imm <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1094;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_port_sig.contents2 <= decodedInstr.imm)) then 
				active_operation <= op_readRegisterFile_8_write_1095;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_port_sig.contents2 <= decodedInstr.imm)) then 
				active_operation <= op_readRegisterFile_8_write_1096;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1097;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1098;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1099;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1100;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1101;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1102;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1103;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1104;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1105;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(decodedInstr.imm <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1106;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (decodedInstr.imm <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1107;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1108;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1109;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1110;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT)) then 
				active_operation <= op_readRegisterFile_8_write_1111;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_port_sig.contents2 <= decodedInstr.imm)) then 
				active_operation <= op_readRegisterFile_8_write_1112;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_port_sig.contents2 <= decodedInstr.imm)) then 
				active_operation <= op_readRegisterFile_8_write_1113;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1114;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT)) then 
				active_operation <= op_readRegisterFile_8_write_1115;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_port_sig.contents2 <= pc_reg)) then 
				active_operation <= op_readRegisterFile_8_write_1116;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_port_sig.contents2 <= pc_reg)) then 
				active_operation <= op_readRegisterFile_8_write_1117;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1118;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1119;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_port_sig.contents2 = x"00000000")) then 
				active_operation <= op_readRegisterFile_8_write_1120;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_port_sig.contents2 = x"00000000")) then 
				active_operation <= op_readRegisterFile_8_write_1121;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1122;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1123;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1124;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1125;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1126;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1127;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1128;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU)) then 
				active_operation <= op_readRegisterFile_8_write_1129;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1130;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1131;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU)) then 
				active_operation <= op_readRegisterFile_8_write_1132;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1133;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg <= decodedInstr.imm)) then 
				active_operation <= op_readRegisterFile_8_write_1134;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg <= decodedInstr.imm)) then 
				active_operation <= op_readRegisterFile_8_write_1135;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT)) then 
				active_operation <= op_readRegisterFile_8_write_1136;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_port_sig.contents2 <= pc_reg)) then 
				active_operation <= op_readRegisterFile_8_write_1137;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_port_sig.contents2 <= pc_reg)) then 
				active_operation <= op_readRegisterFile_8_write_1138;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1139;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(decodedInstr.imm <= pc_reg)) then 
				active_operation <= op_readRegisterFile_8_write_1140;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (decodedInstr.imm <= pc_reg)) then 
				active_operation <= op_readRegisterFile_8_write_1141;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_port_sig.contents2 = x"00000000")) then 
				active_operation <= op_readRegisterFile_8_write_1142;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_port_sig.contents2 = x"00000000")) then 
				active_operation <= op_readRegisterFile_8_write_1143;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1144;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(decodedInstr.imm = x"00000000")) then 
				active_operation <= op_readRegisterFile_8_write_1145;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (decodedInstr.imm = x"00000000")) then 
				active_operation <= op_readRegisterFile_8_write_1146;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1147;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1148;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1149;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1150;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1151;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1152;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg <= decodedInstr.imm)) then 
				active_operation <= op_readRegisterFile_8_write_1153;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg <= decodedInstr.imm)) then 
				active_operation <= op_readRegisterFile_8_write_1154;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1155;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU)) then 
				active_operation <= op_readRegisterFile_8_write_1156;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1157;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1158;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(decodedInstr.imm <= pc_reg)) then 
				active_operation <= op_readRegisterFile_8_write_1159;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (decodedInstr.imm <= pc_reg)) then 
				active_operation <= op_readRegisterFile_8_write_1160;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1161;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT)) then 
				active_operation <= op_readRegisterFile_8_write_1162;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT)) then 
				active_operation <= op_readRegisterFile_8_write_1163;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1164;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(decodedInstr.imm = x"00000000")) then 
				active_operation <= op_readRegisterFile_8_write_1165;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (decodedInstr.imm = x"00000000")) then 
				active_operation <= op_readRegisterFile_8_write_1166;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1167;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and not(pc_reg = x"00000000")) then 
				active_operation <= op_readRegisterFile_8_write_1168;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT) and (pc_reg = x"00000000")) then 
				active_operation <= op_readRegisterFile_8_write_1169;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLT)) then 
				active_operation <= op_readRegisterFile_8_write_1170;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1171;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1172;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1173;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1174;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1175;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1176;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1177;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1178;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1179;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU)) then 
				active_operation <= op_readRegisterFile_8_write_1180;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1181;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU)) then 
				active_operation <= op_readRegisterFile_8_write_1182;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1183;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1184;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1185;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(pc_reg = x"00000000")) then 
				active_operation <= op_readRegisterFile_8_write_1186;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU) and (pc_reg = x"00000000")) then 
				active_operation <= op_readRegisterFile_8_write_1187;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1188;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLTU)) then 
				active_operation <= op_readRegisterFile_8_write_1189;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1190;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1191;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1192;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1193;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1194;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1195;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1196;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1197;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1198;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1199;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1200;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1201;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1202;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1203;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1204;
			elsif ((CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1205;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1206;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1207;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1208;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1209;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1210;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1211;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1212;
			elsif ((CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1213;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1214;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1215;
			end if;
		when st_writeBack_10 =>
			if (true) then 
				active_operation <= op_writeBack_10_write_1216;
			end if;
		end case;
	end process;

	-- Main process
	process (clk, rst)
	begin
		if (rst = '1') then
			decodedInstr.rd_addr <= x"00000000";
			decodedInstr.imm <= x"00000000";
			CtlToMem_port_sig.req <= ME_RD;
			br_en <= false;
			decodedInstr.instrType <= And_Instr;
			memoryAccess.req <= ME_RD;
			active_state <= st_fetch_4;
			CtlToMem_port_sig.addrIn <= x"00000000";
			MemToCtl_port_notify <= false;
			CtlToRegs_data.dst_data <= x"00000000";
			wb_sel <= WB_ALU;
			CtlToRegs_data.src1 <= x"00000000";
			ALUtoCtl_data.ALU_result <= x"00000000";
			CtlToALU_data.op2_sel <= OP_IMM;
			CtlToRegs_port_notify <= false;
			CtlToMem_port_sig.mask <= MT_W;
			fromMemoryData.loadedData <= x"00000000";
			CtlToALU_data.alu_fun <= ALU_ADD;
			CtlToALU_data.op1_sel <= OP_IMM;
			mem_en <= false;
			pc_next <= x"00000000";
			pc_reg <= x"00000000";
			memoryAccess.dataIn <= x"00000000";
			memoryAccess.addrIn <= x"00000000";
			RegsToCtl_data.contents2 <= x"00000000";
			CtlToDec_port_notify <= false;
			RegsToCtl_data.contents1 <= x"00000000";
			wb_en <= false;
			CtlToMem_port_notify <= true;
			memoryAccess.mask <= MT_W;
			CtlToRegs_data.dst <= x"00000000";
			CtlToRegs_data.src2 <= x"00000000";
			CtlToMem_port_sig.dataIn <= x"00000000";
			reg_rd_en <= false;
		elsif (clk = '1' and clk'event) then
			case active_operation is
			when op_wait_fetch_4 =>
				active_state <= st_fetch_4;
				CtlToMem_port_sig.addrIn <= memoryAccess.addrIn;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_sig.dataIn <= memoryAccess.dataIn;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
			when op_fetch_4_write_97 =>
				active_state <= st_fetch_5;
				CtlToMem_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				MemToCtl_port_notify <= true;
			when op_wait_fetch_5 =>
				active_state <= st_fetch_5;
				CtlToMem_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				MemToCtl_port_notify <= true;
			when op_fetch_5_read_98 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_99 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_100 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_101 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_102 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_103 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_104 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_105 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_106 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_107 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_108 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_109 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_110 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_111 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_112 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + DecToCtl_port_sig.imm;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_113 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_114 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_115 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_116 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_117 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_118 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_119 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_120 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_121 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_122 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_123 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_124 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_125 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_126 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_127 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - DecToCtl_port_sig.imm;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_128 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + pc_reg;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_129 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_130 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm - RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_131 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + DecToCtl_port_sig.imm;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_132 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg + RegsToCtl_data.contents2;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_133 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_134 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_135 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents2;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_136 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_137 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_138 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_139 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + DecToCtl_port_sig.imm;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_140 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_141 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_142 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_143 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_144 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_145 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_146 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_147 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_148 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_149 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_150 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_151 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_152 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and DecToCtl_port_sig.imm;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_153 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_154 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_155 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm and RegsToCtl_data.contents2;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_156 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_157 =>
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_158 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_159 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg - RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_160 =>
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_161 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= not(RegsToCtl_data.contents2) + 1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_162 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_163 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_164 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - DecToCtl_port_sig.imm;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_165 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + pc_reg;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_166 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_167 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm - RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_168 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + DecToCtl_port_sig.imm;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_169 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg + RegsToCtl_data.contents2;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_170 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_171 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_172 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents2;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_173 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_174 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_175 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_176 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + DecToCtl_port_sig.imm;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_177 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_178 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_179 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_180 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_181 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_182 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_183 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_184 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and pc_reg;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_185 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_186 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm or RegsToCtl_data.contents2;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_187 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_188 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm - pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_189 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_190 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg and RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_191 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= pc_reg - DecToCtl_port_sig.imm;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_192 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg + pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_193 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_194 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_195 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= not(DecToCtl_port_sig.imm) + 1;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_196 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_197 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_198 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_199 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and DecToCtl_port_sig.imm;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_200 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_201 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_202 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm and RegsToCtl_data.contents2;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_203 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_204 =>
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_205 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_206 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg - RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_207 =>
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_208 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= not(RegsToCtl_data.contents2) + 1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_209 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_210 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_211 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - DecToCtl_port_sig.imm;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_212 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + pc_reg;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_213 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_214 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm - RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_215 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + DecToCtl_port_sig.imm;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_216 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg + RegsToCtl_data.contents2;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_217 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_218 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_219 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents2;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_220 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_221 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_222 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_223 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or pc_reg;
			when op_fetch_5_read_224 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_225 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm xor RegsToCtl_data.contents2;
			when op_fetch_5_read_226 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_227 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm and pc_reg;
			when op_fetch_5_read_228 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_229 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= pc_reg or RegsToCtl_data.contents2;
			when op_fetch_5_read_230 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm and pc_reg;
			when op_fetch_5_read_231 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_232 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_233 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents2;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_234 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_235 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= not(pc_reg) + 1;
			when op_fetch_5_read_236 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_237 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_238 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_239 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and pc_reg;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_240 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_241 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm or RegsToCtl_data.contents2;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_242 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_243 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm - pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_244 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_245 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg and RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_246 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= pc_reg - DecToCtl_port_sig.imm;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_247 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg + pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_248 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_249 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_250 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= not(DecToCtl_port_sig.imm) + 1;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_251 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_252 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_253 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_254 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and DecToCtl_port_sig.imm;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_255 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_256 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_257 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm and RegsToCtl_data.contents2;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_258 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_259 =>
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_260 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_261 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg - RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_262 =>
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_263 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= not(RegsToCtl_data.contents2) + 1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_264 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_265 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_266 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_267 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_268 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_269 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_270 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm or pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_271 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_272 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= pc_reg xor RegsToCtl_data.contents2;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_273 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm or pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_274 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_275 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_276 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents2;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_277 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_278 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_279 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_280 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_281 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or pc_reg;
			when op_fetch_5_read_282 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_283 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm xor RegsToCtl_data.contents2;
			when op_fetch_5_read_284 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_285 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm and pc_reg;
			when op_fetch_5_read_286 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_287 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= pc_reg or RegsToCtl_data.contents2;
			when op_fetch_5_read_288 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm and pc_reg;
			when op_fetch_5_read_289 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_290 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_291 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents2;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_292 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_293 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= not(pc_reg) + 1;
			when op_fetch_5_read_294 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_295 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_296 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_297 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and pc_reg;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_298 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_299 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm or RegsToCtl_data.contents2;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_300 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_301 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm - pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_302 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_303 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg and RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_304 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= pc_reg - DecToCtl_port_sig.imm;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_305 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg + pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_306 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_307 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_308 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= not(DecToCtl_port_sig.imm) + 1;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_309 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_310 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_311 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_312 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_313 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_314 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_315 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_316 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_317 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_318 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm xor pc_reg;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_319 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_320 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm xor pc_reg;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_321 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_322 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_323 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_324 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_325 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_326 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_327 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_328 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_329 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_330 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_331 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm or pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_332 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_333 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= pc_reg xor RegsToCtl_data.contents2;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_334 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm or pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_335 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_336 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_337 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents2;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_338 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_339 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_340 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_341 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_342 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_343 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or pc_reg;
			when op_fetch_5_read_344 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_345 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm xor RegsToCtl_data.contents2;
			when op_fetch_5_read_346 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_347 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm and pc_reg;
			when op_fetch_5_read_348 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_349 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= pc_reg or RegsToCtl_data.contents2;
			when op_fetch_5_read_350 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm and pc_reg;
			when op_fetch_5_read_351 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_352 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_353 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents2;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_354 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_355 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= not(pc_reg) + 1;
			when op_fetch_5_read_356 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_357 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
			when op_fetch_5_read_358 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_359 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_360 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
			when op_fetch_5_read_361 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_362 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_363 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_364 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_365 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_366 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(DecToCtl_port_sig.imm, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_367 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_368 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_369 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_370 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_371 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_372 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_373 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_374 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_375 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_376 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_377 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_378 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_379 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_380 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_381 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_382 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_383 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm xor pc_reg;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_384 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_385 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm xor pc_reg;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_386 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_387 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_388 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_389 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_390 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_391 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_392 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_393 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_394 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_395 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_396 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_397 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_398 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm or pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_399 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_400 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= pc_reg xor RegsToCtl_data.contents2;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_401 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm or pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_402 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_403 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_404 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents2;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_405 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_406 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_407 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_408 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
			when op_fetch_5_read_409 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_410 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_411 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_412 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_413 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_414 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_415 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_416 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_417 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(DecToCtl_port_sig.imm, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_418 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_419 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_420 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_421 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_422 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_423 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_424 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_425 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_426 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_427 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_428 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_429 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_430 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_431 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
			when op_fetch_5_read_432 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_433 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_434 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
			when op_fetch_5_read_435 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_436 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_437 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_438 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_439 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_440 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(DecToCtl_port_sig.imm, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_441 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_442 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_443 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_444 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_445 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_446 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_447 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_448 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_449 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_450 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + RegsToCtl_data.contents2;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_451 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_452 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_453 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_454 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_455 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_456 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_457 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_458 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_459 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_460 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_461 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_462 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_463 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm xor pc_reg;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_464 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_465 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm xor pc_reg;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_466 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_467 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_468 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_469 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_470 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_471 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_472 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_473 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_474 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_475 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_476 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_477 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_478 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_479 =>
				ALUtoCtl_data.ALU_result <= shift_left(DecToCtl_port_sig.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_480 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_481 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_482 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_483 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_484 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_485 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_486 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_487 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_488 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_489 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_490 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_491 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_492 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_493 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_494 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_495 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
			when op_fetch_5_read_496 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_497 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_498 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_499 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_500 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_501 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_502 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_503 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_504 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(DecToCtl_port_sig.imm, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_505 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_506 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_507 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_508 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_509 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_510 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_511 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_512 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_513 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_514 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_515 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_516 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_517 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_518 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_519 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + DecToCtl_port_sig.imm;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_520 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_521 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_522 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_523 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_524 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_525 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
			when op_fetch_5_read_526 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_527 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_528 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
			when op_fetch_5_read_529 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_530 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_531 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_532 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_533 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_534 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(DecToCtl_port_sig.imm, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_535 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_536 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_537 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_538 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_539 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_540 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_541 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_542 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_543 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_544 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_545 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_546 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_547 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_548 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_549 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_550 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_551 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_552 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_553 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_554 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_555 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_556 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_557 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_558 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_559 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_560 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_561 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_562 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_563 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_564 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				CtlToALU_data.op1_sel <= OP_X;
				CtlToALU_data.op2_sel <= OP_X;
				wb_sel <= WB_PC4;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				CtlToALU_data.alu_fun <= ALU_X;
				reg_rd_en <= false;
			when op_fetch_5_read_565 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_566 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_567 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_568 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_569 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_570 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_571 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_572 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_573 =>
				ALUtoCtl_data.ALU_result <= shift_left(DecToCtl_port_sig.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_574 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_575 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_576 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_577 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_578 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_579 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_580 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_581 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_582 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_583 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_584 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_585 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_586 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_587 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_588 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_589 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_590 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - DecToCtl_port_sig.imm;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_591 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + pc_reg;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_592 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_593 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm - RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_594 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + DecToCtl_port_sig.imm;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_595 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg + RegsToCtl_data.contents2;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_596 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_597 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_598 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents2;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_599 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_600 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_601 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
			when op_fetch_5_read_602 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_603 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_604 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_605 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_606 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_607 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_608 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_609 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_610 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(DecToCtl_port_sig.imm, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_611 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_612 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_613 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_614 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_615 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_616 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_617 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_618 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_619 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_620 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_621 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_622 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_623 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_624 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_625 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_626 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_627 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_628 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_629 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_630 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_631 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_632 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_633 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_634 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_635 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_636 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_637 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_638 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_639 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_640 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_641 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_642 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_643 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_644 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_645 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_646 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_647 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_648 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_649 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_650 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_651 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_652 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_653 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_654 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_655 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_656 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_657 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_658 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and DecToCtl_port_sig.imm;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_659 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_660 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_661 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm and RegsToCtl_data.contents2;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_662 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_663 =>
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_664 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_665 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg - RegsToCtl_data.contents2;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_666 =>
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_667 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= not(RegsToCtl_data.contents2) + 1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_668 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_669 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_670 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_671 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_672 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_673 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_674 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_675 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_676 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_677 =>
				ALUtoCtl_data.ALU_result <= shift_left(DecToCtl_port_sig.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_678 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_679 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_680 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_681 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_682 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_683 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_684 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_685 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_686 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_687 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_688 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_689 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_690 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_691 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_692 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_693 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_694 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_695 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_696 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_697 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_698 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_699 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_700 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_701 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_702 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_703 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_704 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_705 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_706 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_707 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_708 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_709 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_710 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_711 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_712 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_713 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_714 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_715 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or DecToCtl_port_sig.imm;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_716 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and pc_reg;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_717 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_718 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm or RegsToCtl_data.contents2;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_719 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_720 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm - pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_721 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_722 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= pc_reg and RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_723 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= pc_reg - DecToCtl_port_sig.imm;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_724 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= pc_reg + pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_725 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_726 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_727 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= not(DecToCtl_port_sig.imm) + 1;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_728 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_729 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_730 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_731 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_732 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_733 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_734 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_735 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_736 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_737 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_738 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_739 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_740 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_741 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_742 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_743 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_744 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_745 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_746 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_747 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_748 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_749 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_750 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_751 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_752 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_753 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_754 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_755 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_756 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_757 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_758 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_759 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_760 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_761 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_762 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_763 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or pc_reg;
			when op_fetch_5_read_764 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_765 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm xor RegsToCtl_data.contents2;
			when op_fetch_5_read_766 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_767 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm and pc_reg;
			when op_fetch_5_read_768 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_769 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
				ALUtoCtl_data.ALU_result <= pc_reg or RegsToCtl_data.contents2;
			when op_fetch_5_read_770 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm and pc_reg;
			when op_fetch_5_read_771 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_772 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_773 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents2;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_774 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_775 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= not(pc_reg) + 1;
				reg_rd_en <= false;
			when op_fetch_5_read_776 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_777 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_778 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_779 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_780 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_781 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_782 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_783 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_784 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_785 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_786 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_787 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_788 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_789 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_790 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_791 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_792 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_793 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_794 =>
				CtlToALU_data.op1_sel <= OP_PC;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				CtlToALU_data.alu_fun <= ALU_ADD;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_795 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_796 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_797 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_798 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_799 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_800 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm or pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_801 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_802 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= pc_reg xor RegsToCtl_data.contents2;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_803 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm or pc_reg;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_804 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_805 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_806 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents2;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_807 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_808 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_809 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_810 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_811 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_812 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_813 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_814 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_815 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_816 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_817 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_818 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_819 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_820 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_821 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_822 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_823 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_824 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_825 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm xor pc_reg;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_826 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_827 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm xor pc_reg;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_828 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_829 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_830 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_831 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_832 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_833 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_834 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_835 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_836 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_837 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				reg_rd_en <= false;
			when op_fetch_5_read_838 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_839 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_840 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
			when op_fetch_5_read_841 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_842 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_843 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_844 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_845 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_846 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_left(DecToCtl_port_sig.imm, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_847 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_848 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_849 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_850 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_851 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_852 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_853 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_854 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_855 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_856 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				reg_rd_en <= false;
			when op_fetch_5_read_857 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_858 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_859 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_860 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_861 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_862 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_863 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_864 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_865 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_left(DecToCtl_port_sig.imm, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_866 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_867 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_868 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_869 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_870 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_871 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_872 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_873 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_874 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_875 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_876 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_877 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_878 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_879 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_880 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_881 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_882 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_883 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_884 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_885 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_886 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_887 =>
				ALUtoCtl_data.ALU_result <= shift_left(DecToCtl_port_sig.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_888 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_889 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_890 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_891 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_892 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_893 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_894 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_895 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_896 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_897 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_898 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_899 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_900 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_901 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_902 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_903 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_904 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_905 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_906 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_907 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_908 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_909 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_910 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_911 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_912 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_913 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_914 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_915 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_916 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_917 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_918 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_919 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_920 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_921 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_922 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_923 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_924 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_925 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_926 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= shift_right(DecToCtl_port_sig.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_927 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_928 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_929 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_930 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_931 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_932 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_933 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_934 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_935 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_936 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_937 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_938 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_939 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_940 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_941 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_942 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_943 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_944 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_945 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				ALUtoCtl_data.ALU_result <= pc_reg;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_946 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_947 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_948 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				CtlToALU_data.op1_sel <= OP_IMM;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				CtlToALU_data.alu_fun <= ALU_COPY1;
				CtlToALU_data.op2_sel <= OP_X;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_949 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_950 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_951 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_952 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_953 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_954 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToALU_data.alu_fun <= ALU_SLT;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_955 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				CtlToALU_data.op1_sel <= OP_X;
				CtlToALU_data.op2_sel <= OP_X;
				wb_sel <= WB_PC4;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				CtlToALU_data.alu_fun <= ALU_X;
			when op_fetch_5_read_956 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToALU_data.alu_fun <= ALU_SUB;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_957 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToALU_data.alu_fun <= ALU_SUB;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_958 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToALU_data.alu_fun <= ALU_SLTU;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_959 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_SLL;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_960 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToALU_data.alu_fun <= ALU_SUB;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_961 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_XOR;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_962 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				mem_en <= true;
				memoryAccess.mask <= MT_B;
				wb_sel <= WB_MEM;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				memoryAccess.req <= ME_RD;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_963 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToALU_data.alu_fun <= ALU_SLT;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_964 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToALU_data.alu_fun <= ALU_SLT;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_965 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_OR;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_966 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				mem_en <= true;
				wb_sel <= WB_MEM;
				memoryAccess.mask <= MT_H;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				memoryAccess.req <= ME_RD;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_967 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToALU_data.alu_fun <= ALU_SLTU;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_968 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToALU_data.alu_fun <= ALU_SLT;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_969 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_AND;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_970 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				mem_en <= true;
				wb_sel <= WB_MEM;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				memoryAccess.req <= ME_RD;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				memoryAccess.mask <= MT_W;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_971 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_XOR;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_972 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToALU_data.alu_fun <= ALU_SLTU;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_973 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_974 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				memoryAccess.req <= ME_WR;
				mem_en <= true;
				memoryAccess.mask <= MT_B;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_975 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_SLL;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_976 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				memoryAccess.mask <= MT_BU;
				mem_en <= true;
				wb_sel <= WB_MEM;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				memoryAccess.req <= ME_RD;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_977 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToALU_data.alu_fun <= ALU_SRL;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_978 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToALU_data.alu_fun <= ALU_SLTU;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_979 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				memoryAccess.req <= ME_WR;
				mem_en <= true;
				memoryAccess.mask <= MT_H;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_980 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				memoryAccess.req <= ME_WR;
				mem_en <= true;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_981 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToALU_data.alu_fun <= ALU_SRL;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_982 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				mem_en <= true;
				wb_sel <= WB_MEM;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				memoryAccess.req <= ME_RD;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				memoryAccess.mask <= MT_HU;
			when op_fetch_5_read_983 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.alu_fun <= ALU_SRA;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_984 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				memoryAccess.req <= ME_WR;
				mem_en <= true;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				memoryAccess.mask <= MT_W;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_985 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.alu_fun <= ALU_SRA;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_986 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_OR;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_987 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_988 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_AND;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_executeALU_2_read_0 =>
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				active_state <= st_executeALU_3;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1004 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1005 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1006 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1007 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 + RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1008 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1009 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1010 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1011 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1012 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1013 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 - RegsToCtl_port_sig.contents2;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1014 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 + decodedInstr.imm;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1015 =>
				ALUtoCtl_data.ALU_result <= decodedInstr.imm + RegsToCtl_port_sig.contents2;
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1016 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1017 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1018 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1019 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1020 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 and RegsToCtl_port_sig.contents2;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1021 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 - decodedInstr.imm;
			when op_readRegisterFile_8_write_1022 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 + pc_reg;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1023 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1024 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm - RegsToCtl_port_sig.contents2;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1025 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm + decodedInstr.imm;
			when op_readRegisterFile_8_write_1026 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg + RegsToCtl_port_sig.contents2;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1027 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1028 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1029 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents2;
			when op_readRegisterFile_8_write_1030 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1031 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1032 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 or RegsToCtl_port_sig.contents2;
			when op_readRegisterFile_8_write_1033 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 and decodedInstr.imm;
			when op_readRegisterFile_8_write_1034 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 - pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1035 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1036 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm and RegsToCtl_port_sig.contents2;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1037 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1038 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				ALUtoCtl_data.ALU_result <= pc_reg + decodedInstr.imm;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1039 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1040 =>
				ALUtoCtl_data.ALU_result <= pc_reg - RegsToCtl_port_sig.contents2;
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1041 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				ALUtoCtl_data.ALU_result <= pc_reg + decodedInstr.imm;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1042 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= not(RegsToCtl_port_sig.contents2) + 1;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1043 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1044 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 xor RegsToCtl_port_sig.contents2;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1045 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 or decodedInstr.imm;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1046 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 and pc_reg;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1047 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1048 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm or RegsToCtl_port_sig.contents2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1049 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1050 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm - pc_reg;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1051 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1052 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= pc_reg and RegsToCtl_port_sig.contents2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1053 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= pc_reg - decodedInstr.imm;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1054 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg + pc_reg;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1055 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1056 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1057 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= not(decodedInstr.imm) + 1;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1058 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1059 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1060 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 xor decodedInstr.imm;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1061 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 or pc_reg;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1062 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1063 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm xor RegsToCtl_port_sig.contents2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1064 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1065 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm and pc_reg;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1066 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1067 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= pc_reg or RegsToCtl_port_sig.contents2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1068 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm and pc_reg;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1069 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1070 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1071 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents2;
			when op_readRegisterFile_8_write_1072 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1073 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= not(pc_reg) + 1;
			when op_readRegisterFile_8_write_1074 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1075 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1076 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1077 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 xor pc_reg;
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1078 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1079 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1080 =>
				ALUtoCtl_data.ALU_result <= decodedInstr.imm or pc_reg;
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1081 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1082 =>
				ALUtoCtl_data.ALU_result <= pc_reg xor RegsToCtl_port_sig.contents2;
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1083 =>
				ALUtoCtl_data.ALU_result <= decodedInstr.imm or pc_reg;
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1084 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1085 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1086 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents2;
			when op_readRegisterFile_8_write_1087 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1088 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1089 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1090 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1091 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1092 =>
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_port_sig.contents1, to_integer(RegsToCtl_port_sig.contents2 and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1093 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1094 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1095 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1096 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1097 =>
				ALUtoCtl_data.ALU_result <= decodedInstr.imm xor pc_reg;
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1098 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1099 =>
				ALUtoCtl_data.ALU_result <= decodedInstr.imm xor pc_reg;
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1100 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1101 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1102 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1103 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1104 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1105 =>
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_port_sig.contents1, to_integer(RegsToCtl_port_sig.contents2 and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1106 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1107 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1108 =>
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_port_sig.contents1, to_integer(decodedInstr.imm and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1109 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1110 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1111 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1112 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1113 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1114 =>
				ALUtoCtl_data.ALU_result <= shift_left(decodedInstr.imm, to_integer(RegsToCtl_port_sig.contents2 and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1115 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1116 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1117 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1118 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1119 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1120 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1121 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1122 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1123 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1124 =>
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_port_sig.contents1, to_integer(RegsToCtl_port_sig.contents2 and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1125 =>
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_port_sig.contents1, to_integer(decodedInstr.imm and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1126 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1127 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1128 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_port_sig.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
			when op_readRegisterFile_8_write_1129 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1130 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1131 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(decodedInstr.imm, to_integer(RegsToCtl_port_sig.contents2 and to_unsigned(31, 32)));
			when op_readRegisterFile_8_write_1132 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1133 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(decodedInstr.imm, to_integer(decodedInstr.imm and to_unsigned(31, 32)));
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1134 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1135 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1136 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1137 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1138 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1139 =>
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(RegsToCtl_port_sig.contents2 and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1140 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1141 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1142 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1143 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1144 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1145 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1146 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1147 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1148 =>
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_port_sig.contents1, to_integer(decodedInstr.imm and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1149 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_port_sig.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1150 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1151 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(decodedInstr.imm, to_integer(RegsToCtl_port_sig.contents2 and to_unsigned(31, 32)));
			when op_readRegisterFile_8_write_1152 =>
				ALUtoCtl_data.ALU_result <= shift_right(decodedInstr.imm, to_integer(decodedInstr.imm and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1153 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1154 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1155 =>
				ALUtoCtl_data.ALU_result <= shift_left(decodedInstr.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1156 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1157 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1158 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(RegsToCtl_port_sig.contents2 and to_unsigned(31, 32)));
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1159 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1160 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1161 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(decodedInstr.imm and to_unsigned(31, 32)));
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1162 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1163 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1164 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1165 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1166 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1167 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1168 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1169 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1170 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1171 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1172 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_port_sig.contents1, to_integer(pc_reg and to_unsigned(31, 32)));
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1173 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1174 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1175 =>
				ALUtoCtl_data.ALU_result <= shift_right(decodedInstr.imm, to_integer(decodedInstr.imm and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1176 =>
				ALUtoCtl_data.ALU_result <= shift_right(decodedInstr.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1177 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1178 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(RegsToCtl_port_sig.contents2 and to_unsigned(31, 32)));
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1179 =>
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(decodedInstr.imm and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1180 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1181 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_left(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1182 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1183 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1184 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1185 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1186 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1187 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1188 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1189 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1190 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1191 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1192 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1193 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1194 =>
				ALUtoCtl_data.ALU_result <= shift_right(decodedInstr.imm, to_integer(pc_reg and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1195 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1196 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1197 =>
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(decodedInstr.imm and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1198 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
			when op_readRegisterFile_8_write_1199 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1200 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1201 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1202 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1203 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1204 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1205 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= decodedInstr.imm;
			when op_readRegisterFile_8_write_1206 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1207 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(pc_reg, to_integer(pc_reg and to_unsigned(31, 32)));
			when op_readRegisterFile_8_write_1208 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1209 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1210 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1211 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1212 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1213 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= pc_reg;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1214 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1215 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_executeALU_3_read_1 =>
				memoryAccess.addrIn <= x"00000004" + pc_reg;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				pc_reg <= x"00000004" + pc_reg;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= x"00000004" + pc_reg;
			when op_executeALU_3_read_2 =>
				memoryAccess.addrIn <= x"00000004" + pc_reg;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				pc_reg <= x"00000004" + pc_reg;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= x"00000004" + pc_reg;
			when op_executeALU_3_read_3 =>
				memoryAccess.addrIn <= x"00000004" + pc_reg;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				pc_reg <= x"00000004" + pc_reg;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= x"00000004" + pc_reg;
			when op_executeALU_3_read_4 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_5 =>
				memoryAccess.addrIn <= x"00000004" + pc_reg;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				pc_reg <= x"00000004" + pc_reg;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= x"00000004" + pc_reg;
			when op_executeALU_3_read_6 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_7 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_8 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_9 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_10 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_11 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_12 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_13 =>
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				memoryAccess.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				pc_reg <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_14 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_15 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_16 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_17 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_18 =>
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				memoryAccess.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				pc_reg <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_19 =>
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				memoryAccess.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				pc_reg <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_20 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_21 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_22 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_23 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_24 =>
				memoryAccess.addrIn <= x"00000004" + pc_reg;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				pc_reg <= x"00000004" + pc_reg;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= x"00000004" + pc_reg;
			when op_executeALU_3_read_25 =>
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				memoryAccess.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				pc_reg <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_26 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_27 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_28 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_29 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_30 =>
				memoryAccess.addrIn <= x"00000004" + pc_reg;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				pc_reg <= x"00000004" + pc_reg;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= x"00000004" + pc_reg;
			when op_executeALU_3_read_31 =>
				memoryAccess.addrIn <= x"00000004" + pc_reg;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				pc_reg <= x"00000004" + pc_reg;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= x"00000004" + pc_reg;
			when op_executeALU_3_read_32 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_33 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_34 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_35 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_36 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_37 =>
				memoryAccess.addrIn <= x"00000004" + pc_reg;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				pc_reg <= x"00000004" + pc_reg;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= x"00000004" + pc_reg;
			when op_executeALU_3_read_38 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_39 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_40 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_41 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_42 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_43 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_44 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_45 =>
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				memoryAccess.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				pc_reg <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_46 =>
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				memoryAccess.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				pc_reg <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_47 =>
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				memoryAccess.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				pc_reg <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_48 =>
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				memoryAccess.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				pc_reg <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_49 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_50 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				pc_next <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_51 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				pc_next <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_52 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				pc_next <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_53 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_54 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				pc_next <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_55 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				pc_next <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_56 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_57 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				pc_next <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_58 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				pc_next <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_59 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				pc_next <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_60 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_61 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= x"00000004" + pc_reg;
			when op_executeALU_3_read_62 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= x"00000004" + pc_reg;
			when op_executeALU_3_read_63 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_64 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= x"00000004" + pc_reg;
			when op_executeALU_3_read_65 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_66 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_67 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_68 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_69 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_70 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_71 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_72 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_73 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_74 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_75 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_76 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_77 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_78 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= x"00000004" + pc_reg;
			when op_executeALU_3_read_79 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_80 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_81 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_82 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_83 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= x"00000004" + pc_reg;
			when op_executeALU_3_read_84 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_85 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_86 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_87 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_88 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= x"00000004" + pc_reg;
			when op_executeALU_3_read_89 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_90 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_91 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_92 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_93 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_94 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_95 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_96 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_memoryOperation_6_write_989 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_memoryOperation_6_write_990 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_memoryOperation_6_write_991 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_memoryOperation_6_write_992 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_wait_memoryOperation_6 =>
				CtlToMem_port_sig.addrIn <= memoryAccess.addrIn;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_sig.dataIn <= memoryAccess.dataIn;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
			when op_memoryOperation_6_write_993 =>
				CtlToMem_port_notify <= false;
				active_state <= st_memoryOperation_7;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				MemToCtl_port_notify <= true;
			when op_memoryOperation_6_write_994 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
			when op_memoryOperation_6_write_995 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst_data <= fromMemoryData.loadedData;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
			when op_memoryOperation_6_write_996 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
			when op_writeBack_10_write_1216 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_memoryOperation_7_read_997 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_memoryOperation_7_read_998 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_memoryOperation_7_read_999 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_memoryOperation_7_read_1000 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_wait_memoryOperation_7 =>
				CtlToMem_port_notify <= false;
				active_state <= st_memoryOperation_7;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				MemToCtl_port_notify <= true;
			when op_memoryOperation_7_read_1001 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
			when op_memoryOperation_7_read_1002 =>
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToRegs_data.dst_data <= MemToCtl_port_sig.loadedData;
				CtlToRegs_port_sig.dst_data <= MemToCtl_port_sig.loadedData;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
			when op_memoryOperation_7_read_1003 =>
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
			end case;
		end if;
	end process;

	-- Assigning state signals that are used by ITL properties for OneSpin
	executeALU_2 <= active_state = st_executeALU_2;
	executeALU_3 <= active_state = st_executeALU_3;
	fetch_4 <= active_state = st_fetch_4;
	fetch_5 <= active_state = st_fetch_5;
	memoryOperation_6 <= active_state = st_memoryOperation_6;
	memoryOperation_7 <= active_state = st_memoryOperation_7;
	readRegisterFile_8 <= active_state = st_readRegisterFile_8;
	writeBack_10 <= active_state = st_writeBack_10;

end ISA_arch;

