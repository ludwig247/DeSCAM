library ieee;
use IEEE.numeric_std.all;

package TestBasic7_types is
end package TestBasic7_types;