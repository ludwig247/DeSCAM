package testarray2_types;

	 import top_level_types::*;
endpackage