library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestArray3_types is
end package TestArray3_types;