package testbasic14_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic14_SECTIONS;

endpackage
