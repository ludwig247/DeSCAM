library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package Component1_types is
-- No local datatypes implemented!


end package Component1_types;