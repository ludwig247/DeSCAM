package testbasic4_types;

	 import top_level_types::*;
endpackage