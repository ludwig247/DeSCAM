library ieee;
use IEEE.numeric_std.all;

package TestBasic6_types is
type TestBasic6_SECTIONS is (run);
end package TestBasic6_types;
