package testarray03_types;

	import top_level_types::*;
// No local datatypes implemented!


endpackage