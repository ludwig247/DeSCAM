library ieee;
use IEEE.numeric_std.all;

package TestBasic8_types is
end package TestBasic8_types;