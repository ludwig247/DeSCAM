package testmasterslave7_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave7_SECTIONS;

endpackage
