package testmasterslave5_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave5_SECTIONS;

endpackage
