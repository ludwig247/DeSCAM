library ieee;
use IEEE.numeric_std.all;

package TestBasic16_types is
type TestBasic16_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic16_types;
