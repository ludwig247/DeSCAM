library ieee;
use IEEE.numeric_std.all;

package TestBasic7_types is
type TestBasic7_SECTIONS is (run);
end package TestBasic7_types;
