package testbasic7_types;

	typedef enum logic {
		run
	} TestBasic7_SECTIONS;

endpackage
