library ieee;
use IEEE.numeric_std.all;

package TestBasic5_types is
type TestBasic5_SECTIONS is (run);
end package TestBasic5_types;
