package testbasic22_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic22_SECTIONS;

endpackage
