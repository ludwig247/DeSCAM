package testbasic20_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic20_SECTIONS;

	typedef enum logic [1:0] {
		green,
		red,
		yellow
	} color_t;

endpackage
