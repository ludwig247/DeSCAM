library ieee;
use IEEE.numeric_std.all;
use work.SCAM_Model_types.all;

package TestFunction1_types is
end package TestFunction1_types;