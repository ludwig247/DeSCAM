package testmasterslave11_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave11_SECTIONS;

endpackage
