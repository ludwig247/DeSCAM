library ieee;
use IEEE.numeric_std.all;

package TestBasic9_types is
type TestBasic9_SECTIONS is (run);
end package TestBasic9_types;
