package testbasic9_types;

	import scam_model_types::*;
endpackage