package testbasic8_types;

	import scam_model_types::*;
endpackage