package testbasic23_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic23_SECTIONS;

endpackage
