library ieee;
use IEEE.numeric_std.all;

package TestBasic19_types is
type TestBasic19_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic19_types;
