library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package Bus_new_types is
-- No local datatypes implemented!


end package Bus_new_types;