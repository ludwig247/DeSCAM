library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave13_types is
type TestMasterSlave13_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave13_types;
