library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestBasic01_types is
type Phases is (SECTION_A, SECTION_B);
end package TestBasic01_types;