library ieee;
use IEEE.numeric_std.all;

package TestBasic4_types is
end package TestBasic4_types;