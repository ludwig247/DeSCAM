package testmasterslave12_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave12_SECTIONS;

endpackage
