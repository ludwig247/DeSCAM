package testbasic1_types;

	typedef enum logic {
		section_a,
		section_b
	} Sections;

endpackage