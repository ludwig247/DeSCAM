-- External data type definition package
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package SCAM_Model_types is
	type ME_MaskType is (MT_B, MT_BU, MT_H, MT_HU, MT_W, MT_X);
	type ME_AccessType is (ME_RD, ME_WR, ME_X);
	type CUtoME_IF is record
		addrIn: unsigned(31 downto 0);
		dataIn: unsigned(31 downto 0);
		mask: ME_MaskType;
		req: ME_AccessType;
	end record;
	type AccessType_Reg is (REG_RD, REG_WR);
	type CtlToRegs_IF is record
		dst: unsigned(31 downto 0);
		dst_data: unsigned(31 downto 0);
		req: AccessType_Reg;
		src1: unsigned(31 downto 0);
		src2: unsigned(31 downto 0);
	end record;
	type EncType is (B, Error_Type, I, J, R, S, U);
	type InstrType is (And_Instr, Or_Instr, Unknown, Xor_Instr, add, addI, andI, auipc, beq, bge, bgeu, blt, bltu, bne, jal, jalr, lb, lbu, lh, lhu, lui, lw, orI, sb, sh, sllI, sll_Instr, slt, sltI, sltIu, sltu, sraI, sra_Instr, srlI, srl_Instr, sub, sw, xorI);
	type DecodedInstr is record
		encType: EncType;
		imm: unsigned(31 downto 0);
		instrType: InstrType;
		rd_addr: unsigned(31 downto 0);
		rs1_addr: unsigned(31 downto 0);
		rs2_addr: unsigned(31 downto 0);
	end record;
	type MEtoCU_IF is record
		loadedData: unsigned(31 downto 0);
	end record;
	type RegsToCtl_IF is record
		contents1: unsigned(31 downto 0);
		contents2: unsigned(31 downto 0);
	end record;
end package SCAM_Model_types;



library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.SCAM_Model_types.all;

entity ISA is
port(	
	CtlToDec_port_sig: out unsigned(31 downto 0);
	CtlToDec_port_notify: out boolean;
	CtlToMem_port_sig: out CUtoME_IF;
	CtlToMem_port_sync: in boolean;
	CtlToMem_port_notify: out boolean;
	CtlToRegs_port_sig: out CtlToRegs_IF;
	CtlToRegs_port_notify: out boolean;
	DecToCtl_port_sig: in DecodedInstr;
	MemToCtl_port_sig: in MEtoCU_IF;
	MemToCtl_port_sync: in boolean;
	MemToCtl_port_notify: out boolean;
	RegsToCtl_port_sig: in RegsToCtl_IF;
	dummy_port_sig: in boolean;
	clk: in std_logic;
	rst: in std_logic
);
end ISA;

architecture ISA_arch of ISA is
	-- Define internal data types
	type ISA_operation_t is (op_wait_fetch_4, op_fetch_4_write_97, op_wait_fetch_5, op_fetch_5_read_98, op_fetch_5_read_101, op_fetch_5_read_102, op_fetch_5_read_110, op_fetch_5_read_111, op_fetch_5_read_112, op_fetch_5_read_118, op_fetch_5_read_126, op_fetch_5_read_131, op_fetch_5_read_137, op_fetch_5_read_138, op_fetch_5_read_139, op_fetch_5_read_145, op_fetch_5_read_151, op_fetch_5_read_152, op_fetch_5_read_160, op_fetch_5_read_163, op_fetch_5_read_168, op_fetch_5_read_174, op_fetch_5_read_175, op_fetch_5_read_176, op_fetch_5_read_182, op_fetch_5_read_183, op_fetch_5_read_198, op_fetch_5_read_199, op_fetch_5_read_207, op_fetch_5_read_210, op_fetch_5_read_215, op_fetch_5_read_221, op_fetch_5_read_222, op_fetch_5_read_237, op_fetch_5_read_238, op_fetch_5_read_253, op_fetch_5_read_254, op_fetch_5_read_262, op_fetch_5_read_265, op_fetch_5_read_266, op_fetch_5_read_280, op_fetch_5_read_295, op_fetch_5_read_296, op_fetch_5_read_311, op_fetch_5_read_312, op_fetch_5_read_313, op_fetch_5_read_314, op_fetch_5_read_315, op_fetch_5_read_326, op_fetch_5_read_327, op_fetch_5_read_341, op_fetch_5_read_342, op_fetch_5_read_357, op_fetch_5_read_358, op_fetch_5_read_359, op_fetch_5_read_360, op_fetch_5_read_376, op_fetch_5_read_377, op_fetch_5_read_378, op_fetch_5_read_379, op_fetch_5_read_380, op_fetch_5_read_393, op_fetch_5_read_394, op_fetch_5_read_408, op_fetch_5_read_409, op_fetch_5_read_431, op_fetch_5_read_432, op_fetch_5_read_433, op_fetch_5_read_434, op_fetch_5_read_450, op_fetch_5_read_456, op_fetch_5_read_457, op_fetch_5_read_458, op_fetch_5_read_459, op_fetch_5_read_460, op_fetch_5_read_471, op_fetch_5_read_472, op_fetch_5_read_495, op_fetch_5_read_496, op_fetch_5_read_518, op_fetch_5_read_519, op_fetch_5_read_525, op_fetch_5_read_526, op_fetch_5_read_527, op_fetch_5_read_528, op_fetch_5_read_564, op_fetch_5_read_565, op_fetch_5_read_566, op_fetch_5_read_589, op_fetch_5_read_594, op_fetch_5_read_600, op_fetch_5_read_601, op_fetch_5_read_602, op_fetch_5_read_657, op_fetch_5_read_658, op_fetch_5_read_666, op_fetch_5_read_669, op_fetch_5_read_670, op_fetch_5_read_694, op_fetch_5_read_714, op_fetch_5_read_715, op_fetch_5_read_755, op_fetch_5_read_762, op_fetch_5_read_794, op_fetch_5_read_795, op_fetch_5_read_796, op_fetch_5_read_811, op_fetch_5_read_818, op_fetch_5_read_819, op_fetch_5_read_820, op_fetch_5_read_821, op_fetch_5_read_822, op_fetch_5_read_837, op_fetch_5_read_838, op_fetch_5_read_839, op_fetch_5_read_840, op_fetch_5_read_856, op_fetch_5_read_857, op_fetch_5_read_879, op_fetch_5_read_880, op_fetch_5_read_937, op_fetch_5_read_948, op_fetch_5_read_949, op_fetch_5_read_950, op_fetch_5_read_951, op_fetch_5_read_952, op_fetch_5_read_953, op_fetch_5_read_954, op_fetch_5_read_955, op_fetch_5_read_956, op_fetch_5_read_957, op_fetch_5_read_958, op_fetch_5_read_959, op_fetch_5_read_960, op_fetch_5_read_961, op_fetch_5_read_962, op_fetch_5_read_963, op_fetch_5_read_964, op_fetch_5_read_965, op_fetch_5_read_966, op_fetch_5_read_967, op_fetch_5_read_968, op_fetch_5_read_969, op_fetch_5_read_970, op_fetch_5_read_971, op_fetch_5_read_972, op_fetch_5_read_973, op_fetch_5_read_974, op_fetch_5_read_975, op_fetch_5_read_976, op_fetch_5_read_977, op_fetch_5_read_978, op_fetch_5_read_979, op_fetch_5_read_980, op_fetch_5_read_981, op_fetch_5_read_982, op_fetch_5_read_983, op_fetch_5_read_984, op_fetch_5_read_985, op_fetch_5_read_986, op_fetch_5_read_987, op_fetch_5_read_988, op_executeALU_2_read_0, op_readRegisterFile_8_write_1004, op_readRegisterFile_8_write_1007, op_readRegisterFile_8_write_1013, op_readRegisterFile_8_write_1014, op_readRegisterFile_8_write_1020, op_readRegisterFile_8_write_1031, op_readRegisterFile_8_write_1032, op_readRegisterFile_8_write_1033, op_readRegisterFile_8_write_1044, op_readRegisterFile_8_write_1045, op_readRegisterFile_8_write_1060, op_readRegisterFile_8_write_1075, op_readRegisterFile_8_write_1076, op_readRegisterFile_8_write_1090, op_readRegisterFile_8_write_1091, op_readRegisterFile_8_write_1092, op_readRegisterFile_8_write_1093, op_readRegisterFile_8_write_1094, op_readRegisterFile_8_write_1105, op_readRegisterFile_8_write_1106, op_readRegisterFile_8_write_1107, op_readRegisterFile_8_write_1108, op_readRegisterFile_8_write_1124, op_readRegisterFile_8_write_1125, op_readRegisterFile_8_write_1147, op_readRegisterFile_8_write_1148, op_executeALU_3_read_1, op_executeALU_3_read_4, op_executeALU_3_read_5, op_executeALU_3_read_10, op_executeALU_3_read_12, op_executeALU_3_read_13, op_executeALU_3_read_16, op_executeALU_3_read_22, op_executeALU_3_read_25, op_executeALU_3_read_28, op_executeALU_3_read_31, op_executeALU_3_read_34, op_executeALU_3_read_40, op_executeALU_3_read_42, op_executeALU_3_read_47, op_executeALU_3_read_49, op_executeALU_3_read_50, op_executeALU_3_read_53, op_executeALU_3_read_61, op_executeALU_3_read_63, op_executeALU_3_read_64, op_executeALU_3_read_69, op_executeALU_3_read_70, op_executeALU_3_read_79, op_memoryOperation_6_write_991, op_wait_memoryOperation_6, op_memoryOperation_6_write_993, op_writeBack_10_write_1216, op_memoryOperation_7_read_998, op_memoryOperation_7_read_999, op_wait_memoryOperation_7, op_memoryOperation_7_read_1002, op_memoryOperation_7_read_1003);
	type ISA_state_t is (st_executeALU_2, st_executeALU_3, st_fetch_4, st_fetch_5, st_memoryOperation_6, st_memoryOperation_7, st_readRegisterFile_8, st_writeBack_10);
	type ALUtoCtl_IF is record
		ALU_result: unsigned(31 downto 0);
	end record;
	type ALU_function is (ALU_ADD, ALU_AND, ALU_COPY1, ALU_OR, ALU_SLL, ALU_SLT, ALU_SLTU, ALU_SRA, ALU_SRL, ALU_SUB, ALU_X, ALU_XOR);
	type ALUopType is (OP_IMM, OP_PC, OP_REG, OP_X);
	type CtlToALU_IF is record
		alu_fun: ALU_function;
		imm: unsigned(31 downto 0);
		op1_sel: ALUopType;
		op2_sel: ALUopType;
		pc_reg: unsigned(31 downto 0);
		reg1_contents: unsigned(31 downto 0);
		reg2_contents: unsigned(31 downto 0);
	end record;
	type WBselType is (WB_ALU, WB_MEM, WB_PC4, WB_X);

	-- Declare signals
	signal active_state: ISA_state_t;
	signal active_operation: ISA_operation_t;
	signal ALUtoCtl_data: ALUtoCtl_IF;
	signal CtlToALU_data: CtlToALU_IF;
	signal CtlToRegs_data: CtlToRegs_IF;
	signal RegsToCtl_data: RegsToCtl_IF;
	signal br_en: boolean;
	signal decodedInstr: DecodedInstr;
	signal fromMemoryData: MEtoCU_IF;
	signal mem_en: boolean;
	signal memoryAccess: CUtoME_IF;
	signal pc_next: unsigned(31 downto 0);
	signal pc_reg: unsigned(31 downto 0);
	signal reg_rd_en: boolean;
	signal wb_en: boolean;
	signal wb_sel: WBselType;

	-- Declare state signals that are used by ITL properties for OneSpin
	signal executeALU_2: boolean;
	signal executeALU_3: boolean;
	signal fetch_4: boolean;
	signal fetch_5: boolean;
	signal memoryOperation_6: boolean;
	signal memoryOperation_7: boolean;
	signal readRegisterFile_8: boolean;
	signal writeBack_10: boolean;


begin
	-- Combinational logic that selects current operation
	process (active_state, CtlToMem_port_sync, MemToCtl_port_sync, DecToCtl_port_sig.instrType, DecToCtl_port_sig.imm, RegsToCtl_port_sig.contents2, RegsToCtl_port_sig.contents1, DecToCtl_port_sig.encType, memoryAccess.req, pc_reg, ALUtoCtl_data.ALU_result, mem_en, CtlToALU_data.alu_fun, wb_sel, CtlToALU_data.op1_sel, CtlToALU_data.op2_sel, decodedInstr.instrType, decodedInstr.rd_addr, decodedInstr.imm, br_en, RegsToCtl_data.contents2, reg_rd_en, wb_en, RegsToCtl_data.contents1)
	begin
	active_operation <= op_wait_fetch_4;
		case active_state is
		when st_executeALU_2 =>
			if (true) then 
				active_operation <= op_executeALU_2_read_0;
			end if;
		when st_executeALU_3 =>
			if (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_1;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_4;
			elsif (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_5;
			elsif (br_en and (decodedInstr.instrType = beq) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_10;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_12;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_ALU) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_13;
			elsif (br_en and (decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000") and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4)) then 
				active_operation <= op_executeALU_3_read_16;
			elsif (br_en and (decodedInstr.instrType = blt) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_22;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_PC4) and not(wb_en and not(decodedInstr.rd_addr = x"00000000"))) then 
				active_operation <= op_executeALU_3_read_25;
			elsif (br_en and (decodedInstr.instrType = bge) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_28;
			elsif (br_en and not((decodedInstr.instrType = beq) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bne) and not(ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = blt) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bge) and (ALUtoCtl_data.ALU_result = x"00000000")) and not((decodedInstr.instrType = bltu) and (ALUtoCtl_data.ALU_result = x"00000001")) and not((decodedInstr.instrType = bgeu) and (ALUtoCtl_data.ALU_result = x"00000000")) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4)) then 
				active_operation <= op_executeALU_3_read_31;
			elsif (br_en and (decodedInstr.instrType = bltu) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and (ALUtoCtl_data.ALU_result = x"00000001")) then 
				active_operation <= op_executeALU_3_read_34;
			elsif (br_en and (decodedInstr.instrType = bgeu) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and (ALUtoCtl_data.ALU_result = x"00000000")) then 
				active_operation <= op_executeALU_3_read_40;
			elsif (br_en and (decodedInstr.instrType = jal) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4)) then 
				active_operation <= op_executeALU_3_read_42;
			elsif (br_en and (decodedInstr.instrType = jalr) and not(mem_en) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4)) then 
				active_operation <= op_executeALU_3_read_47;
			elsif (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and mem_en) then 
				active_operation <= op_executeALU_3_read_49;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and mem_en) then 
				active_operation <= op_executeALU_3_read_50;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and mem_en) then 
				active_operation <= op_executeALU_3_read_53;
			elsif (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_61;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_63;
			elsif (not(br_en) and not(decodedInstr.instrType = jal) and not(decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_64;
			elsif (not(br_en) and (decodedInstr.instrType = jal) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_69;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_ALU) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_70;
			elsif (not(br_en) and (decodedInstr.instrType = jalr) and not(mem_en) and (wb_sel = WB_PC4) and wb_en and not(decodedInstr.rd_addr = x"00000000")) then 
				active_operation <= op_executeALU_3_read_79;
			end if;
		when st_fetch_4 =>
			if (not(CtlToMem_port_sync)) then 
				active_operation <= op_wait_fetch_4;
			elsif (CtlToMem_port_sync) then 
				active_operation <= op_fetch_4_write_97;
			end if;
		when st_fetch_5 =>
			if (not(MemToCtl_port_sync)) then 
				active_operation <= op_wait_fetch_5;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_98;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_101;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_102;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_110;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_111;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_112;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_118;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_126;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_131;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_137;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_138;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_139;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_145;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_151;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_152;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_160;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_163;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_168;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_174;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_175;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_176;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_182;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_183;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_198;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_199;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_207;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_210;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_215;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_221;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_222;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_237;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_238;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_253;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_254;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_262;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_265;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_266;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_280;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_295;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_296;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_311;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_312;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_313;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_314;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_315;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_326;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_327;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_341;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_342;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_357;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_358;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_359;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_360;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_376;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_377;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_378;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_379;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_380;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_393;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_394;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_408;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_409;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_431;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_432;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_433;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_434;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_450;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_456;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_457;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_458;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_459;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_460;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_471;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_472;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_495;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_496;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_518;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_519;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_525;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_526;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_527;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_528;
			elsif ((DecToCtl_port_sig.encType = J) and (DecToCtl_port_sig.instrType = jal) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_564;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_565;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_566;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_589;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_594;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_600;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_601;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_602;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_657;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_658;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_PC) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_666;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_669;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_670;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_694;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_714;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_715;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_755;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_762;
			elsif ((DecToCtl_port_sig.encType = U) and (DecToCtl_port_sig.instrType = auipc) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_794;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_795;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_796;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and not(reg_rd_en) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_811;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_818;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_data.contents2 <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_819;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_820;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_821;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_822;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_837;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_838;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (DecToCtl_port_sig.imm <= RegsToCtl_data.contents1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_839;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_840;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_856;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_857;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_879;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_880;
			elsif ((DecToCtl_port_sig.encType = U) and not(DecToCtl_port_sig.instrType = lui) and not(DecToCtl_port_sig.instrType = auipc) and (CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_COPY1) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_937;
			elsif ((DecToCtl_port_sig.encType = U) and (DecToCtl_port_sig.instrType = lui) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_948;
			elsif ((DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.instrType = addI) and not(DecToCtl_port_sig.instrType = sltI) and not(DecToCtl_port_sig.instrType = sltIu) and not(DecToCtl_port_sig.instrType = xorI) and not(DecToCtl_port_sig.instrType = orI) and not(DecToCtl_port_sig.instrType = andI) and not(DecToCtl_port_sig.instrType = sllI) and not(DecToCtl_port_sig.instrType = srlI) and not(DecToCtl_port_sig.instrType = sraI) and not(DecToCtl_port_sig.instrType = lb) and not(DecToCtl_port_sig.instrType = lh) and not(DecToCtl_port_sig.instrType = lw) and not(DecToCtl_port_sig.instrType = lbu) and not(DecToCtl_port_sig.instrType = lhu) and not(DecToCtl_port_sig.instrType = jalr) and reg_rd_en and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_949;
			elsif ((DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.instrType = jal) and reg_rd_en and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_950;
			elsif (not(DecToCtl_port_sig.encType = I) and not(DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.encType = J) and not(DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.encType = U) and reg_rd_en and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_951;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = addI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_952;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = add) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_953;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = sltI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_954;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = jalr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_955;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = sub) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_956;
			elsif ((DecToCtl_port_sig.encType = B) and (DecToCtl_port_sig.instrType = beq) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_957;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = sltIu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_958;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = sll_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_959;
			elsif ((DecToCtl_port_sig.encType = B) and (DecToCtl_port_sig.instrType = bne) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_960;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = xorI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_961;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = lb) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_962;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = slt) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_963;
			elsif ((DecToCtl_port_sig.encType = B) and (DecToCtl_port_sig.instrType = blt) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_964;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = orI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_965;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = lh) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_966;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = sltu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_967;
			elsif ((DecToCtl_port_sig.encType = B) and (DecToCtl_port_sig.instrType = bge) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_968;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = andI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_969;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = lw) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_970;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = Xor_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_971;
			elsif ((DecToCtl_port_sig.encType = B) and (DecToCtl_port_sig.instrType = bltu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_972;
			elsif ((DecToCtl_port_sig.encType = B) and not(DecToCtl_port_sig.instrType = beq) and not(DecToCtl_port_sig.instrType = bne) and not(DecToCtl_port_sig.instrType = blt) and not(DecToCtl_port_sig.instrType = bge) and not(DecToCtl_port_sig.instrType = bltu) and not(DecToCtl_port_sig.instrType = bgeu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_973;
			elsif ((DecToCtl_port_sig.encType = S) and (DecToCtl_port_sig.instrType = sb) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_974;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = sllI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_975;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = lbu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_976;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = srl_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_977;
			elsif ((DecToCtl_port_sig.encType = B) and (DecToCtl_port_sig.instrType = bgeu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_978;
			elsif ((DecToCtl_port_sig.encType = S) and (DecToCtl_port_sig.instrType = sh) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_979;
			elsif ((DecToCtl_port_sig.encType = S) and not(DecToCtl_port_sig.instrType = sb) and not(DecToCtl_port_sig.instrType = sh) and not(DecToCtl_port_sig.instrType = sw) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_980;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = srlI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_981;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = lhu) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_982;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = sra_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_983;
			elsif ((DecToCtl_port_sig.encType = S) and (DecToCtl_port_sig.instrType = sw) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_984;
			elsif ((DecToCtl_port_sig.encType = I) and (DecToCtl_port_sig.instrType = sraI) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_985;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = Or_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_986;
			elsif ((DecToCtl_port_sig.encType = R) and not(DecToCtl_port_sig.instrType = add) and not(DecToCtl_port_sig.instrType = sub) and not(DecToCtl_port_sig.instrType = sll_Instr) and not(DecToCtl_port_sig.instrType = slt) and not(DecToCtl_port_sig.instrType = sltu) and not(DecToCtl_port_sig.instrType = Xor_Instr) and not(DecToCtl_port_sig.instrType = srl_Instr) and not(DecToCtl_port_sig.instrType = sra_Instr) and not(DecToCtl_port_sig.instrType = Or_Instr) and not(DecToCtl_port_sig.instrType = And_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_987;
			elsif ((DecToCtl_port_sig.encType = R) and (DecToCtl_port_sig.instrType = And_Instr) and MemToCtl_port_sync) then 
				active_operation <= op_fetch_5_read_988;
			end if;
		when st_memoryOperation_6 =>
			elsif (not(memoryAccess.req = ME_RD) and not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and CtlToMem_port_sync) then 
				active_operation <= op_memoryOperation_6_write_991;
			elsif (not(CtlToMem_port_sync)) then 
				active_operation <= op_wait_memoryOperation_6;
			elsif ((memoryAccess.req = ME_RD) and CtlToMem_port_sync) then 
				active_operation <= op_memoryOperation_6_write_993;
			end if;
		when st_memoryOperation_7 =>
			elsif ((wb_sel = WB_MEM) and not(wb_en and not(decodedInstr.rd_addr = x"00000000")) and MemToCtl_port_sync) then 
				active_operation <= op_memoryOperation_7_read_998;
			elsif (not(wb_sel = WB_ALU) and not(wb_sel = WB_MEM) and not(wb_sel = WB_PC4) and MemToCtl_port_sync) then 
				active_operation <= op_memoryOperation_7_read_999;
			elsif (not(MemToCtl_port_sync)) then 
				active_operation <= op_wait_memoryOperation_7;
			elsif ((wb_sel = WB_MEM) and wb_en and not(decodedInstr.rd_addr = x"00000000") and MemToCtl_port_sync) then 
				active_operation <= op_memoryOperation_7_read_1002;
			end if;
		when st_readRegisterFile_8 =>
			if ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1004;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1007;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SUB)) then 
				active_operation <= op_readRegisterFile_8_write_1013;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_ADD)) then 
				active_operation <= op_readRegisterFile_8_write_1014;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1020;
			elsif (not(CtlToALU_data.op1_sel = OP_REG) and not(CtlToALU_data.op1_sel = OP_IMM) and not(CtlToALU_data.op1_sel = OP_PC) and not(CtlToALU_data.op2_sel = OP_REG) and not(CtlToALU_data.op2_sel = OP_IMM) and not(CtlToALU_data.op2_sel = OP_PC) and (CtlToALU_data.alu_fun = ALU_X)) then 
				active_operation <= op_readRegisterFile_8_write_1031;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1032;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_AND)) then 
				active_operation <= op_readRegisterFile_8_write_1033;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1044;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_OR)) then 
				active_operation <= op_readRegisterFile_8_write_1045;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_XOR)) then 
				active_operation <= op_readRegisterFile_8_write_1060;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and not(RegsToCtl_port_sig.contents2 <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1075;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLT) and (RegsToCtl_port_sig.contents2 <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1076;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(RegsToCtl_port_sig.contents2 <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1090;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLTU) and (RegsToCtl_port_sig.contents2 <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1091;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1092;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and not(decodedInstr.imm <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1093;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLT) and (decodedInstr.imm <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1094;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1105;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and not(decodedInstr.imm <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1106;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLTU) and (decodedInstr.imm <= RegsToCtl_port_sig.contents1)) then 
				active_operation <= op_readRegisterFile_8_write_1107;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SLL)) then 
				active_operation <= op_readRegisterFile_8_write_1108;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1124;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRA)) then 
				active_operation <= op_readRegisterFile_8_write_1125;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_REG) and (CtlToALU_data.alu_fun = ALU_COPY1)) then 
				active_operation <= op_readRegisterFile_8_write_1147;
			elsif ((CtlToALU_data.op1_sel = OP_REG) and (CtlToALU_data.op2_sel = OP_IMM) and (CtlToALU_data.alu_fun = ALU_SRL)) then 
				active_operation <= op_readRegisterFile_8_write_1148;
			end if;
		when st_writeBack_10 =>
			if (true) then 
				active_operation <= op_writeBack_10_write_1216;
			end if;
		end case;
	end process;

	-- Main process
	process (clk, rst)
	begin
		if (rst = '1') then
			decodedInstr.rd_addr <= x"00000000";
			decodedInstr.imm <= x"00000000";
			CtlToMem_port_sig.req <= ME_RD;
			br_en <= false;
			decodedInstr.instrType <= And_Instr;
			memoryAccess.req <= ME_RD;
			active_state <= st_fetch_4;
			CtlToMem_port_sig.addrIn <= x"00000000";
			MemToCtl_port_notify <= false;
			CtlToRegs_data.dst_data <= x"00000000";
			wb_sel <= WB_ALU;
			CtlToRegs_data.src1 <= x"00000000";
			ALUtoCtl_data.ALU_result <= x"00000000";
			CtlToALU_data.op2_sel <= OP_IMM;
			CtlToRegs_port_notify <= false;
			CtlToMem_port_sig.mask <= MT_W;
			fromMemoryData.loadedData <= x"00000000";
			CtlToALU_data.alu_fun <= ALU_ADD;
			CtlToALU_data.op1_sel <= OP_IMM;
			mem_en <= false;
			pc_next <= x"00000000";
			pc_reg <= x"00000000";
			memoryAccess.dataIn <= x"00000000";
			memoryAccess.addrIn <= x"00000000";
			RegsToCtl_data.contents2 <= x"00000000";
			CtlToDec_port_notify <= false;
			RegsToCtl_data.contents1 <= x"00000000";
			wb_en <= false;
			CtlToMem_port_notify <= true;
			memoryAccess.mask <= MT_W;
			CtlToRegs_data.dst <= x"00000000";
			CtlToRegs_data.src2 <= x"00000000";
			CtlToMem_port_sig.dataIn <= x"00000000";
			reg_rd_en <= false;
		elsif (clk = '1' and clk'event) then
			case active_operation is
			when op_wait_fetch_4 =>
				active_state <= st_fetch_4;
				CtlToMem_port_sig.addrIn <= memoryAccess.addrIn;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_sig.dataIn <= memoryAccess.dataIn;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
			when op_fetch_4_write_97 =>
				active_state <= st_fetch_5;
				CtlToMem_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				MemToCtl_port_notify <= true;
			when op_wait_fetch_5 =>
				active_state <= st_fetch_5;
				CtlToMem_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				MemToCtl_port_notify <= true;
			when op_fetch_5_read_98 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_101 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_102 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_110 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_111 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_112 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + DecToCtl_port_sig.imm;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_118 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_126 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_131 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + DecToCtl_port_sig.imm;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_137 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_138 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_139 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + DecToCtl_port_sig.imm;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_145 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_151 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_152 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and DecToCtl_port_sig.imm;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_160 =>
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_163 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_168 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + DecToCtl_port_sig.imm;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_174 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_175 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_176 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + DecToCtl_port_sig.imm;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_182 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_183 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_198 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_199 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and DecToCtl_port_sig.imm;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_207 =>
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_210 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_215 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + DecToCtl_port_sig.imm;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_221 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_222 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_237 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_238 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_253 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_254 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and DecToCtl_port_sig.imm;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_262 =>
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_265 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_266 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_280 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_295 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_296 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_311 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_312 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_313 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_314 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_315 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_326 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_327 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_341 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_342 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_357 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
			when op_fetch_5_read_358 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_359 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_360 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
			when op_fetch_5_read_376 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_377 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_378 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_379 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_380 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_393 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_394 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_408 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
			when op_fetch_5_read_409 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_431 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
			when op_fetch_5_read_432 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_433 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_434 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
			when op_fetch_5_read_450 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + RegsToCtl_data.contents2;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_456 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_457 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_458 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_459 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_460 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_471 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_472 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_495 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
			when op_fetch_5_read_496 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_518 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 - RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_519 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 + DecToCtl_port_sig.imm;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_525 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
			when op_fetch_5_read_526 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_527 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_528 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
			when op_fetch_5_read_564 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				CtlToALU_data.op1_sel <= OP_X;
				CtlToALU_data.op2_sel <= OP_X;
				wb_sel <= WB_PC4;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				CtlToALU_data.alu_fun <= ALU_X;
				reg_rd_en <= false;
			when op_fetch_5_read_565 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_566 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_589 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and RegsToCtl_data.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_594 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + DecToCtl_port_sig.imm;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_600 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_601 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
			when op_fetch_5_read_602 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_657 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or RegsToCtl_data.contents2;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_658 =>
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 and DecToCtl_port_sig.imm;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_666 =>
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_669 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_670 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_694 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_714 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor RegsToCtl_data.contents2;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_715 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 or DecToCtl_port_sig.imm;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_755 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_762 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1 xor DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_794 =>
				CtlToALU_data.op1_sel <= OP_PC;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm + pc_reg;
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				CtlToALU_data.alu_fun <= ALU_ADD;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_795 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_796 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_811 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_818 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_819 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_820 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_821 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_822 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_837 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				reg_rd_en <= false;
			when op_fetch_5_read_838 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_839 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				ALUtoCtl_data.ALU_result <= x"00000000";
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_840 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
			when op_fetch_5_read_856 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(RegsToCtl_data.contents2 and to_unsigned(31, 32)));
				reg_rd_en <= false;
			when op_fetch_5_read_857 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_879 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_data.contents1;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_880 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_data.contents1, to_integer(DecToCtl_port_sig.imm and to_unsigned(31, 32)));
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_937 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_948 =>
				active_state <= st_executeALU_2;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_port_notify <= false;
				CtlToALU_data.op1_sel <= OP_IMM;
				mem_en <= false;
				ALUtoCtl_data.ALU_result <= DecToCtl_port_sig.imm;
				CtlToALU_data.alu_fun <= ALU_COPY1;
				CtlToALU_data.op2_sel <= OP_X;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				reg_rd_en <= false;
			when op_fetch_5_read_949 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_950 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_951 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_952 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_953 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_954 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToALU_data.alu_fun <= ALU_SLT;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_955 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				CtlToALU_data.op1_sel <= OP_X;
				CtlToALU_data.op2_sel <= OP_X;
				wb_sel <= WB_PC4;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				CtlToALU_data.alu_fun <= ALU_X;
			when op_fetch_5_read_956 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToALU_data.alu_fun <= ALU_SUB;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_957 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToALU_data.alu_fun <= ALU_SUB;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_958 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToALU_data.alu_fun <= ALU_SLTU;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_959 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_SLL;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_960 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToALU_data.alu_fun <= ALU_SUB;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_961 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_XOR;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_962 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				mem_en <= true;
				memoryAccess.mask <= MT_B;
				wb_sel <= WB_MEM;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				memoryAccess.req <= ME_RD;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_963 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToALU_data.alu_fun <= ALU_SLT;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_964 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToALU_data.alu_fun <= ALU_SLT;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_965 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_OR;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_966 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				mem_en <= true;
				wb_sel <= WB_MEM;
				memoryAccess.mask <= MT_H;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				memoryAccess.req <= ME_RD;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_967 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToALU_data.alu_fun <= ALU_SLTU;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_968 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToALU_data.alu_fun <= ALU_SLT;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_969 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_AND;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_970 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				mem_en <= true;
				wb_sel <= WB_MEM;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				memoryAccess.req <= ME_RD;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				memoryAccess.mask <= MT_W;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_971 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_XOR;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_972 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToALU_data.alu_fun <= ALU_SLTU;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_973 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_974 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				memoryAccess.req <= ME_WR;
				mem_en <= true;
				memoryAccess.mask <= MT_B;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_975 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_SLL;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_976 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				memoryAccess.mask <= MT_BU;
				mem_en <= true;
				wb_sel <= WB_MEM;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				memoryAccess.req <= ME_RD;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_977 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToALU_data.alu_fun <= ALU_SRL;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_978 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= true;
				wb_sel <= WB_X;
				CtlToALU_data.alu_fun <= ALU_SLTU;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_979 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				memoryAccess.req <= ME_WR;
				mem_en <= true;
				memoryAccess.mask <= MT_H;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_980 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				memoryAccess.req <= ME_WR;
				mem_en <= true;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_981 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToALU_data.alu_fun <= ALU_SRL;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_982 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				mem_en <= true;
				wb_sel <= WB_MEM;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				memoryAccess.req <= ME_RD;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
				memoryAccess.mask <= MT_HU;
			when op_fetch_5_read_983 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.alu_fun <= ALU_SRA;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_984 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				memoryAccess.req <= ME_WR;
				mem_en <= true;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				wb_sel <= WB_X;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				CtlToALU_data.alu_fun <= ALU_ADD;
				wb_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				memoryAccess.mask <= MT_W;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_985 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				CtlToALU_data.alu_fun <= ALU_SRA;
				CtlToALU_data.op2_sel <= OP_IMM;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_986 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_OR;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_987 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_fetch_5_read_988 =>
				CtlToRegs_data.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToALU_data.alu_fun <= ALU_AND;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				br_en <= false;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.req <= REG_RD;
				CtlToRegs_port_sig.src1 <= DecToCtl_port_sig.rs1_addr;
				CtlToRegs_port_sig.src2 <= DecToCtl_port_sig.rs2_addr;
				reg_rd_en <= true;
				CtlToALU_data.op1_sel <= OP_REG;
				CtlToALU_data.op2_sel <= OP_REG;
				wb_en <= true;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				wb_sel <= WB_ALU;
				CtlToDec_port_notify <= true;
				decodedInstr.instrType <= DecToCtl_port_sig.instrType;
				decodedInstr.imm <= DecToCtl_port_sig.imm;
				CtlToRegs_data.src2 <= DecToCtl_port_sig.rs2_addr;
				CtlToRegs_port_sig.dst <= CtlToRegs_data.dst;
				CtlToRegs_port_sig.dst_data <= CtlToRegs_data.dst_data;
				mem_en <= false;
				decodedInstr.rd_addr <= DecToCtl_port_sig.rd_addr;
				active_state <= st_readRegisterFile_8;
				CtlToDec_port_sig <= MemToCtl_port_sig.loadedData;
			when op_executeALU_2_read_0 =>
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				active_state <= st_executeALU_3;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1004 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1007 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 + RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1013 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 - RegsToCtl_port_sig.contents2;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1014 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 + decodedInstr.imm;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1020 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 and RegsToCtl_port_sig.contents2;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1031 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1032 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 or RegsToCtl_port_sig.contents2;
			when op_readRegisterFile_8_write_1033 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 and decodedInstr.imm;
			when op_readRegisterFile_8_write_1044 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 xor RegsToCtl_port_sig.contents2;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1045 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 or decodedInstr.imm;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1060 =>
				active_state <= st_executeALU_2;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1 xor decodedInstr.imm;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1075 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1076 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1090 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1091 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1092 =>
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_port_sig.contents1, to_integer(RegsToCtl_port_sig.contents2 and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1093 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1094 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1105 =>
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_port_sig.contents1, to_integer(RegsToCtl_port_sig.contents2 and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1106 =>
				ALUtoCtl_data.ALU_result <= x"00000001";
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1107 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				ALUtoCtl_data.ALU_result <= x"00000000";
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1108 =>
				ALUtoCtl_data.ALU_result <= shift_left(RegsToCtl_port_sig.contents1, to_integer(decodedInstr.imm and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1124 =>
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_port_sig.contents1, to_integer(RegsToCtl_port_sig.contents2 and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1125 =>
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_port_sig.contents1, to_integer(decodedInstr.imm and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1147 =>
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				ALUtoCtl_data.ALU_result <= RegsToCtl_port_sig.contents1;
				CtlToDec_port_notify <= false;
			when op_readRegisterFile_8_write_1148 =>
				ALUtoCtl_data.ALU_result <= shift_right(RegsToCtl_port_sig.contents1, to_integer(decodedInstr.imm and to_unsigned(31, 32)));
				active_state <= st_executeALU_2;
				RegsToCtl_data.contents1 <= RegsToCtl_port_sig.contents1;
				RegsToCtl_data.contents2 <= RegsToCtl_port_sig.contents2;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
			when op_executeALU_3_read_1 =>
				memoryAccess.addrIn <= x"00000004" + pc_reg;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				pc_reg <= x"00000004" + pc_reg;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= x"00000004" + pc_reg;
			when op_executeALU_3_read_4 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_5 =>
				memoryAccess.addrIn <= x"00000004" + pc_reg;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				pc_reg <= x"00000004" + pc_reg;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= x"00000004" + pc_reg;
			when op_executeALU_3_read_10 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_12 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_13 =>
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				memoryAccess.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				pc_reg <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_16 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_22 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_25 =>
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				memoryAccess.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				pc_reg <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_28 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_31 =>
				memoryAccess.addrIn <= x"00000004" + pc_reg;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				pc_reg <= x"00000004" + pc_reg;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= x"00000004" + pc_reg;
			when op_executeALU_3_read_34 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_40 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_42 =>
				pc_reg <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				memoryAccess.addrIn <= pc_reg + decodedInstr.imm;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				CtlToMem_port_sig.addrIn <= pc_reg + decodedInstr.imm;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_47 =>
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				memoryAccess.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.addrIn <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= x"00000000";
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				pc_reg <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_49 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				pc_next <= x"00000004" + pc_reg;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_50 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				pc_next <= pc_reg + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_53 =>
				memoryAccess.addrIn <= ALUtoCtl_data.ALU_result;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
				memoryAccess.dataIn <= RegsToCtl_data.contents2;
				CtlToMem_port_sig.addrIn <= ALUtoCtl_data.ALU_result;
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
				CtlToMem_port_sig.dataIn <= RegsToCtl_data.contents2;
			when op_executeALU_3_read_61 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= x"00000004" + pc_reg;
			when op_executeALU_3_read_63 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_64 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= x"00000004" + pc_reg;
			when op_executeALU_3_read_69 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= pc_reg + decodedInstr.imm;
			when op_executeALU_3_read_70 =>
				CtlToRegs_data.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= ALUtoCtl_data.ALU_result;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_executeALU_3_read_79 =>
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.dst_data <= x"00000004" + pc_reg;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				CtlToRegs_data.dst_data <= x"00000004" + pc_reg;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
				pc_next <= RegsToCtl_data.contents1 + decodedInstr.imm;
			when op_memoryOperation_6_write_991 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_wait_memoryOperation_6 =>
				CtlToMem_port_sig.addrIn <= memoryAccess.addrIn;
				MemToCtl_port_notify <= false;
				active_state <= st_memoryOperation_6;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				CtlToMem_port_sig.dataIn <= memoryAccess.dataIn;
				CtlToMem_port_notify <= true;
				CtlToMem_port_sig.mask <= memoryAccess.mask;
				CtlToMem_port_sig.req <= memoryAccess.req;
			when op_memoryOperation_6_write_993 =>
				CtlToMem_port_notify <= false;
				active_state <= st_memoryOperation_7;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				MemToCtl_port_notify <= true;
			when op_writeBack_10_write_1216 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_memoryOperation_7_read_998 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_memoryOperation_7_read_999 =>
				memoryAccess.addrIn <= pc_next;
				CtlToMem_port_sig.req <= ME_RD;
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				memoryAccess.req <= ME_RD;
				active_state <= st_fetch_4;
				MemToCtl_port_notify <= false;
				pc_reg <= pc_next;
				CtlToRegs_port_notify <= false;
				CtlToMem_port_sig.mask <= MT_W;
				memoryAccess.dataIn <= x"00000000";
				CtlToMem_port_sig.addrIn <= pc_next;
				CtlToDec_port_notify <= false;
				CtlToMem_port_notify <= true;
				memoryAccess.mask <= MT_W;
				CtlToMem_port_sig.dataIn <= x"00000000";
			when op_wait_memoryOperation_7 =>
				CtlToMem_port_notify <= false;
				active_state <= st_memoryOperation_7;
				CtlToRegs_port_notify <= false;
				CtlToDec_port_notify <= false;
				MemToCtl_port_notify <= true;
			when op_memoryOperation_7_read_1002 =>
				fromMemoryData.loadedData <= MemToCtl_port_sig.loadedData;
				CtlToRegs_data.dst_data <= MemToCtl_port_sig.loadedData;
				CtlToRegs_port_sig.dst_data <= MemToCtl_port_sig.loadedData;
				CtlToRegs_port_notify <= true;
				CtlToRegs_port_sig.src1 <= CtlToRegs_data.src1;
				CtlToMem_port_notify <= false;
				MemToCtl_port_notify <= false;
				CtlToRegs_port_sig.req <= REG_WR;
				CtlToRegs_port_sig.src2 <= CtlToRegs_data.src2;
				active_state <= st_writeBack_10;
				CtlToDec_port_notify <= false;
				CtlToRegs_port_sig.dst <= decodedInstr.rd_addr;
				CtlToRegs_data.dst <= decodedInstr.rd_addr;
			end case;
		end if;
	end process;

	-- Assigning state signals that are used by ITL properties for OneSpin
	executeALU_2 <= active_state = st_executeALU_2;
	executeALU_3 <= active_state = st_executeALU_3;
	fetch_4 <= active_state = st_fetch_4;
	fetch_5 <= active_state = st_fetch_5;
	memoryOperation_6 <= active_state = st_memoryOperation_6;
	memoryOperation_7 <= active_state = st_memoryOperation_7;
	readRegisterFile_8 <= active_state = st_readRegisterFile_8;
	writeBack_10 <= active_state = st_writeBack_10;

end ISA_arch;

