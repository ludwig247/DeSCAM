package testbasic18_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic18_SECTIONS;

endpackage
