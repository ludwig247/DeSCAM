library ieee;
use IEEE.numeric_std.all;
use work.SCAM_Model_types.all;

package TestArray0_types is
end package TestArray0_types;