library ieee;
use IEEE.numeric_std.all;

package TestBasic8_types is
type TestBasic8_SECTIONS is (run);
end package TestBasic8_types;
