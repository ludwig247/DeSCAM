library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.SCAM_Model_types.all;

entity Regs is
port(	
	ISAtoRF_port_sig: in RegfileWriteType;
	ISAtoRF_port_sync: in boolean;
	RFtoISA_port_sig: out RegfileType;
	clk: in std_logic;
	rst: in std_logic
);
end Regs;

architecture Regs_arch of Regs is
	-- Define internal data types
	type Regs_operation_t is (op_run_0_write_0, op_run_0_write_1, op_run_0_write_2, op_run_0_write_3, op_run_0_write_4, op_run_0_write_5, op_run_0_write_6, op_run_0_write_7, op_run_0_write_8, op_run_0_write_9, op_run_0_write_10, op_run_0_write_11, op_run_0_write_12, op_run_0_write_13, op_run_0_write_14, op_run_0_write_15, op_run_0_write_16, op_run_0_write_17, op_run_0_write_18, op_run_0_write_19, op_run_0_write_20, op_run_0_write_21, op_run_0_write_22, op_run_0_write_23, op_run_0_write_24, op_run_0_write_25, op_run_0_write_26, op_run_0_write_27, op_run_0_write_28, op_run_0_write_29, op_run_0_write_30, op_run_0_write_31, op_run_0_write_32);
	type Regs_state_t is (st_run_0);

	-- Declare signals
	signal active_state: Regs_state_t;
	signal active_operation: Regs_operation_t;
	signal reg_file_01: unsigned(31 downto 0);
	signal reg_file_02: unsigned(31 downto 0);
	signal reg_file_03: unsigned(31 downto 0);
	signal reg_file_04: unsigned(31 downto 0);
	signal reg_file_05: unsigned(31 downto 0);
	signal reg_file_06: unsigned(31 downto 0);
	signal reg_file_07: unsigned(31 downto 0);
	signal reg_file_08: unsigned(31 downto 0);
	signal reg_file_09: unsigned(31 downto 0);
	signal reg_file_10: unsigned(31 downto 0);
	signal reg_file_11: unsigned(31 downto 0);
	signal reg_file_12: unsigned(31 downto 0);
	signal reg_file_13: unsigned(31 downto 0);
	signal reg_file_14: unsigned(31 downto 0);
	signal reg_file_15: unsigned(31 downto 0);
	signal reg_file_16: unsigned(31 downto 0);
	signal reg_file_17: unsigned(31 downto 0);
	signal reg_file_18: unsigned(31 downto 0);
	signal reg_file_19: unsigned(31 downto 0);
	signal reg_file_20: unsigned(31 downto 0);
	signal reg_file_21: unsigned(31 downto 0);
	signal reg_file_22: unsigned(31 downto 0);
	signal reg_file_23: unsigned(31 downto 0);
	signal reg_file_24: unsigned(31 downto 0);
	signal reg_file_25: unsigned(31 downto 0);
	signal reg_file_26: unsigned(31 downto 0);
	signal reg_file_27: unsigned(31 downto 0);
	signal reg_file_28: unsigned(31 downto 0);
	signal reg_file_29: unsigned(31 downto 0);
	signal reg_file_30: unsigned(31 downto 0);
	signal reg_file_31: unsigned(31 downto 0);

	-- Declare state signals that are used by ITL properties for OneSpin
	signal run_0: boolean;


begin
	-- Combinational logic that selects current operation
	process (active_state, ISAtoRF_port_sync, ISAtoRF_port_sig.dst)
	begin
		case active_state is
		when st_run_0 =>
			if (not(ISAtoRF_port_sync)) then 
				active_operation <= op_run_0_write_0;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000000") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_1;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000001") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_2;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000002") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_3;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000003") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_4;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000004") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_5;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000005") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_6;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000006") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_7;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000007") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_8;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000008") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_9;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000009") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_10;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000000a") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_11;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000000b") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_12;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000000c") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_13;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000000d") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_14;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000000e") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_15;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000000f") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_16;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000010") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_17;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000011") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_18;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000012") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_19;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000013") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_20;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000014") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_21;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000015") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_22;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000016") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_23;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000017") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_24;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000018") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_25;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000019") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_26;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000001a") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_27;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000001b") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_28;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000001c") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_29;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000001d") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_30;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000001e") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_31;
			else--if(ISAtoRF_port_sync and not(ISAtoRF_port_sig.dst = x"00000000") and not(ISAtoRF_port_sig.dst = x"00000001") and not(ISAtoRF_port_sig.dst = x"00000002") and not(ISAtoRF_port_sig.dst = x"00000003") and not(ISAtoRF_port_sig.dst = x"00000004") and not(ISAtoRF_port_sig.dst = x"00000005") and not(ISAtoRF_port_sig.dst = x"00000006") and not(ISAtoRF_port_sig.dst = x"00000007") and not(ISAtoRF_port_sig.dst = x"00000008") and not(ISAtoRF_port_sig.dst = x"00000009") and not(ISAtoRF_port_sig.dst = x"0000000a") and not(ISAtoRF_port_sig.dst = x"0000000b") and not(ISAtoRF_port_sig.dst = x"0000000c") and not(ISAtoRF_port_sig.dst = x"0000000d") and not(ISAtoRF_port_sig.dst = x"0000000e") and not(ISAtoRF_port_sig.dst = x"0000000f") and not(ISAtoRF_port_sig.dst = x"00000010") and not(ISAtoRF_port_sig.dst = x"00000011") and not(ISAtoRF_port_sig.dst = x"00000012") and not(ISAtoRF_port_sig.dst = x"00000013") and not(ISAtoRF_port_sig.dst = x"00000014") and not(ISAtoRF_port_sig.dst = x"00000015") and not(ISAtoRF_port_sig.dst = x"00000016") and not(ISAtoRF_port_sig.dst = x"00000017") and not(ISAtoRF_port_sig.dst = x"00000018") and not(ISAtoRF_port_sig.dst = x"00000019") and not(ISAtoRF_port_sig.dst = x"0000001a") and not(ISAtoRF_port_sig.dst = x"0000001b") and not(ISAtoRF_port_sig.dst = x"0000001c") and not(ISAtoRF_port_sig.dst = x"0000001d") and not(ISAtoRF_port_sig.dst = x"0000001e") and ISAtoRF_port_sync) then 
				active_operation <= op_run_0_write_32;
			end if;
		end case;
	end process;

	-- Main process
	process (clk, rst)
	begin
		if (rst = '1') then
			RFtoISA_port_sig.reg_file_20 <= x"00000000";
			RFtoISA_port_sig.reg_file_18 <= x"00000000";
			RFtoISA_port_sig.reg_file_09 <= x"00000000";
			reg_file_28 <= x"00000000";
			RFtoISA_port_sig.reg_file_13 <= x"00000000";
			RFtoISA_port_sig.reg_file_23 <= x"00000000";
			RFtoISA_port_sig.reg_file_04 <= x"00000000";
			reg_file_11 <= x"00000000";
			reg_file_12 <= x"00000000";
			reg_file_13 <= x"00000000";
			reg_file_14 <= x"00000000";
			RFtoISA_port_sig.reg_file_30 <= x"00000000";
			RFtoISA_port_sig.reg_file_31 <= x"00000000";
			reg_file_04 <= x"00000000";
			reg_file_05 <= x"00000000";
			reg_file_06 <= x"00000000";
			RFtoISA_port_sig.reg_file_22 <= x"00000000";
			reg_file_01 <= x"00000000";
			reg_file_02 <= x"00000000";
			RFtoISA_port_sig.reg_file_19 <= x"00000000";
			reg_file_03 <= x"00000000";
			RFtoISA_port_sig.reg_file_12 <= x"00000000";
			RFtoISA_port_sig.reg_file_01 <= x"00000000";
			RFtoISA_port_sig.reg_file_03 <= x"00000000";
			RFtoISA_port_sig.reg_file_06 <= x"00000000";
			reg_file_22 <= x"00000000";
			reg_file_15 <= x"00000000";
			reg_file_16 <= x"00000000";
			reg_file_31 <= x"00000000";
			reg_file_21 <= x"00000000";
			reg_file_17 <= x"00000000";
			RFtoISA_port_sig.reg_file_24 <= x"00000000";
			RFtoISA_port_sig.reg_file_05 <= x"00000000";
			reg_file_18 <= x"00000000";
			reg_file_19 <= x"00000000";
			reg_file_20 <= x"00000000";
			reg_file_26 <= x"00000000";
			reg_file_27 <= x"00000000";
			reg_file_07 <= x"00000000";
			reg_file_08 <= x"00000000";
			reg_file_09 <= x"00000000";
			reg_file_10 <= x"00000000";
			reg_file_23 <= x"00000000";
			RFtoISA_port_sig.reg_file_17 <= x"00000000";
			RFtoISA_port_sig.reg_file_07 <= x"00000000";
			reg_file_29 <= x"00000000";
			reg_file_30 <= x"00000000";
			RFtoISA_port_sig.reg_file_26 <= x"00000000";
			RFtoISA_port_sig.reg_file_27 <= x"00000000";
			RFtoISA_port_sig.reg_file_08 <= x"00000000";
			RFtoISA_port_sig.reg_file_28 <= x"00000000";
			RFtoISA_port_sig.reg_file_29 <= x"00000000";
			reg_file_25 <= x"00000000";
			active_state <= st_run_0;
			RFtoISA_port_sig.reg_file_14 <= x"00000000";
			RFtoISA_port_sig.reg_file_15 <= x"00000000";
			RFtoISA_port_sig.reg_file_16 <= x"00000000";
			RFtoISA_port_sig.reg_file_25 <= x"00000000";
			RFtoISA_port_sig.reg_file_02 <= x"00000000";
			RFtoISA_port_sig.reg_file_10 <= x"00000000";
			reg_file_24 <= x"00000000";
			RFtoISA_port_sig.reg_file_11 <= x"00000000";
			RFtoISA_port_sig.reg_file_21 <= x"00000000";
		elsif (clk = '1' and clk'event) then
			case active_operation is
			when op_run_0_write_0 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_1 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_2 =>
				RFtoISA_port_sig.reg_file_01 <= ISAtoRF_port_sig.dstData;
				reg_file_01 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_3 =>
				RFtoISA_port_sig.reg_file_02 <= ISAtoRF_port_sig.dstData;
				reg_file_02 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_4 =>
				reg_file_03 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_03 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_5 =>
				RFtoISA_port_sig.reg_file_04 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				reg_file_04 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_6 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_05 <= ISAtoRF_port_sig.dstData;
				reg_file_05 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_7 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				reg_file_06 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_06 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_8 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_07 <= ISAtoRF_port_sig.dstData;
				reg_file_07 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_9 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_08 <= ISAtoRF_port_sig.dstData;
				reg_file_08 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_10 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_09 <= ISAtoRF_port_sig.dstData;
				reg_file_09 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_11 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_10 <= ISAtoRF_port_sig.dstData;
				reg_file_10 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_12 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				reg_file_11 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_11 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_13 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_12 <= ISAtoRF_port_sig.dstData;
				reg_file_12 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_14 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_13 <= ISAtoRF_port_sig.dstData;
				reg_file_13 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_15 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				reg_file_14 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_14 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_16 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_15 <= ISAtoRF_port_sig.dstData;
				reg_file_15 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_17 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_16 <= ISAtoRF_port_sig.dstData;
				reg_file_16 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_18 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_17 <= ISAtoRF_port_sig.dstData;
				reg_file_17 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_19 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_18 <= ISAtoRF_port_sig.dstData;
				reg_file_18 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_20 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_19 <= ISAtoRF_port_sig.dstData;
				reg_file_19 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_21 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_20 <= ISAtoRF_port_sig.dstData;
				reg_file_20 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_22 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				reg_file_21 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_21 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_23 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_22 <= ISAtoRF_port_sig.dstData;
				reg_file_22 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_24 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_23 <= ISAtoRF_port_sig.dstData;
				reg_file_23 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_25 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_24 <= ISAtoRF_port_sig.dstData;
				reg_file_24 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_26 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_25 <= ISAtoRF_port_sig.dstData;
				reg_file_25 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_27 =>
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				reg_file_26 <= ISAtoRF_port_sig.dstData;
				active_state <= st_run_0;
				RFtoISA_port_sig.reg_file_26 <= ISAtoRF_port_sig.dstData;
			when op_run_0_write_28 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				RFtoISA_port_sig.reg_file_27 <= ISAtoRF_port_sig.dstData;
				reg_file_27 <= ISAtoRF_port_sig.dstData;
				active_state <= st_run_0;
			when op_run_0_write_29 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				RFtoISA_port_sig.reg_file_28 <= ISAtoRF_port_sig.dstData;
				reg_file_28 <= ISAtoRF_port_sig.dstData;
				active_state <= st_run_0;
			when op_run_0_write_30 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				reg_file_29 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				RFtoISA_port_sig.reg_file_29 <= ISAtoRF_port_sig.dstData;
				active_state <= st_run_0;
			when op_run_0_write_31 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_31 <= reg_file_31;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_30 <= ISAtoRF_port_sig.dstData;
				reg_file_30 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			when op_run_0_write_32 =>
				RFtoISA_port_sig.reg_file_26 <= reg_file_26;
				RFtoISA_port_sig.reg_file_27 <= reg_file_27;
				RFtoISA_port_sig.reg_file_28 <= reg_file_28;
				RFtoISA_port_sig.reg_file_29 <= reg_file_29;
				RFtoISA_port_sig.reg_file_30 <= reg_file_30;
				RFtoISA_port_sig.reg_file_22 <= reg_file_22;
				RFtoISA_port_sig.reg_file_23 <= reg_file_23;
				RFtoISA_port_sig.reg_file_24 <= reg_file_24;
				RFtoISA_port_sig.reg_file_25 <= reg_file_25;
				RFtoISA_port_sig.reg_file_10 <= reg_file_10;
				RFtoISA_port_sig.reg_file_11 <= reg_file_11;
				RFtoISA_port_sig.reg_file_12 <= reg_file_12;
				RFtoISA_port_sig.reg_file_13 <= reg_file_13;
				RFtoISA_port_sig.reg_file_14 <= reg_file_14;
				RFtoISA_port_sig.reg_file_15 <= reg_file_15;
				RFtoISA_port_sig.reg_file_16 <= reg_file_16;
				RFtoISA_port_sig.reg_file_17 <= reg_file_17;
				RFtoISA_port_sig.reg_file_18 <= reg_file_18;
				RFtoISA_port_sig.reg_file_19 <= reg_file_19;
				RFtoISA_port_sig.reg_file_20 <= reg_file_20;
				RFtoISA_port_sig.reg_file_21 <= reg_file_21;
				RFtoISA_port_sig.reg_file_31 <= ISAtoRF_port_sig.dstData;
				reg_file_31 <= ISAtoRF_port_sig.dstData;
				RFtoISA_port_sig.reg_file_01 <= reg_file_01;
				RFtoISA_port_sig.reg_file_03 <= reg_file_03;
				RFtoISA_port_sig.reg_file_02 <= reg_file_02;
				RFtoISA_port_sig.reg_file_04 <= reg_file_04;
				RFtoISA_port_sig.reg_file_05 <= reg_file_05;
				RFtoISA_port_sig.reg_file_06 <= reg_file_06;
				RFtoISA_port_sig.reg_file_07 <= reg_file_07;
				RFtoISA_port_sig.reg_file_08 <= reg_file_08;
				RFtoISA_port_sig.reg_file_09 <= reg_file_09;
				active_state <= st_run_0;
			end case;
		end if;
	end process;

	-- Assigning state signals that are used by ITL properties for OneSpin
	run_0 <= active_state = st_run_0;

end Regs_arch;

