package testmasterslave6_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave6_SECTIONS;

endpackage
