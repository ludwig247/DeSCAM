package testbasic7_types;

	import scam_model_types::*;
endpackage