library ieee;
use IEEE.numeric_std.all;

package SCAM_Model_types is
type states is (Aw,A,Bw,B);
end package SCAM_Model_types;