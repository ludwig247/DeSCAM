package testarray5_types;

	import scam_model_types::*;
endpackage