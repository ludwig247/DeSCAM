library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave9_types is
type TestMasterSlave9_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave9_types;

