package testfunction0_types;

	import scam_model_types::*;
endpackage