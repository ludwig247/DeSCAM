package testarray3_types;

	 import top_level_types::*;
endpackage