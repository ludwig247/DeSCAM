package testbasic12_types;

	import top_level_types::*;
	typedef enum logic {
		section_a,
		section_b
	} Phases;

endpackage