library ieee;
use IEEE.numeric_std.all;

package TestBasic3_types is
type TestBasic3_SECTIONS is (run);
end package TestBasic3_types;
