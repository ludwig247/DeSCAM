package testbasic3_types;

endpackage