
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_CPU is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type UNSIGNED is array (INTEGER range <>) of std_logic;

end CONV_PACK_CPU;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_53 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_53;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_52 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_52;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_51 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_51;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_50 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_50;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_49 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_49;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_48 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_48;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_47 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_47;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_46 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_46;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_45 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_45;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_44 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_44;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_43 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_43;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_42 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_42;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_41 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_41;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_40 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_40;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_39 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_39;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_38 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_38;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_37 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_37;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_34 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_34;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_33 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_33;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_32 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_32;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_31 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_31;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_30 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_30;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_29 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_29;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_28 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_28;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_27 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_27;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_26 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_26;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_25 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_25;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_24 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_24;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_23 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_23;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_22 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_22;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_21 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_21;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_20 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_20;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_19 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_19;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_18 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_18;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_17 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_17;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_16 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_16;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_15 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_15;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_14 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_14;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_13 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_13;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_12 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_12;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_11 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_11;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_10 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_10;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_9 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_9;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_8 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_8;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_7 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_7;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_6 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_6;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_5 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_5;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_4 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_4;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_3 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_3;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_2 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_2;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_1 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_1;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_36 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_36;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_54 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_54;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_0;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net2468138 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net2468138);
   main_gate : AND2_X1 port map( A1 => net2468138, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity CPU is

   port( clk, rst : in std_logic;  MemToCtl_port : in UNSIGNED (31 downto 0);  
         MemToCtl_port_sync : in std_logic;  MemToCtl_port_notify : out 
         std_logic;  CtlToMem_port_addrIn, CtlToMem_port_dataIn : out UNSIGNED 
         (31 downto 0);  CtlToMem_port_mask : out UNSIGNED (2 downto 0);  
         CtlToMem_port_req : out std_logic;  CtlToMem_port_sync : in std_logic;
         CtlToMem_port_notify : out std_logic);

end CPU;

architecture SYN_CPU_arch of CPU is

   component SNPS_CLOCK_GATE_HIGH_CPU_1
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_2
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_3
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_4
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_5
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_6
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_7
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_8
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_9
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_10
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_11
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_12
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_13
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_14
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_15
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_16
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_17
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_18
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_19
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_20
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_21
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_22
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_23
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_24
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_25
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_26
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_27
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_28
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_29
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_30
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_31
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_32
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_33
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_34
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_36
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_37
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_38
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_39
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_40
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_41
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_42
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_43
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_44
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_45
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_46
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_47
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_48
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_49
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_50
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_51
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_52
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_53
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_54
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal MemToCtl_port_notify_port, CtlToMem_port_notify_port, 
      ALUtoCtl_port_31_port, ALUtoCtl_port_30_port, ALUtoCtl_port_29_port, 
      ALUtoCtl_port_28_port, ALUtoCtl_port_27_port, ALUtoCtl_port_26_port, 
      ALUtoCtl_port_25_port, ALUtoCtl_port_24_port, ALUtoCtl_port_23_port, 
      ALUtoCtl_port_22_port, ALUtoCtl_port_21_port, ALUtoCtl_port_20_port, 
      ALUtoCtl_port_19_port, ALUtoCtl_port_18_port, ALUtoCtl_port_17_port, 
      ALUtoCtl_port_16_port, ALUtoCtl_port_15_port, ALUtoCtl_port_14_port, 
      ALUtoCtl_port_13_port, ALUtoCtl_port_12_port, ALUtoCtl_port_11_port, 
      ALUtoCtl_port_10_port, ALUtoCtl_port_9_port, ALUtoCtl_port_8_port, 
      ALUtoCtl_port_7_port, ALUtoCtl_port_6_port, ALUtoCtl_port_5_port, 
      ALUtoCtl_port_4_port, ALUtoCtl_port_3_port, ALUtoCtl_port_2_port, 
      ALUtoCtl_port_1_port, ALUtoCtl_port_0_port, CtlToALU_port_alu_fun_3_port,
      CtlToALU_port_alu_fun_2_port, CtlToALU_port_alu_fun_1_port, 
      CtlToALU_port_alu_fun_0_port, CtlToALU_port_imm_31_port, 
      CtlToALU_port_imm_30_port, CtlToALU_port_imm_29_port, 
      CtlToALU_port_imm_28_port, CtlToALU_port_imm_27_port, 
      CtlToALU_port_imm_26_port, CtlToALU_port_imm_25_port, 
      CtlToALU_port_imm_24_port, CtlToALU_port_imm_23_port, 
      CtlToALU_port_imm_22_port, CtlToALU_port_imm_21_port, 
      CtlToALU_port_imm_20_port, CtlToALU_port_imm_19_port, 
      CtlToALU_port_imm_18_port, CtlToALU_port_imm_17_port, 
      CtlToALU_port_imm_16_port, CtlToALU_port_imm_15_port, 
      CtlToALU_port_imm_14_port, CtlToALU_port_imm_13_port, 
      CtlToALU_port_imm_12_port, CtlToALU_port_imm_11_port, 
      CtlToALU_port_imm_10_port, CtlToALU_port_imm_9_port, 
      CtlToALU_port_imm_8_port, CtlToALU_port_imm_7_port, 
      CtlToALU_port_imm_6_port, CtlToALU_port_imm_5_port, 
      CtlToALU_port_imm_4_port, CtlToALU_port_imm_3_port, 
      CtlToALU_port_imm_2_port, CtlToALU_port_imm_1_port, 
      CtlToALU_port_imm_0_port, CtlToALU_port_op1_sel_1_port, 
      CtlToALU_port_op1_sel_0_port, CtlToALU_port_op2_sel_1_port, 
      CtlToALU_port_op2_sel_0_port, CtlToALU_port_pc_reg_31_port, 
      CtlToALU_port_pc_reg_30_port, CtlToALU_port_pc_reg_29_port, 
      CtlToALU_port_pc_reg_28_port, CtlToALU_port_pc_reg_27_port, 
      CtlToALU_port_pc_reg_26_port, CtlToALU_port_pc_reg_25_port, 
      CtlToALU_port_pc_reg_24_port, CtlToALU_port_pc_reg_23_port, 
      CtlToALU_port_pc_reg_22_port, CtlToALU_port_pc_reg_21_port, 
      CtlToALU_port_pc_reg_20_port, CtlToALU_port_pc_reg_19_port, 
      CtlToALU_port_pc_reg_18_port, CtlToALU_port_pc_reg_17_port, 
      CtlToALU_port_pc_reg_16_port, CtlToALU_port_pc_reg_15_port, 
      CtlToALU_port_pc_reg_14_port, CtlToALU_port_pc_reg_13_port, 
      CtlToALU_port_pc_reg_12_port, CtlToALU_port_pc_reg_11_port, 
      CtlToALU_port_pc_reg_10_port, CtlToALU_port_pc_reg_9_port, 
      CtlToALU_port_pc_reg_8_port, CtlToALU_port_pc_reg_7_port, 
      CtlToALU_port_pc_reg_6_port, CtlToALU_port_pc_reg_5_port, 
      CtlToALU_port_pc_reg_4_port, CtlToALU_port_pc_reg_3_port, 
      CtlToALU_port_pc_reg_2_port, CtlToALU_port_pc_reg_1_port, 
      CtlToALU_port_pc_reg_0_port, CtlToALU_port_reg1_contents_31_port, 
      CtlToALU_port_reg1_contents_30_port, CtlToALU_port_reg1_contents_29_port,
      CtlToALU_port_reg1_contents_28_port, CtlToALU_port_reg1_contents_27_port,
      CtlToALU_port_reg1_contents_26_port, CtlToALU_port_reg1_contents_25_port,
      CtlToALU_port_reg1_contents_24_port, CtlToALU_port_reg1_contents_23_port,
      CtlToALU_port_reg1_contents_22_port, CtlToALU_port_reg1_contents_21_port,
      CtlToALU_port_reg1_contents_20_port, CtlToALU_port_reg1_contents_19_port,
      CtlToALU_port_reg1_contents_18_port, CtlToALU_port_reg1_contents_17_port,
      CtlToALU_port_reg1_contents_16_port, CtlToALU_port_reg1_contents_15_port,
      CtlToALU_port_reg1_contents_14_port, CtlToALU_port_reg1_contents_13_port,
      CtlToALU_port_reg1_contents_12_port, CtlToALU_port_reg1_contents_11_port,
      CtlToALU_port_reg1_contents_10_port, CtlToALU_port_reg1_contents_9_port, 
      CtlToALU_port_reg1_contents_8_port, CtlToALU_port_reg1_contents_7_port, 
      CtlToALU_port_reg1_contents_6_port, CtlToALU_port_reg1_contents_5_port, 
      CtlToALU_port_reg1_contents_4_port, CtlToALU_port_reg1_contents_3_port, 
      CtlToALU_port_reg1_contents_2_port, CtlToALU_port_reg1_contents_1_port, 
      CtlToALU_port_reg1_contents_0_port, CtlToALU_port_reg2_contents_31_port, 
      CtlToALU_port_reg2_contents_30_port, CtlToALU_port_reg2_contents_29_port,
      CtlToALU_port_reg2_contents_28_port, CtlToALU_port_reg2_contents_27_port,
      CtlToALU_port_reg2_contents_26_port, CtlToALU_port_reg2_contents_25_port,
      CtlToALU_port_reg2_contents_24_port, CtlToALU_port_reg2_contents_23_port,
      CtlToALU_port_reg2_contents_22_port, CtlToALU_port_reg2_contents_21_port,
      CtlToALU_port_reg2_contents_20_port, CtlToALU_port_reg2_contents_19_port,
      CtlToALU_port_reg2_contents_18_port, CtlToALU_port_reg2_contents_17_port,
      CtlToALU_port_reg2_contents_16_port, CtlToALU_port_reg2_contents_15_port,
      CtlToALU_port_reg2_contents_14_port, CtlToALU_port_reg2_contents_13_port,
      CtlToALU_port_reg2_contents_12_port, CtlToALU_port_reg2_contents_11_port,
      CtlToALU_port_reg2_contents_10_port, CtlToALU_port_reg2_contents_9_port, 
      CtlToALU_port_reg2_contents_8_port, CtlToALU_port_reg2_contents_7_port, 
      CtlToALU_port_reg2_contents_6_port, CtlToALU_port_reg2_contents_5_port, 
      CtlToALU_port_reg2_contents_4_port, CtlToALU_port_reg2_contents_3_port, 
      CtlToALU_port_reg2_contents_2_port, CtlToALU_port_reg2_contents_1_port, 
      CtlToALU_port_reg2_contents_0_port, CtlToALU_port_notify, 
      CtlToRegs_port_dst_4_port, CtlToRegs_port_dst_3_port, 
      CtlToRegs_port_dst_2_port, CtlToRegs_port_dst_1_port, 
      CtlToRegs_port_dst_0_port, CtlToRegs_port_dst_data_31_port, 
      CtlToRegs_port_dst_data_30_port, CtlToRegs_port_dst_data_29_port, 
      CtlToRegs_port_dst_data_28_port, CtlToRegs_port_dst_data_27_port, 
      CtlToRegs_port_dst_data_26_port, CtlToRegs_port_dst_data_25_port, 
      CtlToRegs_port_dst_data_24_port, CtlToRegs_port_dst_data_23_port, 
      CtlToRegs_port_dst_data_22_port, CtlToRegs_port_dst_data_21_port, 
      CtlToRegs_port_dst_data_20_port, CtlToRegs_port_dst_data_19_port, 
      CtlToRegs_port_dst_data_18_port, CtlToRegs_port_dst_data_17_port, 
      CtlToRegs_port_dst_data_16_port, CtlToRegs_port_dst_data_15_port, 
      CtlToRegs_port_dst_data_14_port, CtlToRegs_port_dst_data_13_port, 
      CtlToRegs_port_dst_data_12_port, CtlToRegs_port_dst_data_11_port, 
      CtlToRegs_port_dst_data_10_port, CtlToRegs_port_dst_data_9_port, 
      CtlToRegs_port_dst_data_8_port, CtlToRegs_port_dst_data_7_port, 
      CtlToRegs_port_dst_data_6_port, CtlToRegs_port_dst_data_5_port, 
      CtlToRegs_port_dst_data_4_port, CtlToRegs_port_dst_data_3_port, 
      CtlToRegs_port_dst_data_2_port, CtlToRegs_port_dst_data_1_port, 
      CtlToRegs_port_dst_data_0_port, CtlToRegs_port_req, 
      CtlToRegs_port_src1_4_port, CtlToRegs_port_src1_3_port, 
      CtlToRegs_port_src1_2_port, CtlToRegs_port_src1_1_port, 
      CtlToRegs_port_src1_0_port, CtlToRegs_port_src2_4_port, 
      CtlToRegs_port_src2_3_port, CtlToRegs_port_src2_2_port, 
      CtlToRegs_port_src2_0_port, CtlToRegs_port_notify, 
      RegsToCtl_port_contents1_31_port, RegsToCtl_port_contents1_30_port, 
      RegsToCtl_port_contents1_29_port, RegsToCtl_port_contents1_28_port, 
      RegsToCtl_port_contents1_27_port, RegsToCtl_port_contents1_26_port, 
      RegsToCtl_port_contents1_25_port, RegsToCtl_port_contents1_24_port, 
      RegsToCtl_port_contents1_23_port, RegsToCtl_port_contents1_22_port, 
      RegsToCtl_port_contents1_21_port, RegsToCtl_port_contents1_20_port, 
      RegsToCtl_port_contents1_19_port, RegsToCtl_port_contents1_18_port, 
      RegsToCtl_port_contents1_17_port, RegsToCtl_port_contents1_16_port, 
      RegsToCtl_port_contents1_15_port, RegsToCtl_port_contents1_14_port, 
      RegsToCtl_port_contents1_13_port, RegsToCtl_port_contents1_12_port, 
      RegsToCtl_port_contents1_11_port, RegsToCtl_port_contents1_10_port, 
      RegsToCtl_port_contents1_9_port, RegsToCtl_port_contents1_8_port, 
      RegsToCtl_port_contents1_7_port, RegsToCtl_port_contents1_6_port, 
      RegsToCtl_port_contents1_5_port, RegsToCtl_port_contents2_31_port, 
      RegsToCtl_port_contents2_30_port, RegsToCtl_port_contents2_29_port, 
      RegsToCtl_port_contents2_28_port, RegsToCtl_port_contents2_27_port, 
      RegsToCtl_port_contents2_26_port, RegsToCtl_port_contents2_25_port, 
      RegsToCtl_port_contents2_24_port, RegsToCtl_port_contents2_23_port, 
      RegsToCtl_port_contents2_22_port, RegsToCtl_port_contents2_21_port, 
      RegsToCtl_port_contents2_20_port, RegsToCtl_port_contents2_19_port, 
      RegsToCtl_port_contents2_18_port, RegsToCtl_port_contents2_17_port, 
      RegsToCtl_port_contents2_16_port, RegsToCtl_port_contents2_15_port, 
      RegsToCtl_port_contents2_14_port, RegsToCtl_port_contents2_13_port, 
      RegsToCtl_port_contents2_12_port, RegsToCtl_port_contents2_11_port, 
      RegsToCtl_port_contents2_10_port, RegsToCtl_port_contents2_9_port, 
      RegsToCtl_port_contents2_8_port, RegsToCtl_port_contents2_7_port, 
      RegsToCtl_port_contents2_6_port, RegsToCtl_port_contents2_5_port, 
      RegsToCtl_port_contents2_4_port, RegsToCtl_port_contents2_3_port, 
      RegsToCtl_port_contents2_2_port, RegsToCtl_port_contents2_1_port, 
      RegsToCtl_port_contents2_0_port, CtlToDec_port_31_port, 
      CtlToDec_port_30_port, CtlToDec_port_29_port, CtlToDec_port_28_port, 
      CtlToDec_port_27_port, CtlToDec_port_26_port, CtlToDec_port_20_port, 
      CtlToDec_port_14_port, CtlToDec_port_13_port, CtlToDec_port_12_port, 
      CtlToDec_port_7_port, CtlToDec_port_6_port, CtlToDec_port_5_port, 
      CtlToDec_port_4_port, CtlToDec_port_3_port, CtlToDec_port_2_port, 
      CtlToDec_port_1_port, CtlToDec_port_0_port, CtlToDec_port_notify, 
      DecToCtl_port_encType_2_port, DecToCtl_port_encType_1_port, 
      DecToCtl_port_encType_0_port, DecToCtl_port_imm_31_port, 
      DecToCtl_port_imm_30_port, DecToCtl_port_imm_29_port, 
      DecToCtl_port_imm_27_port, DecToCtl_port_imm_26_port, 
      DecToCtl_port_imm_22_port, DecToCtl_port_imm_21_port, 
      DecToCtl_port_imm_20_port, DecToCtl_port_imm_19_port, 
      DecToCtl_port_imm_17_port, DecToCtl_port_imm_15_port, 
      DecToCtl_port_imm_14_port, DecToCtl_port_imm_13_port, 
      DecToCtl_port_imm_12_port, DecToCtl_port_imm_11_port, 
      DecToCtl_port_imm_8_port, DecToCtl_port_imm_6_port, 
      DecToCtl_port_imm_4_port, DecToCtl_port_imm_2_port, 
      DecToCtl_port_imm_1_port, DecToCtl_port_imm_0_port, 
      DecToCtl_port_instrType_5_port, DecToCtl_port_instrType_4_port, 
      DecToCtl_port_instrType_3_port, DecToCtl_port_instrType_2_port, 
      DecToCtl_port_instrType_1_port, DecToCtl_port_instrType_0_port, 
      DecToCtl_port_rd_addr_4_port, DecToCtl_port_rd_addr_3_port, 
      DecToCtl_port_rd_addr_2_port, DecToCtl_port_rd_addr_1_port, 
      DecToCtl_port_rd_addr_0_port, DecToCtl_port_rs1_addr_4_port, 
      DecToCtl_port_rs1_addr_3_port, DecToCtl_port_rs1_addr_2_port, 
      DecToCtl_port_rs1_addr_1_port, DecToCtl_port_rs1_addr_0_port, 
      DecToCtl_port_rs2_addr_4_port, DecToCtl_port_rs2_addr_3_port, 
      DecToCtl_port_rs2_addr_2_port, DecToCtl_port_rs2_addr_1_port, 
      DecToCtl_port_rs2_addr_0_port, IF_ALUxN969, IF_ALUxN968, IF_ALUxN967, 
      IF_ALUxN966, IF_ALUxN965, IF_ALUxN964, IF_ALUxN963, IF_ALUxN962, 
      IF_ALUxN961, IF_ALUxN960, IF_ALUxN959, IF_ALUxN958, IF_ALUxN957, 
      IF_ALUxN956, IF_ALUxN955, IF_ALUxN954, IF_ALUxN953, IF_ALUxN952, 
      IF_ALUxN951, IF_ALUxN950, IF_ALUxN949, IF_ALUxN948, IF_ALUxN947, 
      IF_ALUxN946, IF_ALUxN945, IF_ALUxN944, IF_ALUxN943, IF_ALUxN942, 
      IF_ALUxN941, IF_ALUxN940, IF_ALUxN939, IF_ALUxN938, IF_ALUxN937, 
      IF_ALUxN142, IF_ALUxN141, IF_ALUxN140, IF_ALUxN139, IF_ALUxN138, 
      IF_ALUxN137, IF_ALUxN136, IF_ALUxN135, IF_ALUxN134, IF_ALUxN133, 
      IF_ALUxN132, IF_ALUxN131, IF_ALUxN130, IF_ALUxN129, IF_ALUxN128, 
      IF_ALUxN127, IF_ALUxN126, IF_ALUxN125, IF_ALUxN124, IF_ALUxN123, 
      IF_ALUxN122, IF_ALUxN121, IF_ALUxN120, IF_ALUxN119, IF_ALUxN118, 
      IF_ALUxN117, IF_ALUxN116, IF_ALUxN115, IF_ALUxN114, IF_ALUxN113, 
      IF_ALUxN112, IF_CPathxN2396, IF_CPathxN2394, IF_CPathxN2393, 
      IF_CPathxN2316, IF_CPathxN2310, IF_CPathxN2309, IF_CPathxN2308, 
      IF_CPathxN2274, IF_CPathxN2273, IF_CPathxN2271, IF_CPathxN2270, 
      IF_CPathxN2269, IF_CPathxN2268, IF_CPathxN2267, IF_CPathxN2266, 
      IF_CPathxN2265, IF_CPathxN2264, IF_CPathxN2263, IF_CPathxN2262, 
      IF_CPathxN2261, IF_CPathxN2260, IF_CPathxN2259, IF_CPathxN2258, 
      IF_CPathxN2257, IF_CPathxN2256, IF_CPathxN2255, IF_CPathxN2254, 
      IF_CPathxN2253, IF_CPathxN2252, IF_CPathxN2251, IF_CPathxN2250, 
      IF_CPathxN2249, IF_CPathxN2248, IF_CPathxN2247, IF_CPathxN2246, 
      IF_CPathxN2245, IF_CPathxN2244, IF_CPathxN2243, IF_CPathxN2242, 
      IF_CPathxN2235, IF_CPathxN2233, IF_CPathxN2232, IF_CPathxN2231, 
      IF_CPathxN2230, IF_CPathxN2229, IF_CPathxN2228, IF_CPathxN2227, 
      IF_CPathxN2226, IF_CPathxN2225, IF_CPathxN2224, IF_CPathxN2223, 
      IF_CPathxN2222, IF_CPathxN2221, IF_CPathxN2220, IF_CPathxN2219, 
      IF_CPathxN2218, IF_CPathxN2217, IF_CPathxN2216, IF_CPathxN2215, 
      IF_CPathxN2214, IF_CPathxN2213, IF_CPathxN2212, IF_CPathxN2211, 
      IF_CPathxN2210, IF_CPathxN2209, IF_CPathxN2208, IF_CPathxN2207, 
      IF_CPathxN2206, IF_CPathxN2205, IF_CPathxN2204, IF_CPathxN2203, 
      IF_CPathxN2202, IF_CPathxN2201, IF_CPathxN2200, IF_CPathxN2199, 
      IF_CPathxN2198, IF_CPathxN2197, IF_CPathxN2196, IF_CPathxN2195, 
      IF_CPathxN2194, IF_CPathxN2193, IF_CPathxN2192, IF_CPathxN2191, 
      IF_CPathxN2190, IF_CPathxN2186, IF_CPathxN2183, IF_CPathxN2182, 
      IF_CPathxN2181, IF_CPathxN2176, IF_CPathxN2174, IF_CPathxN2168, 
      IF_CPathxN2167, IF_CPathxN2165, IF_CPathxN2163, IF_CPathxN2162, 
      IF_CPathxN2161, IF_CPathxN2160, IF_CPathxN2159, IF_CPathxN2158, 
      IF_CPathxN2157, IF_CPathxN2155, IF_CPathxN2154, IF_CPathxN2153, 
      IF_CPathxN2152, IF_CPathxN2151, IF_CPathxN2150, IF_CPathxN2149, 
      IF_CPathxN2148, IF_CPathxN2147, IF_CPathxN2146, IF_CPathxN2145, 
      IF_CPathxN2144, IF_CPathxN2143, IF_CPathxN2142, IF_CPathxN2141, 
      IF_CPathxN2140, IF_CPathxN2139, IF_CPathxN2138, IF_CPathxN2137, 
      IF_CPathxN2136, IF_CPathxN2135, IF_CPathxN2134, IF_CPathxN2133, 
      IF_CPathxN2132, IF_CPathxN2131, IF_CPathxN2130, IF_CPathxN2129, 
      IF_CPathxN2128, IF_CPathxN2127, IF_CPathxN2126, IF_CPathxN2125, 
      IF_CPathxN2124, IF_CPathxN2096, IF_CPathxN2095, IF_CPathxN2094, 
      IF_CPathxN2092, IF_CPathxN2091, IF_CPathxN2090, IF_CPathxN2088, 
      IF_CPathxN2087, IF_CPathxN2086, IF_CPathxN2085, IF_CPathxN2084, 
      IF_CPathxN2083, IF_CPathxN2082, IF_CPathxN2081, IF_CPathxN2080, 
      IF_CPathxN2079, IF_CPathxN2078, IF_CPathxN2044, IF_CPathxN2038, 
      IF_CPathxN2037, IF_CPathxN2036, IF_CPathxN2035, IF_CPathxN2034, 
      IF_CPathxN2033, IF_CPathxN2032, IF_CPathxN1967, IF_CPathxN1966, 
      IF_CPathxN1965, IF_CPathxN1964, IF_CPathxN1963, IF_CPathxN1962, 
      IF_CPathxN1961, IF_CPathxN1960, IF_CPathxN1959, IF_CPathxN1958, 
      IF_CPathxN1957, IF_CPathxN1956, IF_CPathxN1955, IF_CPathxN1954, 
      IF_CPathxN1953, IF_CPathxN1952, IF_CPathxN1951, IF_CPathxN1950, 
      IF_CPathxN1949, IF_CPathxN1948, IF_CPathxN1947, IF_CPathxN1946, 
      IF_CPathxN1945, IF_CPathxN1944, IF_CPathxN1943, IF_CPathxN1942, 
      IF_CPathxN1941, IF_CPathxN1940, IF_CPathxN1939, IF_CPathxN1938, 
      IF_CPathxN1937, IF_CPathxN1936, IF_CPathxN1935, IF_CPathxN1932, 
      IF_CPathxN1930, IF_CPathxN1892, IF_CPathxN1891, IF_CPathxN1890, 
      IF_CPathxN1889, IF_CPathxN1888, IF_CPathxN1887, IF_CPathxN1886, 
      IF_CPathxN1885, IF_CPathxN1884, IF_CPathxN1883, IF_CPathxN1882, 
      IF_CPathxN1881, IF_CPathxN1880, IF_CPathxN1879, IF_CPathxN1878, 
      IF_CPathxN1877, IF_CPathxN1876, IF_CPathxN1875, IF_CPathxN1874, 
      IF_CPathxN1873, IF_CPathxN1872, IF_CPathxN1871, IF_CPathxN1870, 
      IF_CPathxN1869, IF_CPathxN1868, IF_CPathxN1867, IF_CPathxN1866, 
      IF_CPathxN1865, IF_CPathxN1864, IF_CPathxN1863, IF_CPathxN1862, 
      IF_CPathxN1861, IF_CPathxN1860, IF_CPathxN1859, IF_CPathxN1858, 
      IF_CPathxN1856, IF_CPathxN1854, IF_CPathxN1668, IF_CPathxN1667, 
      IF_CPathxN1665, IF_CPathxN1664, IF_CPathxN1631, IF_CPathxN1630, 
      IF_CPathxN1629, IF_CPathxN1628, IF_CPathxN896, IF_CPathxN895, 
      IF_CPathxN894, IF_CPathxN893, IF_CPathxN892, IF_CPathxN891, IF_CPathxN890
      , IF_CPathxN889, IF_CPathxN888, IF_CPathxN887, IF_CPathxN886, 
      IF_CPathxN885, IF_CPathxN884, IF_CPathxN883, IF_CPathxN882, IF_CPathxN881
      , IF_CPathxN880, IF_CPathxN879, IF_CPathxN878, IF_CPathxN877, 
      IF_CPathxN876, IF_CPathxN875, IF_CPathxN874, IF_CPathxN873, IF_CPathxN872
      , IF_CPathxN871, IF_CPathxN870, IF_CPathxN869, IF_CPathxN868, 
      IF_CPathxN867, IF_CPathxN866, IF_CPathxwb_sel_signal_0_port, 
      IF_CPathxwb_sel_signal_1_port, IF_CPathxwb_en_signal, 
      IF_CPathxreg_rd_en_signal, IF_CPathxpc_reg_signal_0_port, 
      IF_CPathxpc_reg_signal_1_port, IF_CPathxpc_reg_signal_2_port, 
      IF_CPathxpc_reg_signal_3_port, IF_CPathxpc_reg_signal_4_port, 
      IF_CPathxpc_reg_signal_5_port, IF_CPathxpc_reg_signal_6_port, 
      IF_CPathxpc_reg_signal_7_port, IF_CPathxpc_reg_signal_8_port, 
      IF_CPathxpc_reg_signal_9_port, IF_CPathxpc_reg_signal_10_port, 
      IF_CPathxpc_reg_signal_11_port, IF_CPathxpc_reg_signal_12_port, 
      IF_CPathxpc_reg_signal_13_port, IF_CPathxpc_reg_signal_14_port, 
      IF_CPathxpc_reg_signal_15_port, IF_CPathxpc_reg_signal_16_port, 
      IF_CPathxpc_reg_signal_17_port, IF_CPathxpc_reg_signal_18_port, 
      IF_CPathxpc_reg_signal_19_port, IF_CPathxpc_reg_signal_20_port, 
      IF_CPathxpc_reg_signal_21_port, IF_CPathxpc_reg_signal_22_port, 
      IF_CPathxpc_reg_signal_23_port, IF_CPathxpc_reg_signal_24_port, 
      IF_CPathxpc_reg_signal_25_port, IF_CPathxpc_reg_signal_26_port, 
      IF_CPathxpc_reg_signal_27_port, IF_CPathxpc_reg_signal_28_port, 
      IF_CPathxpc_reg_signal_29_port, IF_CPathxpc_reg_signal_30_port, 
      IF_CPathxpc_reg_signal_31_port, IF_CPathxpc_next_signal_0_port, 
      IF_CPathxpc_next_signal_1_port, IF_CPathxpc_next_signal_2_port, 
      IF_CPathxpc_next_signal_3_port, IF_CPathxpc_next_signal_4_port, 
      IF_CPathxpc_next_signal_5_port, IF_CPathxpc_next_signal_6_port, 
      IF_CPathxpc_next_signal_7_port, IF_CPathxpc_next_signal_8_port, 
      IF_CPathxpc_next_signal_9_port, IF_CPathxpc_next_signal_10_port, 
      IF_CPathxpc_next_signal_11_port, IF_CPathxpc_next_signal_12_port, 
      IF_CPathxpc_next_signal_13_port, IF_CPathxpc_next_signal_14_port, 
      IF_CPathxpc_next_signal_15_port, IF_CPathxpc_next_signal_16_port, 
      IF_CPathxpc_next_signal_17_port, IF_CPathxpc_next_signal_18_port, 
      IF_CPathxpc_next_signal_19_port, IF_CPathxpc_next_signal_20_port, 
      IF_CPathxpc_next_signal_21_port, IF_CPathxpc_next_signal_22_port, 
      IF_CPathxpc_next_signal_23_port, IF_CPathxpc_next_signal_24_port, 
      IF_CPathxpc_next_signal_25_port, IF_CPathxpc_next_signal_26_port, 
      IF_CPathxpc_next_signal_27_port, IF_CPathxpc_next_signal_28_port, 
      IF_CPathxpc_next_signal_29_port, IF_CPathxpc_next_signal_30_port, 
      IF_CPathxpc_next_signal_31_port, IF_CPathxmemoryAccess_signal_mask_0_port
      , IF_CPathxmemoryAccess_signal_mask_1_port, 
      IF_CPathxmemoryAccess_signal_mask_2_port, IF_CPathxmem_en_signal, 
      IF_CPathxMemToCtl_data_signal_0_port, 
      IF_CPathxMemToCtl_data_signal_1_port, 
      IF_CPathxMemToCtl_data_signal_2_port, 
      IF_CPathxMemToCtl_data_signal_3_port, 
      IF_CPathxMemToCtl_data_signal_4_port, 
      IF_CPathxMemToCtl_data_signal_5_port, 
      IF_CPathxMemToCtl_data_signal_6_port, 
      IF_CPathxMemToCtl_data_signal_7_port, 
      IF_CPathxMemToCtl_data_signal_8_port, 
      IF_CPathxMemToCtl_data_signal_9_port, 
      IF_CPathxMemToCtl_data_signal_10_port, 
      IF_CPathxMemToCtl_data_signal_11_port, 
      IF_CPathxMemToCtl_data_signal_12_port, 
      IF_CPathxMemToCtl_data_signal_13_port, 
      IF_CPathxMemToCtl_data_signal_14_port, 
      IF_CPathxMemToCtl_data_signal_15_port, 
      IF_CPathxMemToCtl_data_signal_16_port, 
      IF_CPathxMemToCtl_data_signal_17_port, 
      IF_CPathxMemToCtl_data_signal_18_port, 
      IF_CPathxMemToCtl_data_signal_19_port, 
      IF_CPathxMemToCtl_data_signal_20_port, 
      IF_CPathxMemToCtl_data_signal_21_port, 
      IF_CPathxMemToCtl_data_signal_22_port, 
      IF_CPathxMemToCtl_data_signal_23_port, 
      IF_CPathxMemToCtl_data_signal_24_port, 
      IF_CPathxMemToCtl_data_signal_25_port, 
      IF_CPathxMemToCtl_data_signal_26_port, 
      IF_CPathxMemToCtl_data_signal_27_port, 
      IF_CPathxMemToCtl_data_signal_28_port, 
      IF_CPathxMemToCtl_data_signal_29_port, 
      IF_CPathxMemToCtl_data_signal_30_port, 
      IF_CPathxMemToCtl_data_signal_31_port, 
      IF_CPathxDecToCtl_data_signal_rd_addr_0_port, 
      IF_CPathxDecToCtl_data_signal_rd_addr_1_port, 
      IF_CPathxDecToCtl_data_signal_rd_addr_2_port, 
      IF_CPathxDecToCtl_data_signal_rd_addr_3_port, 
      IF_CPathxDecToCtl_data_signal_rd_addr_4_port, 
      IF_CPathxDecToCtl_data_signal_instrType_0_port, 
      IF_CPathxDecToCtl_data_signal_instrType_1_port, 
      IF_CPathxDecToCtl_data_signal_instrType_2_port, 
      IF_CPathxDecToCtl_data_signal_instrType_4_port, 
      IF_CPathxDecToCtl_data_signal_instrType_5_port, 
      IF_CPathxDecToCtl_data_signal_imm_0_port, 
      IF_CPathxDecToCtl_data_signal_imm_1_port, 
      IF_CPathxDecToCtl_data_signal_imm_2_port, 
      IF_CPathxDecToCtl_data_signal_imm_3_port, 
      IF_CPathxDecToCtl_data_signal_imm_4_port, 
      IF_CPathxDecToCtl_data_signal_imm_5_port, 
      IF_CPathxDecToCtl_data_signal_imm_6_port, 
      IF_CPathxDecToCtl_data_signal_imm_7_port, 
      IF_CPathxDecToCtl_data_signal_imm_8_port, 
      IF_CPathxDecToCtl_data_signal_imm_9_port, 
      IF_CPathxDecToCtl_data_signal_imm_10_port, 
      IF_CPathxDecToCtl_data_signal_imm_11_port, 
      IF_CPathxDecToCtl_data_signal_imm_12_port, 
      IF_CPathxDecToCtl_data_signal_imm_13_port, 
      IF_CPathxDecToCtl_data_signal_imm_14_port, 
      IF_CPathxDecToCtl_data_signal_imm_15_port, 
      IF_CPathxDecToCtl_data_signal_imm_16_port, 
      IF_CPathxDecToCtl_data_signal_imm_17_port, 
      IF_CPathxDecToCtl_data_signal_imm_18_port, 
      IF_CPathxDecToCtl_data_signal_imm_19_port, 
      IF_CPathxDecToCtl_data_signal_imm_20_port, 
      IF_CPathxDecToCtl_data_signal_imm_21_port, 
      IF_CPathxDecToCtl_data_signal_imm_22_port, 
      IF_CPathxDecToCtl_data_signal_imm_23_port, 
      IF_CPathxDecToCtl_data_signal_imm_24_port, 
      IF_CPathxDecToCtl_data_signal_imm_25_port, 
      IF_CPathxDecToCtl_data_signal_imm_26_port, 
      IF_CPathxDecToCtl_data_signal_imm_27_port, 
      IF_CPathxDecToCtl_data_signal_imm_28_port, 
      IF_CPathxDecToCtl_data_signal_imm_29_port, 
      IF_CPathxDecToCtl_data_signal_imm_30_port, 
      IF_CPathxDecToCtl_data_signal_imm_31_port, IF_CPathxbr_en_signal, 
      IF_CPathxRegsToCtl_data_signal_contents1_0_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_1_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_2_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_3_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_4_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_5_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_6_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_7_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_8_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_9_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_10_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_11_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_12_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_13_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_14_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_15_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_16_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_17_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_18_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_19_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_20_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_21_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_22_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_23_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_24_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_25_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_26_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_27_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_28_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_29_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_30_port, 
      IF_CPathxRegsToCtl_data_signal_contents1_31_port, 
      IF_CPathxCtlToRegs_data_signal_src2_0_port, 
      IF_CPathxCtlToRegs_data_signal_src2_1_port, 
      IF_CPathxCtlToRegs_data_signal_src2_2_port, 
      IF_CPathxCtlToRegs_data_signal_src2_3_port, 
      IF_CPathxCtlToRegs_data_signal_src2_4_port, 
      IF_CPathxCtlToRegs_data_signal_src1_0_port, 
      IF_CPathxCtlToRegs_data_signal_src1_1_port, 
      IF_CPathxCtlToRegs_data_signal_src1_2_port, 
      IF_CPathxCtlToRegs_data_signal_src1_3_port, 
      IF_CPathxCtlToRegs_data_signal_src1_4_port, 
      IF_CPathxCtlToRegs_data_signal_dst_0_port, 
      IF_CPathxCtlToRegs_data_signal_dst_1_port, 
      IF_CPathxCtlToRegs_data_signal_dst_2_port, 
      IF_CPathxCtlToRegs_data_signal_dst_3_port, 
      IF_CPathxCtlToRegs_data_signal_dst_4_port, 
      IF_CPathxCtlToALU_data_signal_op2_sel_0_port, 
      IF_CPathxCtlToALU_data_signal_op2_sel_1_port, 
      IF_CPathxCtlToALU_data_signal_op1_sel_0_port, 
      IF_CPathxCtlToALU_data_signal_op1_sel_1_port, 
      IF_CPathxCtlToALU_data_signal_alu_fun_0_port, 
      IF_CPathxCtlToALU_data_signal_alu_fun_1_port, 
      IF_CPathxCtlToALU_data_signal_alu_fun_2_port, 
      IF_CPathxCtlToALU_data_signal_alu_fun_3_port, 
      IF_CPathxALUtoCtl_data_signal_0_port, 
      IF_CPathxALUtoCtl_data_signal_1_port, 
      IF_CPathxALUtoCtl_data_signal_2_port, 
      IF_CPathxALUtoCtl_data_signal_3_port, 
      IF_CPathxALUtoCtl_data_signal_4_port, 
      IF_CPathxALUtoCtl_data_signal_5_port, 
      IF_CPathxALUtoCtl_data_signal_6_port, 
      IF_CPathxALUtoCtl_data_signal_7_port, 
      IF_CPathxALUtoCtl_data_signal_8_port, 
      IF_CPathxALUtoCtl_data_signal_9_port, 
      IF_CPathxALUtoCtl_data_signal_10_port, 
      IF_CPathxALUtoCtl_data_signal_11_port, 
      IF_CPathxALUtoCtl_data_signal_12_port, 
      IF_CPathxALUtoCtl_data_signal_13_port, 
      IF_CPathxALUtoCtl_data_signal_14_port, 
      IF_CPathxALUtoCtl_data_signal_15_port, 
      IF_CPathxALUtoCtl_data_signal_16_port, 
      IF_CPathxALUtoCtl_data_signal_17_port, 
      IF_CPathxALUtoCtl_data_signal_18_port, 
      IF_CPathxALUtoCtl_data_signal_19_port, 
      IF_CPathxALUtoCtl_data_signal_20_port, 
      IF_CPathxALUtoCtl_data_signal_21_port, 
      IF_CPathxALUtoCtl_data_signal_22_port, 
      IF_CPathxALUtoCtl_data_signal_23_port, 
      IF_CPathxALUtoCtl_data_signal_24_port, 
      IF_CPathxALUtoCtl_data_signal_25_port, 
      IF_CPathxALUtoCtl_data_signal_26_port, 
      IF_CPathxALUtoCtl_data_signal_27_port, 
      IF_CPathxALUtoCtl_data_signal_28_port, 
      IF_CPathxALUtoCtl_data_signal_29_port, 
      IF_CPathxALUtoCtl_data_signal_30_port, 
      IF_CPathxALUtoCtl_data_signal_31_port, IF_CPathxsection_0_port, 
      IF_CPathxsection_2_port, IF_CPathxsection_3_port, IF_DecoderxN606, 
      IF_DecoderxN605, IF_DecoderxN604, IF_DecoderxN603, IF_DecoderxN602, 
      IF_DecoderxN601, IF_DecoderxN600, IF_DecoderxN599, IF_DecoderxN598, 
      IF_DecoderxN597, IF_DecoderxN596, IF_DecoderxN595, IF_DecoderxN594, 
      IF_DecoderxN593, IF_DecoderxN592, IF_DecoderxN591, IF_DecoderxN590, 
      IF_DecoderxN589, IF_DecoderxN588, IF_DecoderxN587, IF_DecoderxN586, 
      IF_DecoderxN585, IF_DecoderxN552, IF_DecoderxN551, IF_DecoderxN550, 
      IF_DecoderxN549, IF_RegsxN721, IF_RegsxN720, IF_RegsxN719, IF_RegsxN718, 
      IF_RegsxN717, IF_RegsxN716, IF_RegsxN715, IF_RegsxN714, IF_RegsxN713, 
      IF_RegsxN712, IF_RegsxN711, IF_RegsxN710, IF_RegsxN709, IF_RegsxN708, 
      IF_RegsxN707, IF_RegsxN706, IF_RegsxN705, IF_RegsxN704, IF_RegsxN703, 
      IF_RegsxN702, IF_RegsxN701, IF_RegsxN700, IF_RegsxN699, IF_RegsxN698, 
      IF_RegsxN697, IF_RegsxN696, IF_RegsxN695, IF_RegsxN694, IF_RegsxN693, 
      IF_RegsxN692, IF_RegsxN691, IF_RegsxN690, IF_RegsxN689, IF_RegsxN688, 
      IF_RegsxN687, IF_RegsxN686, IF_RegsxN685, IF_RegsxN684, IF_RegsxN683, 
      IF_RegsxN682, IF_RegsxN681, IF_RegsxN680, IF_RegsxN679, IF_RegsxN678, 
      IF_RegsxN677, IF_RegsxN676, IF_RegsxN675, IF_RegsxN674, IF_RegsxN673, 
      IF_RegsxN672, IF_RegsxN671, IF_RegsxN670, IF_RegsxN669, IF_RegsxN668, 
      IF_RegsxN667, IF_RegsxN666, IF_RegsxN665, IF_RegsxN664, IF_RegsxN663, 
      IF_RegsxN662, IF_RegsxN661, IF_RegsxN660, IF_RegsxN659, IF_RegsxN658, 
      IF_RegsxN657, IF_RegsxN656, IF_RegsxN655, IF_RegsxN654, IF_RegsxN653, 
      IF_RegsxN652, IF_RegsxN651, IF_RegsxN650, IF_RegsxN649, IF_RegsxN648, 
      IF_RegsxN647, IF_RegsxN646, IF_RegsxN645, IF_RegsxN644, IF_RegsxN643, 
      IF_RegsxN642, IF_RegsxN641, IF_RegsxN640, IF_RegsxN639, IF_RegsxN638, 
      IF_RegsxN637, IF_RegsxN636, IF_RegsxN635, IF_RegsxN634, IF_RegsxN633, 
      IF_RegsxN632, IF_RegsxN631, IF_RegsxN630, IF_RegsxN629, IF_RegsxN628, 
      IF_RegsxN627, IF_RegsxN626, IF_RegsxN625, IF_RegsxN624, IF_RegsxN623, 
      IF_RegsxN622, IF_RegsxN621, IF_RegsxN620, IF_RegsxN619, IF_RegsxN618, 
      IF_RegsxN617, IF_RegsxN616, IF_RegsxN615, IF_RegsxN614, IF_RegsxN613, 
      IF_RegsxN612, IF_RegsxN611, IF_RegsxN610, IF_RegsxN609, IF_RegsxN608, 
      IF_RegsxN607, IF_RegsxN606, IF_RegsxN605, IF_RegsxN604, IF_RegsxN603, 
      IF_RegsxN602, IF_RegsxN601, IF_RegsxN600, IF_RegsxN599, IF_RegsxN598, 
      IF_RegsxN597, IF_RegsxN596, IF_RegsxN595, IF_RegsxN594, 
      IF_Regsxreg_file_0_port, IF_Regsxreg_file_1_port, IF_Regsxreg_file_2_port
      , IF_Regsxreg_file_3_port, IF_Regsxreg_file_4_port, 
      IF_Regsxreg_file_5_port, IF_Regsxreg_file_6_port, IF_Regsxreg_file_7_port
      , IF_Regsxreg_file_8_port, IF_Regsxreg_file_9_port, 
      IF_Regsxreg_file_10_port, IF_Regsxreg_file_11_port, 
      IF_Regsxreg_file_12_port, IF_Regsxreg_file_13_port, 
      IF_Regsxreg_file_14_port, IF_Regsxreg_file_15_port, 
      IF_Regsxreg_file_16_port, IF_Regsxreg_file_17_port, 
      IF_Regsxreg_file_18_port, IF_Regsxreg_file_19_port, 
      IF_Regsxreg_file_20_port, IF_Regsxreg_file_21_port, 
      IF_Regsxreg_file_22_port, IF_Regsxreg_file_23_port, 
      IF_Regsxreg_file_24_port, IF_Regsxreg_file_25_port, 
      IF_Regsxreg_file_26_port, IF_Regsxreg_file_27_port, 
      IF_Regsxreg_file_28_port, IF_Regsxreg_file_29_port, 
      IF_Regsxreg_file_30_port, IF_Regsxreg_file_31_port, 
      IF_Regsxreg_file_32_port, IF_Regsxreg_file_33_port, 
      IF_Regsxreg_file_34_port, IF_Regsxreg_file_35_port, 
      IF_Regsxreg_file_36_port, IF_Regsxreg_file_37_port, 
      IF_Regsxreg_file_38_port, IF_Regsxreg_file_39_port, 
      IF_Regsxreg_file_40_port, IF_Regsxreg_file_41_port, 
      IF_Regsxreg_file_42_port, IF_Regsxreg_file_43_port, 
      IF_Regsxreg_file_44_port, IF_Regsxreg_file_45_port, 
      IF_Regsxreg_file_46_port, IF_Regsxreg_file_47_port, 
      IF_Regsxreg_file_48_port, IF_Regsxreg_file_49_port, 
      IF_Regsxreg_file_50_port, IF_Regsxreg_file_51_port, 
      IF_Regsxreg_file_52_port, IF_Regsxreg_file_53_port, 
      IF_Regsxreg_file_54_port, IF_Regsxreg_file_55_port, 
      IF_Regsxreg_file_56_port, IF_Regsxreg_file_57_port, 
      IF_Regsxreg_file_58_port, IF_Regsxreg_file_59_port, 
      IF_Regsxreg_file_60_port, IF_Regsxreg_file_61_port, 
      IF_Regsxreg_file_62_port, IF_Regsxreg_file_63_port, 
      IF_Regsxreg_file_64_port, IF_Regsxreg_file_65_port, 
      IF_Regsxreg_file_66_port, IF_Regsxreg_file_67_port, 
      IF_Regsxreg_file_68_port, IF_Regsxreg_file_69_port, 
      IF_Regsxreg_file_70_port, IF_Regsxreg_file_71_port, 
      IF_Regsxreg_file_72_port, IF_Regsxreg_file_73_port, 
      IF_Regsxreg_file_74_port, IF_Regsxreg_file_75_port, 
      IF_Regsxreg_file_76_port, IF_Regsxreg_file_77_port, 
      IF_Regsxreg_file_78_port, IF_Regsxreg_file_79_port, 
      IF_Regsxreg_file_80_port, IF_Regsxreg_file_81_port, 
      IF_Regsxreg_file_82_port, IF_Regsxreg_file_83_port, 
      IF_Regsxreg_file_84_port, IF_Regsxreg_file_85_port, 
      IF_Regsxreg_file_86_port, IF_Regsxreg_file_87_port, 
      IF_Regsxreg_file_88_port, IF_Regsxreg_file_89_port, 
      IF_Regsxreg_file_90_port, IF_Regsxreg_file_91_port, 
      IF_Regsxreg_file_92_port, IF_Regsxreg_file_93_port, 
      IF_Regsxreg_file_94_port, IF_Regsxreg_file_95_port, 
      IF_Regsxreg_file_96_port, IF_Regsxreg_file_97_port, 
      IF_Regsxreg_file_98_port, IF_Regsxreg_file_99_port, 
      IF_Regsxreg_file_100_port, IF_Regsxreg_file_101_port, 
      IF_Regsxreg_file_102_port, IF_Regsxreg_file_103_port, 
      IF_Regsxreg_file_104_port, IF_Regsxreg_file_105_port, 
      IF_Regsxreg_file_106_port, IF_Regsxreg_file_107_port, 
      IF_Regsxreg_file_108_port, IF_Regsxreg_file_109_port, 
      IF_Regsxreg_file_110_port, IF_Regsxreg_file_111_port, 
      IF_Regsxreg_file_112_port, IF_Regsxreg_file_113_port, 
      IF_Regsxreg_file_114_port, IF_Regsxreg_file_115_port, 
      IF_Regsxreg_file_116_port, IF_Regsxreg_file_117_port, 
      IF_Regsxreg_file_118_port, IF_Regsxreg_file_119_port, 
      IF_Regsxreg_file_120_port, IF_Regsxreg_file_121_port, 
      IF_Regsxreg_file_122_port, IF_Regsxreg_file_123_port, 
      IF_Regsxreg_file_124_port, IF_Regsxreg_file_125_port, 
      IF_Regsxreg_file_126_port, IF_Regsxreg_file_127_port, 
      IF_Regsxreg_file_128_port, IF_Regsxreg_file_129_port, 
      IF_Regsxreg_file_130_port, IF_Regsxreg_file_131_port, 
      IF_Regsxreg_file_132_port, IF_Regsxreg_file_133_port, 
      IF_Regsxreg_file_134_port, IF_Regsxreg_file_135_port, 
      IF_Regsxreg_file_136_port, IF_Regsxreg_file_137_port, 
      IF_Regsxreg_file_138_port, IF_Regsxreg_file_139_port, 
      IF_Regsxreg_file_140_port, IF_Regsxreg_file_141_port, 
      IF_Regsxreg_file_142_port, IF_Regsxreg_file_143_port, 
      IF_Regsxreg_file_144_port, IF_Regsxreg_file_145_port, 
      IF_Regsxreg_file_146_port, IF_Regsxreg_file_147_port, 
      IF_Regsxreg_file_148_port, IF_Regsxreg_file_149_port, 
      IF_Regsxreg_file_150_port, IF_Regsxreg_file_151_port, 
      IF_Regsxreg_file_152_port, IF_Regsxreg_file_153_port, 
      IF_Regsxreg_file_154_port, IF_Regsxreg_file_155_port, 
      IF_Regsxreg_file_156_port, IF_Regsxreg_file_157_port, 
      IF_Regsxreg_file_158_port, IF_Regsxreg_file_159_port, 
      IF_Regsxreg_file_160_port, IF_Regsxreg_file_161_port, 
      IF_Regsxreg_file_162_port, IF_Regsxreg_file_163_port, 
      IF_Regsxreg_file_164_port, IF_Regsxreg_file_165_port, 
      IF_Regsxreg_file_166_port, IF_Regsxreg_file_167_port, 
      IF_Regsxreg_file_168_port, IF_Regsxreg_file_169_port, 
      IF_Regsxreg_file_170_port, IF_Regsxreg_file_171_port, 
      IF_Regsxreg_file_172_port, IF_Regsxreg_file_173_port, 
      IF_Regsxreg_file_174_port, IF_Regsxreg_file_175_port, 
      IF_Regsxreg_file_176_port, IF_Regsxreg_file_177_port, 
      IF_Regsxreg_file_178_port, IF_Regsxreg_file_179_port, 
      IF_Regsxreg_file_180_port, IF_Regsxreg_file_181_port, 
      IF_Regsxreg_file_182_port, IF_Regsxreg_file_183_port, 
      IF_Regsxreg_file_184_port, IF_Regsxreg_file_185_port, 
      IF_Regsxreg_file_186_port, IF_Regsxreg_file_187_port, 
      IF_Regsxreg_file_188_port, IF_Regsxreg_file_189_port, 
      IF_Regsxreg_file_190_port, IF_Regsxreg_file_191_port, 
      IF_Regsxreg_file_192_port, IF_Regsxreg_file_193_port, 
      IF_Regsxreg_file_194_port, IF_Regsxreg_file_195_port, 
      IF_Regsxreg_file_196_port, IF_Regsxreg_file_197_port, 
      IF_Regsxreg_file_198_port, IF_Regsxreg_file_199_port, 
      IF_Regsxreg_file_200_port, IF_Regsxreg_file_201_port, 
      IF_Regsxreg_file_202_port, IF_Regsxreg_file_203_port, 
      IF_Regsxreg_file_204_port, IF_Regsxreg_file_205_port, 
      IF_Regsxreg_file_206_port, IF_Regsxreg_file_207_port, 
      IF_Regsxreg_file_208_port, IF_Regsxreg_file_209_port, 
      IF_Regsxreg_file_210_port, IF_Regsxreg_file_211_port, 
      IF_Regsxreg_file_212_port, IF_Regsxreg_file_213_port, 
      IF_Regsxreg_file_214_port, IF_Regsxreg_file_215_port, 
      IF_Regsxreg_file_216_port, IF_Regsxreg_file_217_port, 
      IF_Regsxreg_file_218_port, IF_Regsxreg_file_219_port, 
      IF_Regsxreg_file_220_port, IF_Regsxreg_file_221_port, 
      IF_Regsxreg_file_222_port, IF_Regsxreg_file_223_port, 
      IF_Regsxreg_file_224_port, IF_Regsxreg_file_225_port, 
      IF_Regsxreg_file_226_port, IF_Regsxreg_file_227_port, 
      IF_Regsxreg_file_228_port, IF_Regsxreg_file_229_port, 
      IF_Regsxreg_file_230_port, IF_Regsxreg_file_231_port, 
      IF_Regsxreg_file_232_port, IF_Regsxreg_file_233_port, 
      IF_Regsxreg_file_234_port, IF_Regsxreg_file_235_port, 
      IF_Regsxreg_file_236_port, IF_Regsxreg_file_237_port, 
      IF_Regsxreg_file_238_port, IF_Regsxreg_file_239_port, 
      IF_Regsxreg_file_240_port, IF_Regsxreg_file_241_port, 
      IF_Regsxreg_file_242_port, IF_Regsxreg_file_243_port, 
      IF_Regsxreg_file_244_port, IF_Regsxreg_file_245_port, 
      IF_Regsxreg_file_246_port, IF_Regsxreg_file_247_port, 
      IF_Regsxreg_file_248_port, IF_Regsxreg_file_249_port, 
      IF_Regsxreg_file_250_port, IF_Regsxreg_file_251_port, 
      IF_Regsxreg_file_252_port, IF_Regsxreg_file_253_port, 
      IF_Regsxreg_file_254_port, IF_Regsxreg_file_255_port, 
      IF_Regsxreg_file_256_port, IF_Regsxreg_file_257_port, 
      IF_Regsxreg_file_258_port, IF_Regsxreg_file_259_port, 
      IF_Regsxreg_file_260_port, IF_Regsxreg_file_261_port, 
      IF_Regsxreg_file_262_port, IF_Regsxreg_file_263_port, 
      IF_Regsxreg_file_264_port, IF_Regsxreg_file_265_port, 
      IF_Regsxreg_file_266_port, IF_Regsxreg_file_267_port, 
      IF_Regsxreg_file_268_port, IF_Regsxreg_file_269_port, 
      IF_Regsxreg_file_270_port, IF_Regsxreg_file_271_port, 
      IF_Regsxreg_file_272_port, IF_Regsxreg_file_273_port, 
      IF_Regsxreg_file_274_port, IF_Regsxreg_file_275_port, 
      IF_Regsxreg_file_276_port, IF_Regsxreg_file_277_port, 
      IF_Regsxreg_file_278_port, IF_Regsxreg_file_279_port, 
      IF_Regsxreg_file_280_port, IF_Regsxreg_file_281_port, 
      IF_Regsxreg_file_282_port, IF_Regsxreg_file_283_port, 
      IF_Regsxreg_file_284_port, IF_Regsxreg_file_285_port, 
      IF_Regsxreg_file_286_port, IF_Regsxreg_file_287_port, 
      IF_Regsxreg_file_288_port, IF_Regsxreg_file_289_port, 
      IF_Regsxreg_file_290_port, IF_Regsxreg_file_291_port, 
      IF_Regsxreg_file_292_port, IF_Regsxreg_file_293_port, 
      IF_Regsxreg_file_294_port, IF_Regsxreg_file_295_port, 
      IF_Regsxreg_file_296_port, IF_Regsxreg_file_297_port, 
      IF_Regsxreg_file_298_port, IF_Regsxreg_file_299_port, 
      IF_Regsxreg_file_300_port, IF_Regsxreg_file_301_port, 
      IF_Regsxreg_file_302_port, IF_Regsxreg_file_303_port, 
      IF_Regsxreg_file_304_port, IF_Regsxreg_file_305_port, 
      IF_Regsxreg_file_306_port, IF_Regsxreg_file_307_port, 
      IF_Regsxreg_file_308_port, IF_Regsxreg_file_309_port, 
      IF_Regsxreg_file_310_port, IF_Regsxreg_file_311_port, 
      IF_Regsxreg_file_312_port, IF_Regsxreg_file_313_port, 
      IF_Regsxreg_file_314_port, IF_Regsxreg_file_315_port, 
      IF_Regsxreg_file_316_port, IF_Regsxreg_file_317_port, 
      IF_Regsxreg_file_318_port, IF_Regsxreg_file_319_port, 
      IF_Regsxreg_file_320_port, IF_Regsxreg_file_321_port, 
      IF_Regsxreg_file_322_port, IF_Regsxreg_file_323_port, 
      IF_Regsxreg_file_324_port, IF_Regsxreg_file_325_port, 
      IF_Regsxreg_file_326_port, IF_Regsxreg_file_327_port, 
      IF_Regsxreg_file_328_port, IF_Regsxreg_file_329_port, 
      IF_Regsxreg_file_330_port, IF_Regsxreg_file_331_port, 
      IF_Regsxreg_file_332_port, IF_Regsxreg_file_333_port, 
      IF_Regsxreg_file_334_port, IF_Regsxreg_file_335_port, 
      IF_Regsxreg_file_336_port, IF_Regsxreg_file_337_port, 
      IF_Regsxreg_file_338_port, IF_Regsxreg_file_339_port, 
      IF_Regsxreg_file_340_port, IF_Regsxreg_file_341_port, 
      IF_Regsxreg_file_342_port, IF_Regsxreg_file_343_port, 
      IF_Regsxreg_file_344_port, IF_Regsxreg_file_345_port, 
      IF_Regsxreg_file_346_port, IF_Regsxreg_file_347_port, 
      IF_Regsxreg_file_348_port, IF_Regsxreg_file_349_port, 
      IF_Regsxreg_file_350_port, IF_Regsxreg_file_351_port, 
      IF_Regsxreg_file_352_port, IF_Regsxreg_file_353_port, 
      IF_Regsxreg_file_354_port, IF_Regsxreg_file_355_port, 
      IF_Regsxreg_file_356_port, IF_Regsxreg_file_357_port, 
      IF_Regsxreg_file_358_port, IF_Regsxreg_file_359_port, 
      IF_Regsxreg_file_360_port, IF_Regsxreg_file_361_port, 
      IF_Regsxreg_file_362_port, IF_Regsxreg_file_363_port, 
      IF_Regsxreg_file_364_port, IF_Regsxreg_file_365_port, 
      IF_Regsxreg_file_366_port, IF_Regsxreg_file_367_port, 
      IF_Regsxreg_file_368_port, IF_Regsxreg_file_369_port, 
      IF_Regsxreg_file_370_port, IF_Regsxreg_file_371_port, 
      IF_Regsxreg_file_372_port, IF_Regsxreg_file_373_port, 
      IF_Regsxreg_file_374_port, IF_Regsxreg_file_375_port, 
      IF_Regsxreg_file_376_port, IF_Regsxreg_file_377_port, 
      IF_Regsxreg_file_378_port, IF_Regsxreg_file_379_port, 
      IF_Regsxreg_file_380_port, IF_Regsxreg_file_381_port, 
      IF_Regsxreg_file_382_port, IF_Regsxreg_file_383_port, 
      IF_Regsxreg_file_384_port, IF_Regsxreg_file_385_port, 
      IF_Regsxreg_file_386_port, IF_Regsxreg_file_387_port, 
      IF_Regsxreg_file_388_port, IF_Regsxreg_file_389_port, 
      IF_Regsxreg_file_390_port, IF_Regsxreg_file_391_port, 
      IF_Regsxreg_file_392_port, IF_Regsxreg_file_393_port, 
      IF_Regsxreg_file_394_port, IF_Regsxreg_file_395_port, 
      IF_Regsxreg_file_396_port, IF_Regsxreg_file_397_port, 
      IF_Regsxreg_file_398_port, IF_Regsxreg_file_399_port, 
      IF_Regsxreg_file_400_port, IF_Regsxreg_file_401_port, 
      IF_Regsxreg_file_402_port, IF_Regsxreg_file_403_port, 
      IF_Regsxreg_file_404_port, IF_Regsxreg_file_405_port, 
      IF_Regsxreg_file_406_port, IF_Regsxreg_file_407_port, 
      IF_Regsxreg_file_408_port, IF_Regsxreg_file_409_port, 
      IF_Regsxreg_file_410_port, IF_Regsxreg_file_411_port, 
      IF_Regsxreg_file_412_port, IF_Regsxreg_file_413_port, 
      IF_Regsxreg_file_414_port, IF_Regsxreg_file_415_port, 
      IF_Regsxreg_file_416_port, IF_Regsxreg_file_417_port, 
      IF_Regsxreg_file_418_port, IF_Regsxreg_file_419_port, 
      IF_Regsxreg_file_420_port, IF_Regsxreg_file_421_port, 
      IF_Regsxreg_file_422_port, IF_Regsxreg_file_423_port, 
      IF_Regsxreg_file_424_port, IF_Regsxreg_file_425_port, 
      IF_Regsxreg_file_426_port, IF_Regsxreg_file_427_port, 
      IF_Regsxreg_file_428_port, IF_Regsxreg_file_429_port, 
      IF_Regsxreg_file_430_port, IF_Regsxreg_file_431_port, 
      IF_Regsxreg_file_432_port, IF_Regsxreg_file_433_port, 
      IF_Regsxreg_file_434_port, IF_Regsxreg_file_435_port, 
      IF_Regsxreg_file_436_port, IF_Regsxreg_file_437_port, 
      IF_Regsxreg_file_438_port, IF_Regsxreg_file_439_port, 
      IF_Regsxreg_file_440_port, IF_Regsxreg_file_441_port, 
      IF_Regsxreg_file_442_port, IF_Regsxreg_file_443_port, 
      IF_Regsxreg_file_444_port, IF_Regsxreg_file_445_port, 
      IF_Regsxreg_file_446_port, IF_Regsxreg_file_447_port, 
      IF_Regsxreg_file_448_port, IF_Regsxreg_file_449_port, 
      IF_Regsxreg_file_450_port, IF_Regsxreg_file_451_port, 
      IF_Regsxreg_file_452_port, IF_Regsxreg_file_453_port, 
      IF_Regsxreg_file_454_port, IF_Regsxreg_file_455_port, 
      IF_Regsxreg_file_456_port, IF_Regsxreg_file_457_port, 
      IF_Regsxreg_file_458_port, IF_Regsxreg_file_459_port, 
      IF_Regsxreg_file_460_port, IF_Regsxreg_file_461_port, 
      IF_Regsxreg_file_462_port, IF_Regsxreg_file_463_port, 
      IF_Regsxreg_file_464_port, IF_Regsxreg_file_465_port, 
      IF_Regsxreg_file_466_port, IF_Regsxreg_file_467_port, 
      IF_Regsxreg_file_468_port, IF_Regsxreg_file_469_port, 
      IF_Regsxreg_file_470_port, IF_Regsxreg_file_471_port, 
      IF_Regsxreg_file_472_port, IF_Regsxreg_file_473_port, 
      IF_Regsxreg_file_474_port, IF_Regsxreg_file_475_port, 
      IF_Regsxreg_file_476_port, IF_Regsxreg_file_477_port, 
      IF_Regsxreg_file_478_port, IF_Regsxreg_file_479_port, 
      IF_Regsxreg_file_480_port, IF_Regsxreg_file_481_port, 
      IF_Regsxreg_file_482_port, IF_Regsxreg_file_483_port, 
      IF_Regsxreg_file_484_port, IF_Regsxreg_file_485_port, 
      IF_Regsxreg_file_486_port, IF_Regsxreg_file_487_port, 
      IF_Regsxreg_file_488_port, IF_Regsxreg_file_489_port, 
      IF_Regsxreg_file_490_port, IF_Regsxreg_file_491_port, 
      IF_Regsxreg_file_492_port, IF_Regsxreg_file_493_port, 
      IF_Regsxreg_file_494_port, IF_Regsxreg_file_495_port, 
      IF_Regsxreg_file_496_port, IF_Regsxreg_file_497_port, 
      IF_Regsxreg_file_498_port, IF_Regsxreg_file_499_port, 
      IF_Regsxreg_file_500_port, IF_Regsxreg_file_501_port, 
      IF_Regsxreg_file_502_port, IF_Regsxreg_file_503_port, 
      IF_Regsxreg_file_504_port, IF_Regsxreg_file_505_port, 
      IF_Regsxreg_file_506_port, IF_Regsxreg_file_507_port, 
      IF_Regsxreg_file_508_port, IF_Regsxreg_file_509_port, 
      IF_Regsxreg_file_510_port, IF_Regsxreg_file_511_port, 
      IF_Regsxreg_file_512_port, IF_Regsxreg_file_513_port, 
      IF_Regsxreg_file_514_port, IF_Regsxreg_file_515_port, 
      IF_Regsxreg_file_516_port, IF_Regsxreg_file_517_port, 
      IF_Regsxreg_file_518_port, IF_Regsxreg_file_519_port, 
      IF_Regsxreg_file_520_port, IF_Regsxreg_file_521_port, 
      IF_Regsxreg_file_522_port, IF_Regsxreg_file_523_port, 
      IF_Regsxreg_file_524_port, IF_Regsxreg_file_525_port, 
      IF_Regsxreg_file_526_port, IF_Regsxreg_file_527_port, 
      IF_Regsxreg_file_528_port, IF_Regsxreg_file_529_port, 
      IF_Regsxreg_file_530_port, IF_Regsxreg_file_531_port, 
      IF_Regsxreg_file_532_port, IF_Regsxreg_file_533_port, 
      IF_Regsxreg_file_534_port, IF_Regsxreg_file_535_port, 
      IF_Regsxreg_file_536_port, IF_Regsxreg_file_537_port, 
      IF_Regsxreg_file_538_port, IF_Regsxreg_file_539_port, 
      IF_Regsxreg_file_540_port, IF_Regsxreg_file_541_port, 
      IF_Regsxreg_file_542_port, IF_Regsxreg_file_543_port, 
      IF_Regsxreg_file_544_port, IF_Regsxreg_file_545_port, 
      IF_Regsxreg_file_546_port, IF_Regsxreg_file_547_port, 
      IF_Regsxreg_file_548_port, IF_Regsxreg_file_549_port, 
      IF_Regsxreg_file_550_port, IF_Regsxreg_file_551_port, 
      IF_Regsxreg_file_552_port, IF_Regsxreg_file_553_port, 
      IF_Regsxreg_file_554_port, IF_Regsxreg_file_555_port, 
      IF_Regsxreg_file_556_port, IF_Regsxreg_file_557_port, 
      IF_Regsxreg_file_558_port, IF_Regsxreg_file_559_port, 
      IF_Regsxreg_file_560_port, IF_Regsxreg_file_561_port, 
      IF_Regsxreg_file_562_port, IF_Regsxreg_file_563_port, 
      IF_Regsxreg_file_564_port, IF_Regsxreg_file_565_port, 
      IF_Regsxreg_file_566_port, IF_Regsxreg_file_567_port, 
      IF_Regsxreg_file_568_port, IF_Regsxreg_file_569_port, 
      IF_Regsxreg_file_570_port, IF_Regsxreg_file_571_port, 
      IF_Regsxreg_file_572_port, IF_Regsxreg_file_573_port, 
      IF_Regsxreg_file_574_port, IF_Regsxreg_file_575_port, 
      IF_Regsxreg_file_576_port, IF_Regsxreg_file_577_port, 
      IF_Regsxreg_file_578_port, IF_Regsxreg_file_579_port, 
      IF_Regsxreg_file_580_port, IF_Regsxreg_file_581_port, 
      IF_Regsxreg_file_582_port, IF_Regsxreg_file_583_port, 
      IF_Regsxreg_file_584_port, IF_Regsxreg_file_585_port, 
      IF_Regsxreg_file_586_port, IF_Regsxreg_file_587_port, 
      IF_Regsxreg_file_588_port, IF_Regsxreg_file_589_port, 
      IF_Regsxreg_file_590_port, IF_Regsxreg_file_591_port, 
      IF_Regsxreg_file_592_port, IF_Regsxreg_file_593_port, 
      IF_Regsxreg_file_594_port, IF_Regsxreg_file_595_port, 
      IF_Regsxreg_file_596_port, IF_Regsxreg_file_597_port, 
      IF_Regsxreg_file_598_port, IF_Regsxreg_file_599_port, 
      IF_Regsxreg_file_600_port, IF_Regsxreg_file_601_port, 
      IF_Regsxreg_file_602_port, IF_Regsxreg_file_603_port, 
      IF_Regsxreg_file_604_port, IF_Regsxreg_file_605_port, 
      IF_Regsxreg_file_606_port, IF_Regsxreg_file_607_port, 
      IF_Regsxreg_file_608_port, IF_Regsxreg_file_609_port, 
      IF_Regsxreg_file_610_port, IF_Regsxreg_file_611_port, 
      IF_Regsxreg_file_612_port, IF_Regsxreg_file_613_port, 
      IF_Regsxreg_file_614_port, IF_Regsxreg_file_615_port, 
      IF_Regsxreg_file_616_port, IF_Regsxreg_file_617_port, 
      IF_Regsxreg_file_618_port, IF_Regsxreg_file_619_port, 
      IF_Regsxreg_file_620_port, IF_Regsxreg_file_621_port, 
      IF_Regsxreg_file_622_port, IF_Regsxreg_file_623_port, 
      IF_Regsxreg_file_624_port, IF_Regsxreg_file_625_port, 
      IF_Regsxreg_file_626_port, IF_Regsxreg_file_627_port, 
      IF_Regsxreg_file_628_port, IF_Regsxreg_file_629_port, 
      IF_Regsxreg_file_630_port, IF_Regsxreg_file_631_port, 
      IF_Regsxreg_file_632_port, IF_Regsxreg_file_633_port, 
      IF_Regsxreg_file_634_port, IF_Regsxreg_file_635_port, 
      IF_Regsxreg_file_636_port, IF_Regsxreg_file_637_port, 
      IF_Regsxreg_file_638_port, IF_Regsxreg_file_639_port, 
      IF_Regsxreg_file_640_port, IF_Regsxreg_file_641_port, 
      IF_Regsxreg_file_642_port, IF_Regsxreg_file_643_port, 
      IF_Regsxreg_file_644_port, IF_Regsxreg_file_645_port, 
      IF_Regsxreg_file_646_port, IF_Regsxreg_file_647_port, 
      IF_Regsxreg_file_648_port, IF_Regsxreg_file_649_port, 
      IF_Regsxreg_file_650_port, IF_Regsxreg_file_651_port, 
      IF_Regsxreg_file_652_port, IF_Regsxreg_file_653_port, 
      IF_Regsxreg_file_654_port, IF_Regsxreg_file_655_port, 
      IF_Regsxreg_file_656_port, IF_Regsxreg_file_657_port, 
      IF_Regsxreg_file_658_port, IF_Regsxreg_file_659_port, 
      IF_Regsxreg_file_660_port, IF_Regsxreg_file_661_port, 
      IF_Regsxreg_file_662_port, IF_Regsxreg_file_663_port, 
      IF_Regsxreg_file_664_port, IF_Regsxreg_file_665_port, 
      IF_Regsxreg_file_666_port, IF_Regsxreg_file_667_port, 
      IF_Regsxreg_file_668_port, IF_Regsxreg_file_669_port, 
      IF_Regsxreg_file_670_port, IF_Regsxreg_file_671_port, 
      IF_Regsxreg_file_672_port, IF_Regsxreg_file_673_port, 
      IF_Regsxreg_file_674_port, IF_Regsxreg_file_675_port, 
      IF_Regsxreg_file_676_port, IF_Regsxreg_file_677_port, 
      IF_Regsxreg_file_678_port, IF_Regsxreg_file_679_port, 
      IF_Regsxreg_file_680_port, IF_Regsxreg_file_681_port, 
      IF_Regsxreg_file_682_port, IF_Regsxreg_file_683_port, 
      IF_Regsxreg_file_684_port, IF_Regsxreg_file_685_port, 
      IF_Regsxreg_file_686_port, IF_Regsxreg_file_687_port, 
      IF_Regsxreg_file_688_port, IF_Regsxreg_file_689_port, 
      IF_Regsxreg_file_690_port, IF_Regsxreg_file_691_port, 
      IF_Regsxreg_file_692_port, IF_Regsxreg_file_693_port, 
      IF_Regsxreg_file_694_port, IF_Regsxreg_file_695_port, 
      IF_Regsxreg_file_696_port, IF_Regsxreg_file_697_port, 
      IF_Regsxreg_file_698_port, IF_Regsxreg_file_699_port, 
      IF_Regsxreg_file_700_port, IF_Regsxreg_file_701_port, 
      IF_Regsxreg_file_702_port, IF_Regsxreg_file_703_port, 
      IF_Regsxreg_file_704_port, IF_Regsxreg_file_705_port, 
      IF_Regsxreg_file_706_port, IF_Regsxreg_file_707_port, 
      IF_Regsxreg_file_708_port, IF_Regsxreg_file_709_port, 
      IF_Regsxreg_file_710_port, IF_Regsxreg_file_711_port, 
      IF_Regsxreg_file_712_port, IF_Regsxreg_file_713_port, 
      IF_Regsxreg_file_714_port, IF_Regsxreg_file_715_port, 
      IF_Regsxreg_file_716_port, IF_Regsxreg_file_717_port, 
      IF_Regsxreg_file_718_port, IF_Regsxreg_file_719_port, 
      IF_Regsxreg_file_720_port, IF_Regsxreg_file_721_port, 
      IF_Regsxreg_file_722_port, IF_Regsxreg_file_723_port, 
      IF_Regsxreg_file_724_port, IF_Regsxreg_file_725_port, 
      IF_Regsxreg_file_726_port, IF_Regsxreg_file_727_port, 
      IF_Regsxreg_file_728_port, IF_Regsxreg_file_729_port, 
      IF_Regsxreg_file_730_port, IF_Regsxreg_file_731_port, 
      IF_Regsxreg_file_732_port, IF_Regsxreg_file_733_port, 
      IF_Regsxreg_file_734_port, IF_Regsxreg_file_735_port, 
      IF_Regsxreg_file_736_port, IF_Regsxreg_file_737_port, 
      IF_Regsxreg_file_738_port, IF_Regsxreg_file_739_port, 
      IF_Regsxreg_file_740_port, IF_Regsxreg_file_741_port, 
      IF_Regsxreg_file_742_port, IF_Regsxreg_file_743_port, 
      IF_Regsxreg_file_744_port, IF_Regsxreg_file_745_port, 
      IF_Regsxreg_file_746_port, IF_Regsxreg_file_747_port, 
      IF_Regsxreg_file_748_port, IF_Regsxreg_file_749_port, 
      IF_Regsxreg_file_750_port, IF_Regsxreg_file_751_port, 
      IF_Regsxreg_file_752_port, IF_Regsxreg_file_753_port, 
      IF_Regsxreg_file_754_port, IF_Regsxreg_file_755_port, 
      IF_Regsxreg_file_756_port, IF_Regsxreg_file_757_port, 
      IF_Regsxreg_file_758_port, IF_Regsxreg_file_759_port, 
      IF_Regsxreg_file_760_port, IF_Regsxreg_file_761_port, 
      IF_Regsxreg_file_762_port, IF_Regsxreg_file_763_port, 
      IF_Regsxreg_file_764_port, IF_Regsxreg_file_765_port, 
      IF_Regsxreg_file_766_port, IF_Regsxreg_file_767_port, 
      IF_Regsxreg_file_768_port, IF_Regsxreg_file_769_port, 
      IF_Regsxreg_file_770_port, IF_Regsxreg_file_771_port, 
      IF_Regsxreg_file_772_port, IF_Regsxreg_file_773_port, 
      IF_Regsxreg_file_774_port, IF_Regsxreg_file_775_port, 
      IF_Regsxreg_file_776_port, IF_Regsxreg_file_777_port, 
      IF_Regsxreg_file_778_port, IF_Regsxreg_file_779_port, 
      IF_Regsxreg_file_780_port, IF_Regsxreg_file_781_port, 
      IF_Regsxreg_file_782_port, IF_Regsxreg_file_783_port, 
      IF_Regsxreg_file_784_port, IF_Regsxreg_file_785_port, 
      IF_Regsxreg_file_786_port, IF_Regsxreg_file_787_port, 
      IF_Regsxreg_file_788_port, IF_Regsxreg_file_789_port, 
      IF_Regsxreg_file_790_port, IF_Regsxreg_file_791_port, 
      IF_Regsxreg_file_792_port, IF_Regsxreg_file_793_port, 
      IF_Regsxreg_file_794_port, IF_Regsxreg_file_795_port, 
      IF_Regsxreg_file_796_port, IF_Regsxreg_file_797_port, 
      IF_Regsxreg_file_798_port, IF_Regsxreg_file_799_port, 
      IF_Regsxreg_file_800_port, IF_Regsxreg_file_801_port, 
      IF_Regsxreg_file_802_port, IF_Regsxreg_file_803_port, 
      IF_Regsxreg_file_804_port, IF_Regsxreg_file_805_port, 
      IF_Regsxreg_file_806_port, IF_Regsxreg_file_807_port, 
      IF_Regsxreg_file_808_port, IF_Regsxreg_file_809_port, 
      IF_Regsxreg_file_810_port, IF_Regsxreg_file_811_port, 
      IF_Regsxreg_file_812_port, IF_Regsxreg_file_813_port, 
      IF_Regsxreg_file_814_port, IF_Regsxreg_file_815_port, 
      IF_Regsxreg_file_816_port, IF_Regsxreg_file_817_port, 
      IF_Regsxreg_file_818_port, IF_Regsxreg_file_819_port, 
      IF_Regsxreg_file_820_port, IF_Regsxreg_file_821_port, 
      IF_Regsxreg_file_822_port, IF_Regsxreg_file_823_port, 
      IF_Regsxreg_file_824_port, IF_Regsxreg_file_825_port, 
      IF_Regsxreg_file_826_port, IF_Regsxreg_file_827_port, 
      IF_Regsxreg_file_828_port, IF_Regsxreg_file_829_port, 
      IF_Regsxreg_file_830_port, IF_Regsxreg_file_831_port, 
      IF_Regsxreg_file_832_port, IF_Regsxreg_file_833_port, 
      IF_Regsxreg_file_834_port, IF_Regsxreg_file_835_port, 
      IF_Regsxreg_file_836_port, IF_Regsxreg_file_837_port, 
      IF_Regsxreg_file_838_port, IF_Regsxreg_file_839_port, 
      IF_Regsxreg_file_840_port, IF_Regsxreg_file_841_port, 
      IF_Regsxreg_file_842_port, IF_Regsxreg_file_843_port, 
      IF_Regsxreg_file_844_port, IF_Regsxreg_file_845_port, 
      IF_Regsxreg_file_846_port, IF_Regsxreg_file_847_port, 
      IF_Regsxreg_file_848_port, IF_Regsxreg_file_849_port, 
      IF_Regsxreg_file_850_port, IF_Regsxreg_file_851_port, 
      IF_Regsxreg_file_852_port, IF_Regsxreg_file_853_port, 
      IF_Regsxreg_file_854_port, IF_Regsxreg_file_855_port, 
      IF_Regsxreg_file_856_port, IF_Regsxreg_file_857_port, 
      IF_Regsxreg_file_858_port, IF_Regsxreg_file_859_port, 
      IF_Regsxreg_file_860_port, IF_Regsxreg_file_861_port, 
      IF_Regsxreg_file_862_port, IF_Regsxreg_file_863_port, 
      IF_Regsxreg_file_864_port, IF_Regsxreg_file_865_port, 
      IF_Regsxreg_file_866_port, IF_Regsxreg_file_867_port, 
      IF_Regsxreg_file_868_port, IF_Regsxreg_file_869_port, 
      IF_Regsxreg_file_870_port, IF_Regsxreg_file_871_port, 
      IF_Regsxreg_file_872_port, IF_Regsxreg_file_873_port, 
      IF_Regsxreg_file_874_port, IF_Regsxreg_file_875_port, 
      IF_Regsxreg_file_876_port, IF_Regsxreg_file_877_port, 
      IF_Regsxreg_file_878_port, IF_Regsxreg_file_879_port, 
      IF_Regsxreg_file_880_port, IF_Regsxreg_file_881_port, 
      IF_Regsxreg_file_882_port, IF_Regsxreg_file_883_port, 
      IF_Regsxreg_file_884_port, IF_Regsxreg_file_885_port, 
      IF_Regsxreg_file_886_port, IF_Regsxreg_file_887_port, 
      IF_Regsxreg_file_888_port, IF_Regsxreg_file_889_port, 
      IF_Regsxreg_file_890_port, IF_Regsxreg_file_891_port, 
      IF_Regsxreg_file_892_port, IF_Regsxreg_file_893_port, 
      IF_Regsxreg_file_894_port, IF_Regsxreg_file_895_port, 
      IF_Regsxreg_file_896_port, IF_Regsxreg_file_897_port, 
      IF_Regsxreg_file_898_port, IF_Regsxreg_file_899_port, 
      IF_Regsxreg_file_900_port, IF_Regsxreg_file_901_port, 
      IF_Regsxreg_file_902_port, IF_Regsxreg_file_903_port, 
      IF_Regsxreg_file_904_port, IF_Regsxreg_file_905_port, 
      IF_Regsxreg_file_906_port, IF_Regsxreg_file_907_port, 
      IF_Regsxreg_file_908_port, IF_Regsxreg_file_909_port, 
      IF_Regsxreg_file_910_port, IF_Regsxreg_file_911_port, 
      IF_Regsxreg_file_912_port, IF_Regsxreg_file_913_port, 
      IF_Regsxreg_file_914_port, IF_Regsxreg_file_915_port, 
      IF_Regsxreg_file_916_port, IF_Regsxreg_file_917_port, 
      IF_Regsxreg_file_918_port, IF_Regsxreg_file_919_port, 
      IF_Regsxreg_file_920_port, IF_Regsxreg_file_921_port, 
      IF_Regsxreg_file_922_port, IF_Regsxreg_file_923_port, 
      IF_Regsxreg_file_924_port, IF_Regsxreg_file_925_port, 
      IF_Regsxreg_file_926_port, IF_Regsxreg_file_927_port, 
      IF_Regsxreg_file_928_port, IF_Regsxreg_file_929_port, 
      IF_Regsxreg_file_930_port, IF_Regsxreg_file_931_port, 
      IF_Regsxreg_file_932_port, IF_Regsxreg_file_933_port, 
      IF_Regsxreg_file_934_port, IF_Regsxreg_file_935_port, 
      IF_Regsxreg_file_936_port, IF_Regsxreg_file_937_port, 
      IF_Regsxreg_file_938_port, IF_Regsxreg_file_939_port, 
      IF_Regsxreg_file_940_port, IF_Regsxreg_file_941_port, 
      IF_Regsxreg_file_942_port, IF_Regsxreg_file_943_port, 
      IF_Regsxreg_file_944_port, IF_Regsxreg_file_945_port, 
      IF_Regsxreg_file_946_port, IF_Regsxreg_file_947_port, 
      IF_Regsxreg_file_948_port, IF_Regsxreg_file_949_port, 
      IF_Regsxreg_file_950_port, IF_Regsxreg_file_951_port, 
      IF_Regsxreg_file_952_port, IF_Regsxreg_file_953_port, 
      IF_Regsxreg_file_954_port, IF_Regsxreg_file_955_port, 
      IF_Regsxreg_file_956_port, IF_Regsxreg_file_957_port, 
      IF_Regsxreg_file_958_port, IF_Regsxreg_file_959_port, 
      IF_Regsxreg_file_960_port, IF_Regsxreg_file_961_port, 
      IF_Regsxreg_file_962_port, IF_Regsxreg_file_963_port, 
      IF_Regsxreg_file_964_port, IF_Regsxreg_file_965_port, 
      IF_Regsxreg_file_966_port, IF_Regsxreg_file_967_port, 
      IF_Regsxreg_file_968_port, IF_Regsxreg_file_969_port, 
      IF_Regsxreg_file_970_port, IF_Regsxreg_file_971_port, 
      IF_Regsxreg_file_972_port, IF_Regsxreg_file_973_port, 
      IF_Regsxreg_file_974_port, IF_Regsxreg_file_975_port, 
      IF_Regsxreg_file_976_port, IF_Regsxreg_file_977_port, 
      IF_Regsxreg_file_978_port, IF_Regsxreg_file_979_port, 
      IF_Regsxreg_file_980_port, IF_Regsxreg_file_981_port, 
      IF_Regsxreg_file_982_port, IF_Regsxreg_file_983_port, 
      IF_Regsxreg_file_984_port, IF_Regsxreg_file_985_port, 
      IF_Regsxreg_file_986_port, IF_Regsxreg_file_987_port, 
      IF_Regsxreg_file_988_port, IF_Regsxreg_file_989_port, 
      IF_Regsxreg_file_990_port, IF_Regsxreg_file_991_port, net2468144, 
      net2468149, net2468154, net2468159, net2468164, net2468169, net2468174, 
      net2468179, net2468184, net2468189, net2468194, net2468199, net2468204, 
      net2468209, net2468214, net2468219, net2468224, net2468229, net2468234, 
      net2468239, net2468249, net2468254, net2468259, net2468264, net2468269, 
      net2468274, net2468279, net2468284, net2468289, net2468294, net2468299, 
      net2468304, net2468309, net2468314, net2468319, net2468324, net2468329, 
      net2468334, net2468339, net2468344, net2468349, net2468354, net2468359, 
      net2468364, net2468369, net2468374, net2468379, net2468384, net2468389, 
      net2468394, net2468399, net2468404, net2468409, net2468414, C596xDATA2_0,
      C596xDATA2_1, C596xDATA2_2, C596xDATA2_3, C596xDATA2_4, C596xDATA2_5, 
      C596xDATA2_6, C596xDATA2_7, C596xDATA2_8, C596xDATA2_9, C596xDATA2_10, 
      C596xDATA2_11, C596xDATA2_12, C596xDATA2_13, C596xDATA2_14, C596xDATA2_15
      , C596xDATA2_16, C596xDATA2_17, C596xDATA2_18, C596xDATA2_19, 
      C596xDATA2_20, C596xDATA2_21, C596xDATA2_22, C596xDATA2_23, C596xDATA2_24
      , C596xDATA2_25, C596xDATA2_26, C596xDATA2_27, C596xDATA2_28, 
      C596xDATA2_29, C596xDATA2_30, n2944, n2946, DP_OP_1698J95_122_4028xn68, 
      DP_OP_1698J95_122_4028xn67, DP_OP_1698J95_122_4028xn66, 
      DP_OP_1698J95_122_4028xn65, DP_OP_1698J95_122_4028xn64, 
      DP_OP_1698J95_122_4028xn63, DP_OP_1698J95_122_4028xn62, 
      DP_OP_1698J95_122_4028xn61, DP_OP_1698J95_122_4028xn60, 
      DP_OP_1698J95_122_4028xn59, DP_OP_1698J95_122_4028xn58, 
      DP_OP_1698J95_122_4028xn57, DP_OP_1698J95_122_4028xn56, 
      DP_OP_1698J95_122_4028xn55, DP_OP_1698J95_122_4028xn54, 
      DP_OP_1698J95_122_4028xn53, DP_OP_1698J95_122_4028xn52, 
      DP_OP_1698J95_122_4028xn51, DP_OP_1698J95_122_4028xn50, 
      DP_OP_1698J95_122_4028xn49, DP_OP_1698J95_122_4028xn48, 
      DP_OP_1698J95_122_4028xn47, DP_OP_1698J95_122_4028xn46, 
      DP_OP_1698J95_122_4028xn45, DP_OP_1698J95_122_4028xn44, 
      DP_OP_1698J95_122_4028xn43, DP_OP_1698J95_122_4028xn42, 
      DP_OP_1698J95_122_4028xn41, DP_OP_1698J95_122_4028xn40, 
      DP_OP_1698J95_122_4028xn39, DP_OP_1698J95_122_4028xn38, 
      DP_OP_1698J95_122_4028xn32, DP_OP_1698J95_122_4028xn31, 
      DP_OP_1698J95_122_4028xn30, DP_OP_1698J95_122_4028xn29, 
      DP_OP_1698J95_122_4028xn28, DP_OP_1698J95_122_4028xn27, 
      DP_OP_1698J95_122_4028xn26, DP_OP_1698J95_122_4028xn25, 
      DP_OP_1698J95_122_4028xn24, DP_OP_1698J95_122_4028xn23, 
      DP_OP_1698J95_122_4028xn22, DP_OP_1698J95_122_4028xn21, 
      DP_OP_1698J95_122_4028xn20, DP_OP_1698J95_122_4028xn19, 
      DP_OP_1698J95_122_4028xn18, DP_OP_1698J95_122_4028xn17, 
      DP_OP_1698J95_122_4028xn16, DP_OP_1698J95_122_4028xn15, 
      DP_OP_1698J95_122_4028xn14, DP_OP_1698J95_122_4028xn13, 
      DP_OP_1698J95_122_4028xn12, DP_OP_1698J95_122_4028xn11, 
      DP_OP_1698J95_122_4028xn10, DP_OP_1698J95_122_4028xn9, 
      DP_OP_1698J95_122_4028xn8, DP_OP_1698J95_122_4028xn7, 
      DP_OP_1698J95_122_4028xn6, DP_OP_1698J95_122_4028xn5, 
      DP_OP_1698J95_122_4028xn4, DP_OP_1698J95_122_4028xn3, 
      DP_OP_1698J95_122_4028xn2, DP_OP_1703J95_125_7309xn131, 
      DP_OP_1703J95_125_7309xn130, DP_OP_1703J95_125_7309xn129, 
      DP_OP_1703J95_125_7309xn128, DP_OP_1703J95_125_7309xn127, 
      DP_OP_1703J95_125_7309xn126, DP_OP_1703J95_125_7309xn125, 
      DP_OP_1703J95_125_7309xn124, DP_OP_1703J95_125_7309xn123, 
      DP_OP_1703J95_125_7309xn122, DP_OP_1703J95_125_7309xn121, 
      DP_OP_1703J95_125_7309xn120, DP_OP_1703J95_125_7309xn119, 
      DP_OP_1703J95_125_7309xn118, DP_OP_1703J95_125_7309xn117, 
      DP_OP_1703J95_125_7309xn116, DP_OP_1703J95_125_7309xn115, 
      DP_OP_1703J95_125_7309xn114, DP_OP_1703J95_125_7309xn113, 
      DP_OP_1703J95_125_7309xn112, DP_OP_1703J95_125_7309xn111, 
      DP_OP_1703J95_125_7309xn110, DP_OP_1703J95_125_7309xn109, 
      DP_OP_1703J95_125_7309xn108, DP_OP_1703J95_125_7309xn107, 
      DP_OP_1703J95_125_7309xn106, DP_OP_1703J95_125_7309xn105, 
      DP_OP_1703J95_125_7309xn104, DP_OP_1703J95_125_7309xn103, 
      DP_OP_1703J95_125_7309xn102, DP_OP_1703J95_125_7309xn101, 
      DP_OP_1703J95_125_7309xn32, DP_OP_1703J95_125_7309xn31, 
      DP_OP_1703J95_125_7309xn30, DP_OP_1703J95_125_7309xn29, 
      DP_OP_1703J95_125_7309xn28, DP_OP_1703J95_125_7309xn27, 
      DP_OP_1703J95_125_7309xn26, DP_OP_1703J95_125_7309xn25, 
      DP_OP_1703J95_125_7309xn24, DP_OP_1703J95_125_7309xn23, 
      DP_OP_1703J95_125_7309xn22, DP_OP_1703J95_125_7309xn21, 
      DP_OP_1703J95_125_7309xn20, DP_OP_1703J95_125_7309xn19, 
      DP_OP_1703J95_125_7309xn18, DP_OP_1703J95_125_7309xn17, 
      DP_OP_1703J95_125_7309xn16, DP_OP_1703J95_125_7309xn15, 
      DP_OP_1703J95_125_7309xn14, DP_OP_1703J95_125_7309xn13, 
      DP_OP_1703J95_125_7309xn12, DP_OP_1703J95_125_7309xn11, 
      DP_OP_1703J95_125_7309xn10, DP_OP_1703J95_125_7309xn9, 
      DP_OP_1703J95_125_7309xn8, DP_OP_1703J95_125_7309xn7, 
      DP_OP_1703J95_125_7309xn6, DP_OP_1703J95_125_7309xn5, 
      DP_OP_1703J95_125_7309xn4, DP_OP_1703J95_125_7309xn3, 
      DP_OP_1703J95_125_7309xn2, n2952, n2953, n2954, n2955, n2956, n2957, 
      n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, 
      n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, 
      n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, 
      n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, 
      n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, 
      n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, 
      n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, 
      n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, 
      n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, 
      n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, 
      n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, 
      n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, 
      n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, 
      n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, 
      n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, 
      n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, 
      n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, 
      n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, 
      n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, 
      n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, 
      n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, 
      n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, 
      n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, 
      n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, 
      n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, 
      n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, 
      n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, 
      n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, 
      n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, 
      n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, 
      n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, 
      n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, 
      n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, 
      n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, 
      n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, 
      n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, 
      n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, 
      n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, 
      n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, 
      n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, 
      n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, 
      n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, 
      n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, 
      n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, 
      n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, 
      n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, 
      n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, 
      n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, 
      n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, 
      n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, 
      n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, 
      n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, 
      n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, 
      n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, 
      n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, 
      n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, 
      n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, 
      n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, 
      n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, 
      n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, 
      n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, 
      n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, 
      n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, 
      n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, 
      n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, 
      n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, 
      n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, 
      n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, 
      n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, 
      n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, 
      n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, 
      n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, 
      n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, 
      n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, 
      n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, 
      n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, 
      n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, 
      n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, 
      n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, 
      n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, 
      n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, 
      n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, 
      n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, 
      n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, 
      n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, 
      n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, 
      n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, 
      n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, 
      n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, 
      n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, 
      n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, 
      n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, 
      n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, 
      n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, 
      n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, 
      n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, 
      n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, 
      n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, 
      n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, 
      n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, 
      n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, 
      n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, 
      n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, 
      n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, 
      n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, 
      n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, 
      n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, 
      n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, 
      n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, 
      n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, 
      n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, 
      n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, 
      n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, 
      n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, 
      n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, 
      n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, 
      n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, 
      n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, 
      n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, 
      n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, 
      n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, 
      n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, 
      n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, 
      n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
      n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, 
      n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, 
      n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, 
      n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, 
      n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, 
      n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, 
      n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, 
      n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, 
      n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, 
      n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, 
      n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, 
      n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, 
      n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, 
      n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, 
      n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, 
      n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, 
      n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, 
      n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, 
      n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, 
      n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, 
      n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, 
      n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, 
      n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, 
      n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, 
      n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, 
      n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, 
      n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, 
      n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, 
      n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, 
      n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, 
      n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, 
      n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, 
      n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, 
      n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, 
      n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, 
      n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, 
      n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, 
      n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, 
      n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, 
      n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, 
      n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, 
      n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, 
      n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, 
      n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, 
      n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, 
      n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, 
      n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, 
      n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, 
      n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, 
      n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, 
      n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, 
      n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, 
      n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, 
      n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, 
      n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, 
      n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, 
      n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, 
      n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, 
      n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, 
      n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, 
      n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, 
      n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, 
      n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, 
      n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, 
      n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, 
      n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, 
      n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, 
      n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, 
      n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, 
      n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, 
      n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, 
      n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, 
      n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, 
      n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, 
      n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, 
      n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, 
      n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, 
      n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, 
      n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, 
      n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, 
      n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, 
      n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, 
      n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, 
      n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, 
      n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, 
      n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, 
      n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, 
      n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, 
      n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, 
      n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, 
      n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, 
      n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, 
      n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, 
      n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, 
      n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, 
      n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, 
      n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, 
      n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, 
      n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, 
      n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, 
      n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, 
      n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, 
      n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, 
      n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, 
      n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, 
      n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, 
      n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, 
      n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, 
      n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, 
      n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, 
      n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, 
      n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, 
      n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, 
      n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, 
      n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, 
      n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, 
      n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, 
      n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, 
      n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, 
      n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, 
      n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, 
      n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, 
      n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, 
      n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, 
      n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, 
      n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, 
      n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, 
      n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, 
      n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, 
      n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, 
      n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, 
      n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, 
      n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, 
      n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, 
      n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, 
      n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, 
      n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, 
      n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, 
      n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, 
      n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, 
      n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, 
      n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, 
      n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, 
      n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, 
      n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, 
      n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, 
      n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, 
      n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, 
      n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, 
      n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, 
      n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, 
      n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, 
      n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, 
      n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, 
      n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, 
      n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, 
      n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, 
      n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, 
      n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, 
      n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, 
      n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, 
      n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, 
      n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, 
      n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, 
      n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, 
      n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, 
      n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, 
      n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, 
      n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, 
      n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, 
      n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, 
      n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, 
      n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, 
      n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, 
      n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, 
      n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, 
      n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, 
      n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, 
      n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, 
      n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, 
      n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, 
      n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, 
      n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, 
      n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, 
      n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, 
      n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, 
      n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, 
      n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, 
      n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, 
      n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, 
      n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, 
      n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, 
      n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, 
      n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, 
      n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, 
      n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, 
      n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, 
      n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, 
      n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, 
      n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, 
      n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, 
      n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, 
      n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, 
      n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, 
      n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, 
      n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, 
      n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, 
      n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, 
      n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, 
      n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, 
      n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, 
      n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, 
      n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, 
      n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, 
      n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, 
      n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, 
      n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, 
      n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, 
      n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, 
      n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, 
      n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, 
      n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, 
      n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, 
      n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, 
      n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, 
      n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, 
      n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, 
      n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, 
      n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, 
      n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, 
      n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, 
      n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, 
      n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, 
      n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, 
      n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, 
      n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, 
      n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, 
      n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, 
      n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, 
      n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, 
      n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, 
      n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, 
      n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, 
      n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, 
      n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, 
      n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, 
      n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, 
      n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, 
      n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, 
      n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, 
      n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, 
      n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, 
      n6718, n6719, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, 
      n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, 
      n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, 
      n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, 
      n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, 
      n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, 
      n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, 
      n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, 
      n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, 
      n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, 
      n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, 
      n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, 
      n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, 
      n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, 
      n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, 
      n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, 
      n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, 
      n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, 
      n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, 
      n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, 
      n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, 
      n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, 
      n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, 
      n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, 
      n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, 
      n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, 
      n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, 
      n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, 
      n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, 
      n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, 
      n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, 
      n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, 
      n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, 
      n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, 
      n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, 
      n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, 
      n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, 
      n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, 
      n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, 
      n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, 
      n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, 
      n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, 
      n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, 
      n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, 
      n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, 
      n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, 
      n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, 
      n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, 
      n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, 
      n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, 
      n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, 
      n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, 
      n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, 
      n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, 
      n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, 
      n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, 
      n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, 
      n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, 
      n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, 
      n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, 
      n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, 
      n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, 
      n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, 
      n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, 
      n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, 
      n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, 
      n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, 
      n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, 
      n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, 
      n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, 
      n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, 
      n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, 
      n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, 
      n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, 
      n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, 
      n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, 
      n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, 
      n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, 
      n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, 
      n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, 
      n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, 
      n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, 
      n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, 
      n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, 
      n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, 
      n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, 
      n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, 
      n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, 
      n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, 
      n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, 
      n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, 
      n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, 
      n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, 
      n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, 
      n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, 
      n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, 
      n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, 
      n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, 
      n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, 
      n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, 
      n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, 
      n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, 
      n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, 
      n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, 
      n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, 
      n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, 
      n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, 
      n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, 
      n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, 
      n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, 
      n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, 
      n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, 
      n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, 
      n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, 
      n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, 
      n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, 
      n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, 
      n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, 
      n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, 
      n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, 
      n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, 
      n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, 
      n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, 
      n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, 
      n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, 
      n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, 
      n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, 
      n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, 
      n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, 
      n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, 
      n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, 
      n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, 
      n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, 
      n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, 
      n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, 
      n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, 
      n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, 
      n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, 
      n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, 
      n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, 
      n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, 
      n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, 
      n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, 
      n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, 
      n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, 
      n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, 
      n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, 
      n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, 
      n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, 
      n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, 
      n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, 
      n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, 
      n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, 
      n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, 
      n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, 
      n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, 
      n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, 
      n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, 
      n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, 
      n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, 
      n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, 
      n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, 
      n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, 
      n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, 
      n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, 
      n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, 
      n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, 
      n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, 
      n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, 
      n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, 
      n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, 
      n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, 
      n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, 
      n_2555, n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, 
      n_2564, n_2565, n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, 
      n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, n_2579 : std_logic;

begin
   MemToCtl_port_notify <= MemToCtl_port_notify_port;
   CtlToMem_port_notify <= CtlToMem_port_notify_port;
   
   IF_DecoderxDecToCtl_port_encType_regx2x : DFF_X1 port map( D => 
                           IF_DecoderxN551, CK => net2468249, Q => 
                           DecToCtl_port_encType_2_port, QN => n6230);
   IF_CPathxsection_regx1x : DFF_X1 port map( D => IF_CPathxN1856, CK => 
                           net2468239, Q => n6207, QN => n6227);
   IF_CPathxCtlToDec_port_notify_reg : DFF_X1 port map( D => n2946, CK => 
                           net2468239, Q => CtlToDec_port_notify, QN => n_1000)
                           ;
   IF_CPathxmem_en_signal_reg : DFF_X1 port map( D => n6505, CK => net2468169, 
                           Q => IF_CPathxmem_en_signal, QN => n6199);
   IF_CPathxsection_regx3x : DFF_X1 port map( D => IF_CPathxN1858, CK => 
                           net2468239, Q => IF_CPathxsection_3_port, QN => 
                           n6228);
   IF_CPathxsection_regx0x : DFF_X1 port map( D => n6687, CK => net2468239, Q 
                           => IF_CPathxsection_0_port, QN => n_1001);
   IF_CPathxCtlToDec_port_regx0x : DFF_X1 port map( D => MemToCtl_port(0), CK 
                           => net2468159, Q => CtlToDec_port_0_port, QN => 
                           n_1002);
   IF_CPathxCtlToDec_port_regx1x : DFF_X1 port map( D => MemToCtl_port(1), CK 
                           => net2468159, Q => CtlToDec_port_1_port, QN => 
                           n_1003);
   IF_CPathxCtlToDec_port_regx2x : DFF_X1 port map( D => MemToCtl_port(2), CK 
                           => net2468159, Q => CtlToDec_port_2_port, QN => 
                           n6229);
   IF_CPathxCtlToDec_port_regx3x : DFF_X1 port map( D => MemToCtl_port(3), CK 
                           => net2468159, Q => CtlToDec_port_3_port, QN => 
                           n6231);
   IF_CPathxCtlToDec_port_regx4x : DFF_X1 port map( D => MemToCtl_port(4), CK 
                           => net2468159, Q => CtlToDec_port_4_port, QN => 
                           n6234);
   IF_CPathxCtlToDec_port_regx5x : DFF_X1 port map( D => MemToCtl_port(5), CK 
                           => net2468159, Q => CtlToDec_port_5_port, QN => 
                           n_1004);
   IF_CPathxCtlToDec_port_regx6x : DFF_X1 port map( D => MemToCtl_port(6), CK 
                           => net2468159, Q => CtlToDec_port_6_port, QN => 
                           n_1005);
   IF_DecoderxDecToCtl_port_encType_regx0x : DFF_X1 port map( D => 
                           IF_DecoderxN549, CK => net2468249, Q => 
                           DecToCtl_port_encType_0_port, QN => n6197);
   IF_CPathxCtlToDec_port_regx7x : DFF_X1 port map( D => MemToCtl_port(7), CK 
                           => net2468159, Q => CtlToDec_port_7_port, QN => 
                           n_1006);
   IF_DecoderxDecToCtl_port_rd_addr_regx0x : DFF_X1 port map( D => 
                           IF_DecoderxN591, CK => net2468249, Q => 
                           DecToCtl_port_rd_addr_0_port, QN => n_1007);
   IF_CPathxCtlToDec_port_regx8x : DFF_X1 port map( D => MemToCtl_port(8), CK 
                           => net2468159, Q => n_1008, QN => n6319);
   IF_DecoderxDecToCtl_port_rd_addr_regx1x : DFF_X1 port map( D => 
                           IF_DecoderxN592, CK => net2468249, Q => 
                           DecToCtl_port_rd_addr_1_port, QN => n_1009);
   IF_CPathxCtlToDec_port_regx9x : DFF_X1 port map( D => MemToCtl_port(9), CK 
                           => net2468159, Q => n_1010, QN => n6320);
   IF_DecoderxDecToCtl_port_rd_addr_regx2x : DFF_X1 port map( D => 
                           IF_DecoderxN593, CK => net2468249, Q => 
                           DecToCtl_port_rd_addr_2_port, QN => n_1011);
   IF_CPathxCtlToDec_port_regx10x : DFF_X1 port map( D => MemToCtl_port(10), CK
                           => net2468159, Q => n_1012, QN => n6321);
   IF_DecoderxDecToCtl_port_rd_addr_regx3x : DFF_X1 port map( D => 
                           IF_DecoderxN594, CK => net2468249, Q => 
                           DecToCtl_port_rd_addr_3_port, QN => n_1013);
   IF_CPathxCtlToDec_port_regx11x : DFF_X1 port map( D => MemToCtl_port(11), CK
                           => net2468159, Q => n_1014, QN => n6322);
   IF_DecoderxDecToCtl_port_rd_addr_regx4x : DFF_X1 port map( D => 
                           IF_DecoderxN595, CK => net2468249, Q => 
                           DecToCtl_port_rd_addr_4_port, QN => n_1015);
   IF_CPathxCtlToDec_port_regx12x : DFF_X1 port map( D => MemToCtl_port(12), CK
                           => net2468159, Q => CtlToDec_port_12_port, QN => 
                           n6259);
   IF_CPathxCtlToDec_port_regx13x : DFF_X1 port map( D => MemToCtl_port(13), CK
                           => net2468159, Q => CtlToDec_port_13_port, QN => 
                           n6208);
   IF_CPathxCtlToDec_port_regx14x : DFF_X1 port map( D => MemToCtl_port(14), CK
                           => net2468159, Q => CtlToDec_port_14_port, QN => 
                           n6261);
   IF_CPathxCtlToDec_port_regx15x : DFF_X1 port map( D => MemToCtl_port(15), CK
                           => net2468159, Q => n_1016, QN => n6324);
   IF_DecoderxDecToCtl_port_rs1_addr_regx0x : DFF_X1 port map( D => 
                           IF_DecoderxN597, CK => net2468249, Q => 
                           DecToCtl_port_rs1_addr_0_port, QN => n_1017);
   IF_CPathxCtlToDec_port_regx16x : DFF_X1 port map( D => MemToCtl_port(16), CK
                           => net2468159, Q => n_1018, QN => n6325);
   IF_DecoderxDecToCtl_port_rs1_addr_regx1x : DFF_X1 port map( D => 
                           IF_DecoderxN598, CK => net2468249, Q => 
                           DecToCtl_port_rs1_addr_1_port, QN => n_1019);
   IF_CPathxCtlToDec_port_regx17x : DFF_X1 port map( D => MemToCtl_port(17), CK
                           => net2468159, Q => n_1020, QN => n6326);
   IF_DecoderxDecToCtl_port_rs1_addr_regx2x : DFF_X1 port map( D => 
                           IF_DecoderxN599, CK => net2468249, Q => 
                           DecToCtl_port_rs1_addr_2_port, QN => n_1021);
   IF_CPathxCtlToDec_port_regx18x : DFF_X1 port map( D => MemToCtl_port(18), CK
                           => net2468159, Q => n_1022, QN => n6327);
   IF_DecoderxDecToCtl_port_rs1_addr_regx3x : DFF_X1 port map( D => 
                           IF_DecoderxN600, CK => net2468249, Q => 
                           DecToCtl_port_rs1_addr_3_port, QN => n_1023);
   IF_CPathxCtlToDec_port_regx19x : DFF_X1 port map( D => MemToCtl_port(19), CK
                           => net2468159, Q => n_1024, QN => n6328);
   IF_DecoderxDecToCtl_port_rs1_addr_regx4x : DFF_X1 port map( D => 
                           IF_DecoderxN601, CK => net2468249, Q => 
                           DecToCtl_port_rs1_addr_4_port, QN => n_1025);
   IF_CPathxCtlToDec_port_regx20x : DFF_X1 port map( D => MemToCtl_port(20), CK
                           => net2468159, Q => CtlToDec_port_20_port, QN => 
                           n6274);
   IF_DecoderxDecToCtl_port_rs2_addr_regx0x : DFF_X1 port map( D => 
                           IF_DecoderxN602, CK => net2468249, Q => 
                           DecToCtl_port_rs2_addr_0_port, QN => n_1026);
   IF_CPathxCtlToDec_port_regx21x : DFF_X1 port map( D => MemToCtl_port(21), CK
                           => net2468159, Q => n_1027, QN => n6210);
   IF_DecoderxDecToCtl_port_rs2_addr_regx1x : DFF_X1 port map( D => 
                           IF_DecoderxN603, CK => net2468249, Q => 
                           DecToCtl_port_rs2_addr_1_port, QN => n_1028);
   IF_CPathxCtlToDec_port_regx22x : DFF_X1 port map( D => MemToCtl_port(22), CK
                           => net2468159, Q => n_1029, QN => n6211);
   IF_DecoderxDecToCtl_port_rs2_addr_regx2x : DFF_X1 port map( D => 
                           IF_DecoderxN604, CK => net2468249, Q => 
                           DecToCtl_port_rs2_addr_2_port, QN => n_1030);
   IF_CPathxCtlToDec_port_regx23x : DFF_X1 port map( D => MemToCtl_port(23), CK
                           => net2468159, Q => n_1031, QN => n6212);
   IF_DecoderxDecToCtl_port_rs2_addr_regx3x : DFF_X1 port map( D => 
                           IF_DecoderxN605, CK => net2468249, Q => 
                           DecToCtl_port_rs2_addr_3_port, QN => n_1032);
   IF_CPathxCtlToDec_port_regx24x : DFF_X1 port map( D => MemToCtl_port(24), CK
                           => net2468159, Q => n_1033, QN => n6213);
   IF_DecoderxDecToCtl_port_rs2_addr_regx4x : DFF_X1 port map( D => 
                           IF_DecoderxN606, CK => net2468249, Q => 
                           DecToCtl_port_rs2_addr_4_port, QN => n_1034);
   IF_CPathxCtlToDec_port_regx25x : DFF_X1 port map( D => MemToCtl_port(25), CK
                           => net2468159, Q => n_1035, QN => n6264);
   IF_CPathxCtlToDec_port_regx26x : DFF_X1 port map( D => MemToCtl_port(26), CK
                           => net2468159, Q => CtlToDec_port_26_port, QN => 
                           n6273);
   IF_CPathxCtlToDec_port_regx27x : DFF_X1 port map( D => MemToCtl_port(27), CK
                           => net2468159, Q => CtlToDec_port_27_port, QN => 
                           n6271);
   IF_CPathxCtlToDec_port_regx28x : DFF_X1 port map( D => MemToCtl_port(28), CK
                           => net2468159, Q => CtlToDec_port_28_port, QN => 
                           n6272);
   IF_CPathxCtlToDec_port_regx29x : DFF_X1 port map( D => MemToCtl_port(29), CK
                           => net2468159, Q => CtlToDec_port_29_port, QN => 
                           n6270);
   IF_CPathxCtlToDec_port_regx30x : DFF_X1 port map( D => MemToCtl_port(30), CK
                           => net2468159, Q => CtlToDec_port_30_port, QN => 
                           n6260);
   IF_CPathxCtlToDec_port_regx31x : DFF_X1 port map( D => MemToCtl_port(31), CK
                           => net2468159, Q => CtlToDec_port_31_port, QN => 
                           n6209);
   IF_DecoderxDecToCtl_port_instrType_regx1x : DFF_X1 port map( D => 
                           IF_DecoderxN586, CK => net2468249, Q => 
                           DecToCtl_port_instrType_1_port, QN => n2953);
   IF_DecoderxDecToCtl_port_instrType_regx3x : DFF_X1 port map( D => 
                           IF_DecoderxN588, CK => net2468249, Q => 
                           DecToCtl_port_instrType_3_port, QN => n6189);
   IF_DecoderxDecToCtl_port_instrType_regx5x : DFF_X1 port map( D => 
                           IF_DecoderxN590, CK => net2468249, Q => 
                           DecToCtl_port_instrType_5_port, QN => n6226);
   IF_DecoderxDecToCtl_port_instrType_regx0x : DFF_X1 port map( D => 
                           IF_DecoderxN585, CK => net2468249, Q => 
                           DecToCtl_port_instrType_0_port, QN => n6232);
   IF_CPathxsection_regx2x : DFF_X1 port map( D => n6686, CK => net2468239, Q 
                           => IF_CPathxsection_2_port, QN => n6196);
   IF_CPathxDecToCtl_data_signal_rd_addr_regx0x : DFF_X1 port map( D => 
                           IF_CPathxN2196, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_rd_addr_0_port, QN => 
                           n6236);
   IF_CPathxDecToCtl_data_signal_rd_addr_regx1x : DFF_X1 port map( D => 
                           IF_CPathxN2197, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_rd_addr_1_port, QN => 
                           n6200);
   IF_CPathxDecToCtl_data_signal_rd_addr_regx2x : DFF_X1 port map( D => 
                           IF_CPathxN2198, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_rd_addr_2_port, QN => 
                           n6192);
   IF_CPathxDecToCtl_data_signal_rd_addr_regx3x : DFF_X1 port map( D => 
                           IF_CPathxN2199, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_rd_addr_3_port, QN => 
                           n6190);
   IF_CPathxDecToCtl_data_signal_rd_addr_regx4x : DFF_X1 port map( D => 
                           IF_CPathxN2200, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_rd_addr_4_port, QN => 
                           n_1036);
   IF_CPathxDecToCtl_data_signal_instrType_regx0x : DFF_X1 port map( D => 
                           IF_CPathxN2190, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_instrType_0_port, QN 
                           => n_1037);
   IF_CPathxDecToCtl_data_signal_instrType_regx1x : DFF_X1 port map( D => 
                           IF_CPathxN2191, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_instrType_1_port, QN 
                           => n6240);
   IF_CPathxDecToCtl_data_signal_instrType_regx2x : DFF_X1 port map( D => 
                           IF_CPathxN2192, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_instrType_2_port, QN 
                           => n_1038);
   IF_CPathxDecToCtl_data_signal_instrType_regx3x : DFF_X1 port map( D => 
                           IF_CPathxN2193, CK => net2468194, Q => n_1039, QN =>
                           n6239);
   IF_CPathxDecToCtl_data_signal_instrType_regx4x : DFF_X1 port map( D => 
                           IF_CPathxN2194, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_instrType_4_port, QN 
                           => n_1040);
   IF_CPathxDecToCtl_data_signal_instrType_regx5x : DFF_X1 port map( D => 
                           IF_CPathxN2195, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_instrType_5_port, QN 
                           => n_1041);
   IF_CPathxCtlToRegs_data_signal_src2_regx0x : DFF_X1 port map( D => 
                           IF_CPathxN2084, CK => net2468204, Q => 
                           IF_CPathxCtlToRegs_data_signal_src2_0_port, QN => 
                           n_1042);
   IF_CPathxCtlToRegs_data_signal_src2_regx1x : DFF_X1 port map( D => 
                           IF_CPathxN2085, CK => net2468204, Q => 
                           IF_CPathxCtlToRegs_data_signal_src2_1_port, QN => 
                           n_1043);
   IF_CPathxCtlToRegs_data_signal_src2_regx2x : DFF_X1 port map( D => 
                           IF_CPathxN2086, CK => net2468204, Q => 
                           IF_CPathxCtlToRegs_data_signal_src2_2_port, QN => 
                           n_1044);
   IF_CPathxCtlToRegs_data_signal_src2_regx3x : DFF_X1 port map( D => 
                           IF_CPathxN2087, CK => net2468204, Q => 
                           IF_CPathxCtlToRegs_data_signal_src2_3_port, QN => 
                           n_1045);
   IF_CPathxCtlToRegs_data_signal_src2_regx4x : DFF_X1 port map( D => 
                           IF_CPathxN2088, CK => net2468204, Q => 
                           IF_CPathxCtlToRegs_data_signal_src2_4_port, QN => 
                           n_1046);
   IF_CPathxCtlToRegs_data_signal_src1_regx0x : DFF_X1 port map( D => 
                           IF_CPathxN2079, CK => net2468204, Q => 
                           IF_CPathxCtlToRegs_data_signal_src1_0_port, QN => 
                           n_1047);
   IF_CPathxCtlToRegs_data_signal_src1_regx1x : DFF_X1 port map( D => 
                           IF_CPathxN2080, CK => net2468204, Q => 
                           IF_CPathxCtlToRegs_data_signal_src1_1_port, QN => 
                           n_1048);
   IF_CPathxCtlToRegs_data_signal_src1_regx2x : DFF_X1 port map( D => 
                           IF_CPathxN2081, CK => net2468204, Q => 
                           IF_CPathxCtlToRegs_data_signal_src1_2_port, QN => 
                           n_1049);
   IF_CPathxCtlToRegs_data_signal_src1_regx3x : DFF_X1 port map( D => 
                           IF_CPathxN2082, CK => net2468204, Q => 
                           IF_CPathxCtlToRegs_data_signal_src1_3_port, QN => 
                           n_1050);
   IF_CPathxCtlToRegs_data_signal_src1_regx4x : DFF_X1 port map( D => 
                           IF_CPathxN2083, CK => net2468204, Q => 
                           IF_CPathxCtlToRegs_data_signal_src1_4_port, QN => 
                           n_1051);
   IF_CPathxwb_sel_signal_regx0x : DFF_X1 port map( D => n6504, CK => 
                           net2468169, Q => IF_CPathxwb_sel_signal_0_port, QN 
                           => n6269);
   IF_CPathxwb_sel_signal_regx1x : DFF_X1 port map( D => n6503, CK => 
                           net2468169, Q => IF_CPathxwb_sel_signal_1_port, QN 
                           => n_1052);
   IF_CPathxwb_en_signal_reg : DFF_X1 port map( D => IF_CPathxN2309, CK => 
                           net2468169, Q => IF_CPathxwb_en_signal, QN => n_1053
                           );
   IF_CPathxreg_rd_en_signal_reg : DFF_X1 port map( D => IF_CPathxN2308, CK => 
                           net2468169, Q => IF_CPathxreg_rd_en_signal, QN => 
                           n_1054);
   IF_CPathxbr_en_signal_reg : DFF_X1 port map( D => n6502, CK => net2468169, Q
                           => IF_CPathxbr_en_signal, QN => n_1055);
   IF_CPathxCtlToALU_data_signal_op2_sel_regx0x : DFF_X1 port map( D => n6677, 
                           CK => net2468229, Q => 
                           IF_CPathxCtlToALU_data_signal_op2_sel_0_port, QN => 
                           n_1056);
   IF_CPathxCtlToALU_port_op2_sel_regx0x : DFF_X1 port map( D => IF_CPathxN1667
                           , CK => net2468149, Q => 
                           CtlToALU_port_op2_sel_0_port, QN => n6241);
   IF_CPathxCtlToALU_data_signal_op2_sel_regx1x : DFF_X1 port map( D => n6676, 
                           CK => net2468229, Q => 
                           IF_CPathxCtlToALU_data_signal_op2_sel_1_port, QN => 
                           n_1057);
   IF_CPathxCtlToALU_port_op2_sel_regx1x : DFF_X1 port map( D => IF_CPathxN1668
                           , CK => net2468149, Q => 
                           CtlToALU_port_op2_sel_1_port, QN => n6202);
   IF_CPathxCtlToALU_data_signal_op1_sel_regx0x : DFF_X1 port map( D => n6675, 
                           CK => net2468229, Q => 
                           IF_CPathxCtlToALU_data_signal_op1_sel_0_port, QN => 
                           n6345);
   IF_CPathxCtlToALU_port_op1_sel_regx0x : DFF_X1 port map( D => IF_CPathxN1664
                           , CK => net2468149, Q => 
                           CtlToALU_port_op1_sel_0_port, QN => n6242);
   IF_CPathxCtlToALU_data_signal_op1_sel_regx1x : DFF_X1 port map( D => 
                           IF_CPathxN1932, CK => net2468229, Q => 
                           IF_CPathxCtlToALU_data_signal_op1_sel_1_port, QN => 
                           n_1058);
   IF_CPathxCtlToALU_port_op1_sel_regx1x : DFF_X1 port map( D => IF_CPathxN1665
                           , CK => net2468149, Q => 
                           CtlToALU_port_op1_sel_1_port, QN => n6203);
   IF_CPathxCtlToALU_data_signal_alu_fun_regx0x : DFF_X1 port map( D => n6681, 
                           CK => net2468234, Q => 
                           IF_CPathxCtlToALU_data_signal_alu_fun_0_port, QN => 
                           n_1059);
   IF_CPathxCtlToALU_data_signal_alu_fun_regx1x : DFF_X1 port map( D => n6680, 
                           CK => net2468234, Q => 
                           IF_CPathxCtlToALU_data_signal_alu_fun_1_port, QN => 
                           n_1060);
   IF_CPathxCtlToALU_port_alu_fun_regx1x : DFF_X1 port map( D => IF_CPathxN1629
                           , CK => net2468149, Q => 
                           CtlToALU_port_alu_fun_1_port, QN => n6246);
   IF_CPathxCtlToALU_data_signal_alu_fun_regx2x : DFF_X1 port map( D => n6679, 
                           CK => net2468234, Q => 
                           IF_CPathxCtlToALU_data_signal_alu_fun_2_port, QN => 
                           n_1061);
   IF_CPathxCtlToALU_port_alu_fun_regx2x : DFF_X1 port map( D => IF_CPathxN1630
                           , CK => net2468149, Q => 
                           CtlToALU_port_alu_fun_2_port, QN => n6268);
   IF_CPathxCtlToALU_data_signal_alu_fun_regx3x : DFF_X1 port map( D => n6678, 
                           CK => net2468234, Q => 
                           IF_CPathxCtlToALU_data_signal_alu_fun_3_port, QN => 
                           n_1062);
   IF_CPathxCtlToALU_port_alu_fun_regx3x : DFF_X1 port map( D => IF_CPathxN1631
                           , CK => net2468149, Q => 
                           CtlToALU_port_alu_fun_3_port, QN => n6193);
   IF_CPathxmemoryAccess_signal_mask_regx0x : DFF_X1 port map( D => n6540, CK 
                           => net2468184, Q => 
                           IF_CPathxmemoryAccess_signal_mask_0_port, QN => 
                           n_1063);
   IF_CPathxmemoryAccess_signal_mask_regx1x : DFF_X1 port map( D => n6539, CK 
                           => net2468184, Q => 
                           IF_CPathxmemoryAccess_signal_mask_1_port, QN => 
                           n_1064);
   IF_CPathxmemoryAccess_signal_mask_regx2x : DFF_X1 port map( D => n6538, CK 
                           => net2468184, Q => 
                           IF_CPathxmemoryAccess_signal_mask_2_port, QN => 
                           n_1065);
   IF_CPathxMemToCtl_data_signal_regx0x : DFF_X1 port map( D => IF_CPathxN2202,
                           CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_0_port, QN => n_1066);
   IF_CPathxMemToCtl_data_signal_regx1x : DFF_X1 port map( D => IF_CPathxN2203,
                           CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_1_port, QN => n_1067);
   IF_CPathxMemToCtl_data_signal_regx2x : DFF_X1 port map( D => IF_CPathxN2204,
                           CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_2_port, QN => n_1068);
   IF_CPathxMemToCtl_data_signal_regx3x : DFF_X1 port map( D => IF_CPathxN2205,
                           CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_3_port, QN => n_1069);
   IF_CPathxMemToCtl_data_signal_regx4x : DFF_X1 port map( D => IF_CPathxN2206,
                           CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_4_port, QN => n_1070);
   IF_CPathxMemToCtl_data_signal_regx5x : DFF_X1 port map( D => IF_CPathxN2207,
                           CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_5_port, QN => n_1071);
   IF_CPathxMemToCtl_data_signal_regx6x : DFF_X1 port map( D => IF_CPathxN2208,
                           CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_6_port, QN => n_1072);
   IF_CPathxMemToCtl_data_signal_regx7x : DFF_X1 port map( D => IF_CPathxN2209,
                           CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_7_port, QN => n_1073);
   IF_CPathxMemToCtl_data_signal_regx8x : DFF_X1 port map( D => IF_CPathxN2210,
                           CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_8_port, QN => n_1074);
   IF_CPathxMemToCtl_data_signal_regx9x : DFF_X1 port map( D => IF_CPathxN2211,
                           CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_9_port, QN => n_1075);
   IF_CPathxMemToCtl_data_signal_regx10x : DFF_X1 port map( D => IF_CPathxN2212
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_10_port, QN => n_1076)
                           ;
   IF_CPathxMemToCtl_data_signal_regx11x : DFF_X1 port map( D => IF_CPathxN2213
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_11_port, QN => n_1077)
                           ;
   IF_CPathxMemToCtl_data_signal_regx12x : DFF_X1 port map( D => IF_CPathxN2214
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_12_port, QN => n_1078)
                           ;
   IF_CPathxMemToCtl_data_signal_regx13x : DFF_X1 port map( D => IF_CPathxN2215
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_13_port, QN => n_1079)
                           ;
   IF_CPathxMemToCtl_data_signal_regx14x : DFF_X1 port map( D => IF_CPathxN2216
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_14_port, QN => n_1080)
                           ;
   IF_CPathxMemToCtl_data_signal_regx15x : DFF_X1 port map( D => IF_CPathxN2217
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_15_port, QN => n_1081)
                           ;
   IF_CPathxMemToCtl_data_signal_regx16x : DFF_X1 port map( D => IF_CPathxN2218
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_16_port, QN => n_1082)
                           ;
   IF_CPathxMemToCtl_data_signal_regx17x : DFF_X1 port map( D => IF_CPathxN2219
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_17_port, QN => n_1083)
                           ;
   IF_CPathxMemToCtl_data_signal_regx18x : DFF_X1 port map( D => IF_CPathxN2220
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_18_port, QN => n_1084)
                           ;
   IF_CPathxMemToCtl_data_signal_regx19x : DFF_X1 port map( D => IF_CPathxN2221
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_19_port, QN => n_1085)
                           ;
   IF_CPathxMemToCtl_data_signal_regx20x : DFF_X1 port map( D => IF_CPathxN2222
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_20_port, QN => n_1086)
                           ;
   IF_CPathxMemToCtl_data_signal_regx21x : DFF_X1 port map( D => IF_CPathxN2223
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_21_port, QN => n_1087)
                           ;
   IF_CPathxMemToCtl_data_signal_regx22x : DFF_X1 port map( D => IF_CPathxN2224
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_22_port, QN => n_1088)
                           ;
   IF_CPathxMemToCtl_data_signal_regx23x : DFF_X1 port map( D => IF_CPathxN2225
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_23_port, QN => n_1089)
                           ;
   IF_CPathxMemToCtl_data_signal_regx24x : DFF_X1 port map( D => IF_CPathxN2226
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_24_port, QN => n_1090)
                           ;
   IF_CPathxMemToCtl_data_signal_regx25x : DFF_X1 port map( D => IF_CPathxN2227
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_25_port, QN => n_1091)
                           ;
   IF_CPathxMemToCtl_data_signal_regx26x : DFF_X1 port map( D => IF_CPathxN2228
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_26_port, QN => n_1092)
                           ;
   IF_CPathxMemToCtl_data_signal_regx27x : DFF_X1 port map( D => IF_CPathxN2229
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_27_port, QN => n_1093)
                           ;
   IF_CPathxMemToCtl_data_signal_regx28x : DFF_X1 port map( D => IF_CPathxN2230
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_28_port, QN => n_1094)
                           ;
   IF_CPathxMemToCtl_data_signal_regx29x : DFF_X1 port map( D => IF_CPathxN2231
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_29_port, QN => n_1095)
                           ;
   IF_CPathxMemToCtl_data_signal_regx30x : DFF_X1 port map( D => IF_CPathxN2232
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_30_port, QN => n_1096)
                           ;
   IF_CPathxMemToCtl_data_signal_regx31x : DFF_X1 port map( D => IF_CPathxN2233
                           , CK => net2468189, Q => 
                           IF_CPathxMemToCtl_data_signal_31_port, QN => n_1097)
                           ;
   IF_CPathxCtlToRegs_port_src2_regx0x : DFF_X1 port map( D => n6433, CK => 
                           net2468154, Q => CtlToRegs_port_src2_0_port, QN => 
                           n6266);
   IF_CPathxCtlToRegs_port_src2_regx1x : DFF_X1 port map( D => n6432, CK => 
                           net2468154, Q => n_1098, QN => n2952);
   IF_CPathxCtlToRegs_port_src2_regx2x : DFF_X1 port map( D => n6431, CK => 
                           net2468154, Q => CtlToRegs_port_src2_2_port, QN => 
                           n6257);
   IF_CPathxCtlToRegs_port_src2_regx3x : DFF_X1 port map( D => n6430, CK => 
                           net2468154, Q => CtlToRegs_port_src2_3_port, QN => 
                           n6265);
   IF_CPathxCtlToRegs_port_src2_regx4x : DFF_X1 port map( D => n6429, CK => 
                           net2468154, Q => CtlToRegs_port_src2_4_port, QN => 
                           n6206);
   IF_CPathxCtlToRegs_port_src1_regx0x : DFF_X1 port map( D => n6428, CK => 
                           net2468154, Q => CtlToRegs_port_src1_0_port, QN => 
                           n6267);
   IF_CPathxCtlToRegs_port_src1_regx1x : DFF_X1 port map( D => n6427, CK => 
                           net2468154, Q => CtlToRegs_port_src1_1_port, QN => 
                           n6194);
   IF_CPathxCtlToRegs_port_src1_regx2x : DFF_X1 port map( D => n6426, CK => 
                           net2468154, Q => CtlToRegs_port_src1_2_port, QN => 
                           n6258);
   IF_CPathxCtlToRegs_port_src1_regx3x : DFF_X1 port map( D => n6425, CK => 
                           net2468154, Q => CtlToRegs_port_src1_3_port, QN => 
                           n6256);
   IF_CPathxCtlToRegs_port_src1_regx4x : DFF_X1 port map( D => n6424, CK => 
                           net2468154, Q => CtlToRegs_port_src1_4_port, QN => 
                           n6205);
   IF_CPathxCtlToRegs_port_req_reg : DFF_X1 port map( D => n6546, CK => 
                           net2468209, Q => CtlToRegs_port_req, QN => n_1099);
   IF_CPathxCtlToRegs_data_signal_dst_regx0x : DFF_X1 port map( D => 
                           IF_CPathxN2033, CK => net2468219, Q => 
                           IF_CPathxCtlToRegs_data_signal_dst_0_port, QN => 
                           n_1100);
   IF_CPathxCtlToRegs_port_dst_regx0x : DFF_X1 port map( D => n6545, CK => 
                           net2468209, Q => CtlToRegs_port_dst_0_port, QN => 
                           n6233);
   IF_CPathxCtlToRegs_data_signal_dst_regx1x : DFF_X1 port map( D => 
                           IF_CPathxN2034, CK => net2468219, Q => 
                           IF_CPathxCtlToRegs_data_signal_dst_1_port, QN => 
                           n_1101);
   IF_CPathxCtlToRegs_port_dst_regx1x : DFF_X1 port map( D => n6544, CK => 
                           net2468209, Q => CtlToRegs_port_dst_1_port, QN => 
                           n6198);
   IF_CPathxCtlToRegs_data_signal_dst_regx2x : DFF_X1 port map( D => 
                           IF_CPathxN2035, CK => net2468219, Q => 
                           IF_CPathxCtlToRegs_data_signal_dst_2_port, QN => 
                           n_1102);
   IF_CPathxCtlToRegs_port_dst_regx2x : DFF_X1 port map( D => n6543, CK => 
                           net2468209, Q => CtlToRegs_port_dst_2_port, QN => 
                           n_1103);
   IF_CPathxCtlToRegs_data_signal_dst_regx3x : DFF_X1 port map( D => 
                           IF_CPathxN2036, CK => net2468219, Q => 
                           IF_CPathxCtlToRegs_data_signal_dst_3_port, QN => 
                           n_1104);
   IF_CPathxCtlToRegs_port_dst_regx3x : DFF_X1 port map( D => n6542, CK => 
                           net2468209, Q => CtlToRegs_port_dst_3_port, QN => 
                           n_1105);
   IF_CPathxCtlToRegs_data_signal_dst_regx4x : DFF_X1 port map( D => 
                           IF_CPathxN2037, CK => net2468219, Q => 
                           IF_CPathxCtlToRegs_data_signal_dst_4_port, QN => 
                           n_1106);
   IF_CPathxCtlToRegs_port_dst_regx4x : DFF_X1 port map( D => n6541, CK => 
                           net2468209, Q => CtlToRegs_port_dst_4_port, QN => 
                           n6235);
   IF_CPathxCtlToMem_port_mask_regx0x : DFF_X1 port map( D => n6501, CK => 
                           net2468164, Q => CtlToMem_port_mask(0), QN => n_1107
                           );
   IF_CPathxCtlToMem_port_mask_regx1x : DFF_X1 port map( D => n6500, CK => 
                           net2468164, Q => CtlToMem_port_mask(1), QN => n_1108
                           );
   IF_CPathxCtlToMem_port_mask_regx2x : DFF_X1 port map( D => n6499, CK => 
                           net2468164, Q => CtlToMem_port_mask(2), QN => n_1109
                           );
   IF_DecoderxDecToCtl_port_imm_regx0x : DFF_X1 port map( D => n6719, CK => 
                           net2468254, Q => DecToCtl_port_imm_0_port, QN => 
                           n_1110);
   IF_CPathxDecToCtl_data_signal_imm_regx0x : DFF_X1 port map( D => 
                           IF_CPathxN2158, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_0_port, QN => 
                           n_1111);
   IF_CPathxCtlToALU_port_imm_regx0x : DFF_X1 port map( D => n6674, CK => 
                           net2468224, Q => CtlToALU_port_imm_0_port, QN => 
                           n_1112);
   IF_DecoderxDecToCtl_port_imm_regx1x : DFF_X1 port map( D => n6718, CK => 
                           net2468254, Q => DecToCtl_port_imm_1_port, QN => 
                           n_1113);
   IF_CPathxDecToCtl_data_signal_imm_regx1x : DFF_X1 port map( D => 
                           IF_CPathxN2159, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_1_port, QN => 
                           n_1114);
   IF_CPathxCtlToALU_port_imm_regx1x : DFF_X1 port map( D => n6673, CK => 
                           net2468224, Q => CtlToALU_port_imm_1_port, QN => 
                           n_1115);
   IF_DecoderxDecToCtl_port_imm_regx2x : DFF_X1 port map( D => n6717, CK => 
                           net2468254, Q => DecToCtl_port_imm_2_port, QN => 
                           n_1116);
   IF_CPathxDecToCtl_data_signal_imm_regx2x : DFF_X1 port map( D => 
                           IF_CPathxN2160, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_2_port, QN => 
                           n_1117);
   IF_CPathxCtlToALU_port_imm_regx2x : DFF_X1 port map( D => n6672, CK => 
                           net2468224, Q => CtlToALU_port_imm_2_port, QN => 
                           n_1118);
   IF_DecoderxDecToCtl_port_imm_regx3x : DFF_X1 port map( D => n6716, CK => 
                           net2468254, Q => n_1119, QN => n6224);
   IF_CPathxDecToCtl_data_signal_imm_regx3x : DFF_X1 port map( D => 
                           IF_CPathxN2161, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_3_port, QN => 
                           n6329);
   IF_CPathxCtlToALU_port_imm_regx3x : DFF_X1 port map( D => n6671, CK => 
                           net2468224, Q => CtlToALU_port_imm_3_port, QN => 
                           n_1120);
   IF_DecoderxDecToCtl_port_imm_regx4x : DFF_X1 port map( D => n6715, CK => 
                           net2468254, Q => DecToCtl_port_imm_4_port, QN => 
                           n_1121);
   IF_CPathxDecToCtl_data_signal_imm_regx4x : DFF_X1 port map( D => 
                           IF_CPathxN2162, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_4_port, QN => 
                           n_1122);
   IF_CPathxCtlToALU_port_imm_regx4x : DFF_X1 port map( D => n6670, CK => 
                           net2468224, Q => CtlToALU_port_imm_4_port, QN => 
                           n_1123);
   IF_DecoderxDecToCtl_port_imm_regx5x : DFF_X1 port map( D => n6714, CK => 
                           net2468254, Q => n_1124, QN => n6218);
   IF_CPathxDecToCtl_data_signal_imm_regx5x : DFF_X1 port map( D => 
                           IF_CPathxN2163, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_5_port, QN => 
                           n6334);
   IF_CPathxCtlToALU_port_imm_regx5x : DFF_X1 port map( D => n6669, CK => 
                           net2468224, Q => CtlToALU_port_imm_5_port, QN => 
                           n_1125);
   IF_DecoderxDecToCtl_port_imm_regx6x : DFF_X1 port map( D => n6713, CK => 
                           net2468254, Q => DecToCtl_port_imm_6_port, QN => 
                           n_1126);
   IF_CPathxDecToCtl_data_signal_imm_regx6x : DFF_X1 port map( D => n6406, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_6_port, QN => 
                           n_1127);
   IF_CPathxCtlToALU_port_imm_regx6x : DFF_X1 port map( D => n6668, CK => 
                           net2468224, Q => CtlToALU_port_imm_6_port, QN => 
                           n_1128);
   IF_DecoderxDecToCtl_port_imm_regx7x : DFF_X1 port map( D => n6712, CK => 
                           net2468254, Q => n_1129, QN => n6219);
   IF_CPathxDecToCtl_data_signal_imm_regx7x : DFF_X1 port map( D => 
                           IF_CPathxN2165, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_7_port, QN => 
                           n6335);
   IF_CPathxCtlToALU_port_imm_regx7x : DFF_X1 port map( D => n6667, CK => 
                           net2468224, Q => CtlToALU_port_imm_7_port, QN => 
                           n_1130);
   IF_DecoderxDecToCtl_port_imm_regx8x : DFF_X1 port map( D => n6711, CK => 
                           net2468254, Q => DecToCtl_port_imm_8_port, QN => 
                           n_1131);
   IF_CPathxDecToCtl_data_signal_imm_regx8x : DFF_X1 port map( D => n6407, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_8_port, QN => 
                           n_1132);
   IF_CPathxCtlToALU_port_imm_regx8x : DFF_X1 port map( D => n6666, CK => 
                           net2468224, Q => CtlToALU_port_imm_8_port, QN => 
                           n_1133);
   IF_DecoderxDecToCtl_port_imm_regx9x : DFF_X1 port map( D => n6710, CK => 
                           net2468254, Q => n_1134, QN => n6217);
   IF_CPathxDecToCtl_data_signal_imm_regx9x : DFF_X1 port map( D => 
                           IF_CPathxN2167, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_9_port, QN => 
                           n6333);
   IF_CPathxCtlToALU_port_imm_regx9x : DFF_X1 port map( D => n6665, CK => 
                           net2468224, Q => CtlToALU_port_imm_9_port, QN => 
                           n_1135);
   IF_DecoderxDecToCtl_port_imm_regx10x : DFF_X1 port map( D => n6709, CK => 
                           net2468254, Q => n_1136, QN => n6220);
   IF_CPathxDecToCtl_data_signal_imm_regx10x : DFF_X1 port map( D => 
                           IF_CPathxN2168, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_10_port, QN => 
                           n6336);
   IF_CPathxCtlToALU_port_imm_regx10x : DFF_X1 port map( D => n6664, CK => 
                           net2468224, Q => CtlToALU_port_imm_10_port, QN => 
                           n_1137);
   IF_DecoderxDecToCtl_port_imm_regx11x : DFF_X1 port map( D => n6708, CK => 
                           net2468254, Q => DecToCtl_port_imm_11_port, QN => 
                           n_1138);
   IF_CPathxDecToCtl_data_signal_imm_regx11x : DFF_X1 port map( D => n6408, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_11_port, QN => 
                           n_1139);
   IF_CPathxCtlToALU_port_imm_regx11x : DFF_X1 port map( D => n6663, CK => 
                           net2468224, Q => CtlToALU_port_imm_11_port, QN => 
                           n_1140);
   IF_DecoderxDecToCtl_port_imm_regx12x : DFF_X1 port map( D => n6707, CK => 
                           net2468254, Q => DecToCtl_port_imm_12_port, QN => 
                           n_1141);
   IF_CPathxDecToCtl_data_signal_imm_regx12x : DFF_X1 port map( D => n6409, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_12_port, QN => 
                           n_1142);
   IF_CPathxCtlToALU_port_imm_regx12x : DFF_X1 port map( D => n6662, CK => 
                           net2468224, Q => CtlToALU_port_imm_12_port, QN => 
                           n_1143);
   IF_DecoderxDecToCtl_port_imm_regx13x : DFF_X1 port map( D => n6706, CK => 
                           net2468254, Q => DecToCtl_port_imm_13_port, QN => 
                           n_1144);
   IF_CPathxDecToCtl_data_signal_imm_regx13x : DFF_X1 port map( D => n6410, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_13_port, QN => 
                           n_1145);
   IF_CPathxCtlToALU_port_imm_regx13x : DFF_X1 port map( D => n6661, CK => 
                           net2468224, Q => CtlToALU_port_imm_13_port, QN => 
                           n_1146);
   IF_DecoderxDecToCtl_port_imm_regx14x : DFF_X1 port map( D => n6705, CK => 
                           net2468254, Q => DecToCtl_port_imm_14_port, QN => 
                           n_1147);
   IF_CPathxDecToCtl_data_signal_imm_regx14x : DFF_X1 port map( D => n6411, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_14_port, QN => 
                           n_1148);
   IF_CPathxCtlToALU_port_imm_regx14x : DFF_X1 port map( D => n6660, CK => 
                           net2468224, Q => CtlToALU_port_imm_14_port, QN => 
                           n_1149);
   IF_DecoderxDecToCtl_port_imm_regx15x : DFF_X1 port map( D => n6704, CK => 
                           net2468254, Q => DecToCtl_port_imm_15_port, QN => 
                           n_1150);
   IF_CPathxDecToCtl_data_signal_imm_regx15x : DFF_X1 port map( D => n6412, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_15_port, QN => 
                           n_1151);
   IF_CPathxCtlToALU_port_imm_regx15x : DFF_X1 port map( D => n6659, CK => 
                           net2468224, Q => CtlToALU_port_imm_15_port, QN => 
                           n_1152);
   IF_DecoderxDecToCtl_port_imm_regx16x : DFF_X1 port map( D => n6703, CK => 
                           net2468254, Q => n_1153, QN => n6221);
   IF_CPathxDecToCtl_data_signal_imm_regx16x : DFF_X1 port map( D => 
                           IF_CPathxN2174, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_16_port, QN => 
                           n6337);
   IF_CPathxCtlToALU_port_imm_regx16x : DFF_X1 port map( D => n6658, CK => 
                           net2468224, Q => CtlToALU_port_imm_16_port, QN => 
                           n_1154);
   IF_DecoderxDecToCtl_port_imm_regx17x : DFF_X1 port map( D => n6702, CK => 
                           net2468254, Q => DecToCtl_port_imm_17_port, QN => 
                           n_1155);
   IF_CPathxDecToCtl_data_signal_imm_regx17x : DFF_X1 port map( D => n6413, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_17_port, QN => 
                           n_1156);
   IF_CPathxCtlToALU_port_imm_regx17x : DFF_X1 port map( D => n6657, CK => 
                           net2468224, Q => CtlToALU_port_imm_17_port, QN => 
                           n_1157);
   IF_DecoderxDecToCtl_port_imm_regx18x : DFF_X1 port map( D => n6701, CK => 
                           net2468254, Q => n_1158, QN => n6222);
   IF_CPathxDecToCtl_data_signal_imm_regx18x : DFF_X1 port map( D => 
                           IF_CPathxN2176, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_18_port, QN => 
                           n6338);
   IF_CPathxCtlToALU_port_imm_regx18x : DFF_X1 port map( D => n6656, CK => 
                           net2468224, Q => CtlToALU_port_imm_18_port, QN => 
                           n_1159);
   IF_DecoderxDecToCtl_port_imm_regx19x : DFF_X1 port map( D => n6700, CK => 
                           net2468254, Q => DecToCtl_port_imm_19_port, QN => 
                           n_1160);
   IF_CPathxDecToCtl_data_signal_imm_regx19x : DFF_X1 port map( D => n6414, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_19_port, QN => 
                           n_1161);
   IF_CPathxCtlToALU_port_imm_regx19x : DFF_X1 port map( D => n6655, CK => 
                           net2468224, Q => CtlToALU_port_imm_19_port, QN => 
                           n_1162);
   IF_DecoderxDecToCtl_port_imm_regx20x : DFF_X1 port map( D => n6699, CK => 
                           net2468254, Q => DecToCtl_port_imm_20_port, QN => 
                           n_1163);
   IF_CPathxDecToCtl_data_signal_imm_regx20x : DFF_X1 port map( D => n6415, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_20_port, QN => 
                           n_1164);
   IF_CPathxCtlToALU_port_imm_regx20x : DFF_X1 port map( D => n6654, CK => 
                           net2468224, Q => CtlToALU_port_imm_20_port, QN => 
                           n_1165);
   IF_DecoderxDecToCtl_port_imm_regx21x : DFF_X1 port map( D => n6698, CK => 
                           net2468254, Q => DecToCtl_port_imm_21_port, QN => 
                           n_1166);
   IF_CPathxDecToCtl_data_signal_imm_regx21x : DFF_X1 port map( D => n6416, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_21_port, QN => 
                           n_1167);
   IF_CPathxCtlToALU_port_imm_regx21x : DFF_X1 port map( D => n6653, CK => 
                           net2468224, Q => CtlToALU_port_imm_21_port, QN => 
                           n_1168);
   IF_DecoderxDecToCtl_port_imm_regx22x : DFF_X1 port map( D => n6697, CK => 
                           net2468254, Q => DecToCtl_port_imm_22_port, QN => 
                           n_1169);
   IF_CPathxDecToCtl_data_signal_imm_regx22x : DFF_X1 port map( D => n6417, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_22_port, QN => 
                           n_1170);
   IF_CPathxCtlToALU_port_imm_regx22x : DFF_X1 port map( D => n6652, CK => 
                           net2468224, Q => CtlToALU_port_imm_22_port, QN => 
                           n_1171);
   IF_DecoderxDecToCtl_port_imm_regx23x : DFF_X1 port map( D => n6696, CK => 
                           net2468254, Q => n_1172, QN => n6215);
   IF_CPathxDecToCtl_data_signal_imm_regx23x : DFF_X1 port map( D => 
                           IF_CPathxN2181, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_23_port, QN => 
                           n6331);
   IF_CPathxCtlToALU_port_imm_regx23x : DFF_X1 port map( D => n6651, CK => 
                           net2468224, Q => CtlToALU_port_imm_23_port, QN => 
                           n_1173);
   IF_DecoderxDecToCtl_port_imm_regx24x : DFF_X1 port map( D => n6695, CK => 
                           net2468254, Q => n_1174, QN => n6216);
   IF_CPathxDecToCtl_data_signal_imm_regx24x : DFF_X1 port map( D => 
                           IF_CPathxN2182, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_24_port, QN => 
                           n6332);
   IF_CPathxCtlToALU_port_imm_regx24x : DFF_X1 port map( D => n6650, CK => 
                           net2468224, Q => CtlToALU_port_imm_24_port, QN => 
                           n_1175);
   IF_DecoderxDecToCtl_port_imm_regx25x : DFF_X1 port map( D => n6694, CK => 
                           net2468254, Q => n_1176, QN => n6214);
   IF_CPathxDecToCtl_data_signal_imm_regx25x : DFF_X1 port map( D => 
                           IF_CPathxN2183, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_25_port, QN => 
                           n6330);
   IF_CPathxCtlToALU_port_imm_regx25x : DFF_X1 port map( D => n6649, CK => 
                           net2468224, Q => CtlToALU_port_imm_25_port, QN => 
                           n_1177);
   IF_DecoderxDecToCtl_port_imm_regx26x : DFF_X1 port map( D => n6693, CK => 
                           net2468254, Q => DecToCtl_port_imm_26_port, QN => 
                           n_1178);
   IF_CPathxDecToCtl_data_signal_imm_regx26x : DFF_X1 port map( D => n6418, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_26_port, QN => 
                           n_1179);
   IF_CPathxCtlToALU_port_imm_regx26x : DFF_X1 port map( D => n6648, CK => 
                           net2468224, Q => CtlToALU_port_imm_26_port, QN => 
                           n_1180);
   IF_DecoderxDecToCtl_port_imm_regx27x : DFF_X1 port map( D => n6692, CK => 
                           net2468254, Q => DecToCtl_port_imm_27_port, QN => 
                           n_1181);
   IF_CPathxDecToCtl_data_signal_imm_regx27x : DFF_X1 port map( D => n6419, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_27_port, QN => 
                           n_1182);
   IF_CPathxCtlToALU_port_imm_regx27x : DFF_X1 port map( D => n6647, CK => 
                           net2468224, Q => CtlToALU_port_imm_27_port, QN => 
                           n_1183);
   IF_DecoderxDecToCtl_port_imm_regx28x : DFF_X1 port map( D => n6691, CK => 
                           net2468254, Q => n_1184, QN => n6223);
   IF_CPathxDecToCtl_data_signal_imm_regx28x : DFF_X1 port map( D => 
                           IF_CPathxN2186, CK => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_28_port, QN => 
                           n6339);
   IF_CPathxCtlToALU_port_imm_regx28x : DFF_X1 port map( D => n6646, CK => 
                           net2468224, Q => CtlToALU_port_imm_28_port, QN => 
                           n_1185);
   IF_DecoderxDecToCtl_port_imm_regx29x : DFF_X1 port map( D => n6690, CK => 
                           net2468254, Q => DecToCtl_port_imm_29_port, QN => 
                           n_1186);
   IF_CPathxDecToCtl_data_signal_imm_regx29x : DFF_X1 port map( D => n6420, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_29_port, QN => 
                           n_1187);
   IF_CPathxCtlToALU_port_imm_regx29x : DFF_X1 port map( D => n6645, CK => 
                           net2468224, Q => CtlToALU_port_imm_29_port, QN => 
                           n_1188);
   IF_DecoderxDecToCtl_port_imm_regx30x : DFF_X1 port map( D => n6689, CK => 
                           net2468254, Q => DecToCtl_port_imm_30_port, QN => 
                           n_1189);
   IF_CPathxDecToCtl_data_signal_imm_regx30x : DFF_X1 port map( D => n6421, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_30_port, QN => 
                           n_1190);
   IF_CPathxCtlToALU_port_imm_regx30x : DFF_X1 port map( D => n6644, CK => 
                           net2468224, Q => CtlToALU_port_imm_30_port, QN => 
                           n_1191);
   IF_DecoderxDecToCtl_port_imm_regx31x : DFF_X1 port map( D => n6688, CK => 
                           net2468254, Q => DecToCtl_port_imm_31_port, QN => 
                           n_1192);
   IF_CPathxDecToCtl_data_signal_imm_regx31x : DFF_X1 port map( D => n6422, CK 
                           => net2468194, Q => 
                           IF_CPathxDecToCtl_data_signal_imm_31_port, QN => 
                           n_1193);
   IF_CPathxCtlToALU_port_imm_regx31x : DFF_X1 port map( D => n6643, CK => 
                           net2468224, Q => CtlToALU_port_imm_31_port, QN => 
                           n_1194);
   IF_CPathxmemoryAccess_signal_req_reg : DFF_X1 port map( D => n6685, CK => 
                           net2468239, Q => n_1195, QN => n6286);
   IF_CPathxCtlToMem_port_req_reg : DFF_X1 port map( D => n6498, CK => 
                           net2468164, Q => CtlToMem_port_req, QN => n_1196);
   IF_CPathxMemToCtl_port_notify_reg : DFF_X1 port map( D => n2944, CK => 
                           net2468239, Q => MemToCtl_port_notify_port, QN => 
                           n_1197);
   IF_CPathxCtlToMem_port_notify_reg : DFF_X1 port map( D => n6684, CK => 
                           net2468239, Q => CtlToMem_port_notify_port, QN => 
                           n_1198);
   IF_CPathxCtlToALU_port_notify_reg : DFF_X1 port map( D => n6683, CK => 
                           net2468239, Q => CtlToALU_port_notify, QN => n_1199)
                           ;
   IF_CPathxCtlToRegs_port_notify_reg : DFF_X1 port map( D => n6682, CK => 
                           net2468239, Q => CtlToRegs_port_notify, QN => n6237)
                           ;
   IF_RegsxRegsToCtl_port_contents1_regx31x : DFF_X1 port map( D => 
                           IF_RegsxN626, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_31_port, QN => n_1200);
   IF_CPathxRegsToCtl_data_signal_contents1_regx31x : DFF_X1 port map( D => 
                           n6405, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_31_port, QN
                           => n6346);
   IF_CPathxCtlToALU_port_reg1_contents_regx31x : DFF_X1 port map( D => n6642, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_31_port, QN => n_1201);
   IF_ALUxALUtoCtl_port_regx31x : DFF_X1 port map( D => IF_ALUxN969, CK => 
                           net2468144, Q => ALUtoCtl_port_31_port, QN => n6279)
                           ;
   IF_CPathxpc_next_signal_regx0x : DFF_X1 port map( D => IF_CPathxN2242, CK =>
                           net2468179, Q => IF_CPathxpc_next_signal_0_port, QN 
                           => n_1202);
   IF_CPathxpc_reg_signal_regx0x : DFF_X1 port map( D => n6537, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_0_port, QN 
                           => n_1203);
   IF_CPathxCtlToALU_port_pc_reg_regx0x : DFF_X1 port map( D => IF_CPathxN1936,
                           CK => net2468224, Q => CtlToALU_port_pc_reg_0_port, 
                           QN => n_1204);
   IF_CPathxpc_next_signal_regx1x : DFF_X1 port map( D => IF_CPathxN2243, CK =>
                           net2468179, Q => IF_CPathxpc_next_signal_1_port, QN 
                           => n_1205);
   IF_CPathxpc_reg_signal_regx1x : DFF_X1 port map( D => n6536, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_1_port, QN 
                           => n6323);
   IF_CPathxCtlToALU_port_pc_reg_regx1x : DFF_X1 port map( D => IF_CPathxN1937,
                           CK => net2468224, Q => CtlToALU_port_pc_reg_1_port, 
                           QN => n_1206);
   IF_CPathxpc_next_signal_regx2x : DFF_X1 port map( D => IF_CPathxN2244, CK =>
                           net2468179, Q => IF_CPathxpc_next_signal_2_port, QN 
                           => n_1207);
   IF_CPathxpc_reg_signal_regx2x : DFF_X1 port map( D => n6535, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_2_port, QN 
                           => n6245);
   IF_CPathxCtlToALU_port_pc_reg_regx2x : DFF_X1 port map( D => IF_CPathxN1938,
                           CK => net2468224, Q => CtlToALU_port_pc_reg_2_port, 
                           QN => n_1208);
   IF_CPathxpc_next_signal_regx3x : DFF_X1 port map( D => IF_CPathxN2245, CK =>
                           net2468179, Q => IF_CPathxpc_next_signal_3_port, QN 
                           => n_1209);
   IF_CPathxpc_reg_signal_regx3x : DFF_X1 port map( D => n6534, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_3_port, QN 
                           => n6204);
   IF_CPathxCtlToALU_port_pc_reg_regx3x : DFF_X1 port map( D => IF_CPathxN1939,
                           CK => net2468224, Q => CtlToALU_port_pc_reg_3_port, 
                           QN => n_1210);
   IF_CPathxpc_next_signal_regx4x : DFF_X1 port map( D => IF_CPathxN2246, CK =>
                           net2468179, Q => IF_CPathxpc_next_signal_4_port, QN 
                           => n_1211);
   IF_CPathxpc_reg_signal_regx4x : DFF_X1 port map( D => n6533, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_4_port, QN 
                           => n_1212);
   IF_CPathxCtlToALU_port_pc_reg_regx4x : DFF_X1 port map( D => IF_CPathxN1940,
                           CK => net2468224, Q => CtlToALU_port_pc_reg_4_port, 
                           QN => n_1213);
   IF_CPathxpc_next_signal_regx5x : DFF_X1 port map( D => IF_CPathxN2247, CK =>
                           net2468179, Q => IF_CPathxpc_next_signal_5_port, QN 
                           => n_1214);
   IF_CPathxpc_reg_signal_regx5x : DFF_X1 port map( D => n6532, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_5_port, QN 
                           => n6243);
   IF_CPathxCtlToALU_port_pc_reg_regx5x : DFF_X1 port map( D => IF_CPathxN1941,
                           CK => net2468224, Q => CtlToALU_port_pc_reg_5_port, 
                           QN => n_1215);
   IF_CPathxpc_next_signal_regx6x : DFF_X1 port map( D => IF_CPathxN2248, CK =>
                           net2468179, Q => IF_CPathxpc_next_signal_6_port, QN 
                           => n_1216);
   IF_CPathxpc_reg_signal_regx6x : DFF_X1 port map( D => n6531, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_6_port, QN 
                           => n_1217);
   IF_CPathxCtlToALU_port_pc_reg_regx6x : DFF_X1 port map( D => IF_CPathxN1942,
                           CK => net2468224, Q => CtlToALU_port_pc_reg_6_port, 
                           QN => n_1218);
   IF_CPathxpc_next_signal_regx7x : DFF_X1 port map( D => IF_CPathxN2249, CK =>
                           net2468179, Q => IF_CPathxpc_next_signal_7_port, QN 
                           => n_1219);
   IF_CPathxpc_reg_signal_regx7x : DFF_X1 port map( D => n6530, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_7_port, QN 
                           => n6244);
   IF_CPathxCtlToALU_port_pc_reg_regx7x : DFF_X1 port map( D => IF_CPathxN1943,
                           CK => net2468224, Q => CtlToALU_port_pc_reg_7_port, 
                           QN => n_1220);
   IF_CPathxpc_next_signal_regx8x : DFF_X1 port map( D => IF_CPathxN2250, CK =>
                           net2468179, Q => IF_CPathxpc_next_signal_8_port, QN 
                           => n_1221);
   IF_CPathxpc_reg_signal_regx8x : DFF_X1 port map( D => n6529, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_8_port, QN 
                           => n_1222);
   IF_CPathxCtlToALU_port_pc_reg_regx8x : DFF_X1 port map( D => IF_CPathxN1944,
                           CK => net2468224, Q => CtlToALU_port_pc_reg_8_port, 
                           QN => n_1223);
   IF_CPathxpc_next_signal_regx9x : DFF_X1 port map( D => IF_CPathxN2251, CK =>
                           net2468179, Q => IF_CPathxpc_next_signal_9_port, QN 
                           => n_1224);
   IF_CPathxpc_reg_signal_regx9x : DFF_X1 port map( D => n6528, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_9_port, QN 
                           => n6247);
   IF_CPathxCtlToALU_port_pc_reg_regx9x : DFF_X1 port map( D => IF_CPathxN1945,
                           CK => net2468224, Q => CtlToALU_port_pc_reg_9_port, 
                           QN => n_1225);
   IF_CPathxpc_next_signal_regx10x : DFF_X1 port map( D => IF_CPathxN2252, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_10_port,
                           QN => n_1226);
   IF_CPathxpc_reg_signal_regx10x : DFF_X1 port map( D => n6527, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_10_port, QN 
                           => n_1227);
   IF_CPathxCtlToALU_port_pc_reg_regx10x : DFF_X1 port map( D => IF_CPathxN1946
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_10_port, QN => n_1228);
   IF_CPathxpc_next_signal_regx11x : DFF_X1 port map( D => IF_CPathxN2253, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_11_port,
                           QN => n_1229);
   IF_CPathxpc_reg_signal_regx11x : DFF_X1 port map( D => n6526, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_11_port, QN 
                           => n6248);
   IF_CPathxCtlToALU_port_pc_reg_regx11x : DFF_X1 port map( D => IF_CPathxN1947
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_11_port, QN => n_1230);
   IF_CPathxpc_next_signal_regx12x : DFF_X1 port map( D => IF_CPathxN2254, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_12_port,
                           QN => n_1231);
   IF_CPathxpc_reg_signal_regx12x : DFF_X1 port map( D => n6525, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_12_port, QN 
                           => n_1232);
   IF_CPathxCtlToALU_port_pc_reg_regx12x : DFF_X1 port map( D => IF_CPathxN1948
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_12_port, QN => n_1233);
   IF_CPathxpc_next_signal_regx13x : DFF_X1 port map( D => IF_CPathxN2255, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_13_port,
                           QN => n_1234);
   IF_CPathxpc_reg_signal_regx13x : DFF_X1 port map( D => n6524, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_13_port, QN 
                           => n6249);
   IF_CPathxCtlToALU_port_pc_reg_regx13x : DFF_X1 port map( D => IF_CPathxN1949
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_13_port, QN => n_1235);
   IF_CPathxpc_next_signal_regx14x : DFF_X1 port map( D => IF_CPathxN2256, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_14_port,
                           QN => n_1236);
   IF_CPathxpc_reg_signal_regx14x : DFF_X1 port map( D => n6523, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_14_port, QN 
                           => n_1237);
   IF_CPathxCtlToALU_port_pc_reg_regx14x : DFF_X1 port map( D => IF_CPathxN1950
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_14_port, QN => n_1238);
   IF_CPathxpc_next_signal_regx15x : DFF_X1 port map( D => IF_CPathxN2257, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_15_port,
                           QN => n_1239);
   IF_CPathxpc_reg_signal_regx15x : DFF_X1 port map( D => n6522, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_15_port, QN 
                           => n6250);
   IF_CPathxCtlToALU_port_pc_reg_regx15x : DFF_X1 port map( D => IF_CPathxN1951
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_15_port, QN => n_1240);
   IF_CPathxpc_next_signal_regx16x : DFF_X1 port map( D => IF_CPathxN2258, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_16_port,
                           QN => n_1241);
   IF_CPathxpc_reg_signal_regx16x : DFF_X1 port map( D => n6521, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_16_port, QN 
                           => n_1242);
   IF_CPathxCtlToALU_port_pc_reg_regx16x : DFF_X1 port map( D => IF_CPathxN1952
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_16_port, QN => n_1243);
   IF_CPathxpc_next_signal_regx17x : DFF_X1 port map( D => IF_CPathxN2259, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_17_port,
                           QN => n_1244);
   IF_CPathxpc_reg_signal_regx17x : DFF_X1 port map( D => n6520, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_17_port, QN 
                           => n6251);
   IF_CPathxCtlToALU_port_pc_reg_regx17x : DFF_X1 port map( D => IF_CPathxN1953
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_17_port, QN => n_1245);
   IF_CPathxpc_next_signal_regx18x : DFF_X1 port map( D => IF_CPathxN2260, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_18_port,
                           QN => n_1246);
   IF_CPathxpc_reg_signal_regx18x : DFF_X1 port map( D => n6519, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_18_port, QN 
                           => n_1247);
   IF_CPathxCtlToALU_port_pc_reg_regx18x : DFF_X1 port map( D => IF_CPathxN1954
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_18_port, QN => n_1248);
   IF_CPathxpc_next_signal_regx19x : DFF_X1 port map( D => IF_CPathxN2261, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_19_port,
                           QN => n_1249);
   IF_CPathxpc_reg_signal_regx19x : DFF_X1 port map( D => n6518, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_19_port, QN 
                           => n6252);
   IF_CPathxCtlToALU_port_pc_reg_regx19x : DFF_X1 port map( D => IF_CPathxN1955
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_19_port, QN => n_1250);
   IF_CPathxpc_next_signal_regx20x : DFF_X1 port map( D => IF_CPathxN2262, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_20_port,
                           QN => n_1251);
   IF_CPathxpc_reg_signal_regx20x : DFF_X1 port map( D => n6517, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_20_port, QN 
                           => n_1252);
   IF_CPathxCtlToALU_port_pc_reg_regx20x : DFF_X1 port map( D => IF_CPathxN1956
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_20_port, QN => n_1253);
   IF_CPathxpc_next_signal_regx21x : DFF_X1 port map( D => IF_CPathxN2263, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_21_port,
                           QN => n_1254);
   IF_CPathxpc_reg_signal_regx21x : DFF_X1 port map( D => n6516, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_21_port, QN 
                           => n6253);
   IF_CPathxCtlToALU_port_pc_reg_regx21x : DFF_X1 port map( D => IF_CPathxN1957
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_21_port, QN => n_1255);
   IF_CPathxpc_next_signal_regx22x : DFF_X1 port map( D => IF_CPathxN2264, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_22_port,
                           QN => n_1256);
   IF_CPathxpc_reg_signal_regx22x : DFF_X1 port map( D => n6515, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_22_port, QN 
                           => n_1257);
   IF_CPathxCtlToALU_port_pc_reg_regx22x : DFF_X1 port map( D => IF_CPathxN1958
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_22_port, QN => n_1258);
   IF_CPathxpc_next_signal_regx23x : DFF_X1 port map( D => IF_CPathxN2265, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_23_port,
                           QN => n_1259);
   IF_CPathxpc_reg_signal_regx23x : DFF_X1 port map( D => n6514, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_23_port, QN 
                           => n6254);
   IF_CPathxCtlToALU_port_pc_reg_regx23x : DFF_X1 port map( D => IF_CPathxN1959
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_23_port, QN => n_1260);
   IF_CPathxpc_next_signal_regx24x : DFF_X1 port map( D => IF_CPathxN2266, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_24_port,
                           QN => n_1261);
   IF_CPathxpc_reg_signal_regx24x : DFF_X1 port map( D => n6513, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_24_port, QN 
                           => n_1262);
   IF_CPathxCtlToALU_port_pc_reg_regx24x : DFF_X1 port map( D => IF_CPathxN1960
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_24_port, QN => n_1263);
   IF_CPathxpc_next_signal_regx25x : DFF_X1 port map( D => IF_CPathxN2267, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_25_port,
                           QN => n_1264);
   IF_CPathxpc_reg_signal_regx25x : DFF_X1 port map( D => n6512, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_25_port, QN 
                           => n6255);
   IF_CPathxCtlToALU_port_pc_reg_regx25x : DFF_X1 port map( D => IF_CPathxN1961
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_25_port, QN => n_1265);
   IF_CPathxpc_next_signal_regx26x : DFF_X1 port map( D => IF_CPathxN2268, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_26_port,
                           QN => n_1266);
   IF_CPathxpc_reg_signal_regx26x : DFF_X1 port map( D => n6511, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_26_port, QN 
                           => n_1267);
   IF_CPathxCtlToALU_port_pc_reg_regx26x : DFF_X1 port map( D => IF_CPathxN1962
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_26_port, QN => n_1268);
   IF_CPathxpc_next_signal_regx27x : DFF_X1 port map( D => IF_CPathxN2269, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_27_port,
                           QN => n_1269);
   IF_CPathxpc_reg_signal_regx27x : DFF_X1 port map( D => n6510, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_27_port, QN 
                           => n6262);
   IF_CPathxCtlToALU_port_pc_reg_regx27x : DFF_X1 port map( D => IF_CPathxN1963
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_27_port, QN => n_1270);
   IF_CPathxpc_next_signal_regx28x : DFF_X1 port map( D => IF_CPathxN2270, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_28_port,
                           QN => n_1271);
   IF_CPathxpc_reg_signal_regx28x : DFF_X1 port map( D => n6509, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_28_port, QN 
                           => n_1272);
   IF_CPathxCtlToALU_port_pc_reg_regx28x : DFF_X1 port map( D => IF_CPathxN1964
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_28_port, QN => n_1273);
   IF_CPathxpc_next_signal_regx29x : DFF_X1 port map( D => IF_CPathxN2271, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_29_port,
                           QN => n_1274);
   IF_CPathxpc_reg_signal_regx29x : DFF_X1 port map( D => n6508, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_29_port, QN 
                           => n6263);
   IF_CPathxCtlToALU_port_pc_reg_regx29x : DFF_X1 port map( D => IF_CPathxN1965
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_29_port, QN => n_1275);
   IF_CPathxpc_next_signal_regx30x : DFF_X1 port map( D => n6423, CK => 
                           net2468179, Q => IF_CPathxpc_next_signal_30_port, QN
                           => n_1276);
   IF_CPathxpc_reg_signal_regx30x : DFF_X1 port map( D => n6507, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_30_port, QN 
                           => n_1277);
   IF_CPathxCtlToALU_port_pc_reg_regx30x : DFF_X1 port map( D => IF_CPathxN1966
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_30_port, QN => n_1278);
   IF_ALUxALUtoCtl_port_regx0x : DFF_X1 port map( D => IF_ALUxN938, CK => 
                           net2468144, Q => ALUtoCtl_port_0_port, QN => n6238);
   IF_CPathxALUtoCtl_data_signal_regx0x : DFF_X1 port map( D => IF_CPathxN1860,
                           CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_0_port, QN => n_1279);
   IF_CPathxCtlToMem_port_addrIn_regx0x : DFF_X1 port map( D => n6497, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(0), QN => 
                           n_1280);
   IF_CPathxCtlToRegs_port_dst_data_regx0x : DFF_X1 port map( D => n6578, CK =>
                           net2468214, Q => CtlToRegs_port_dst_data_0_port, QN 
                           => n_1281);
   IF_Regsxreg_file_regx31xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468259, Q => IF_Regsxreg_file_0_port, QN => 
                           n_1282);
   IF_Regsxreg_file_regx1xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468409, Q => IF_Regsxreg_file_960_port, QN => 
                           n_1283);
   IF_Regsxreg_file_regx2xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468404, Q => IF_Regsxreg_file_928_port, QN => 
                           n_1284);
   IF_Regsxreg_file_regx3xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468399, Q => IF_Regsxreg_file_896_port, QN => 
                           n_1285);
   IF_Regsxreg_file_regx4xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468394, Q => IF_Regsxreg_file_864_port, QN => 
                           n_1286);
   IF_Regsxreg_file_regx5xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468389, Q => IF_Regsxreg_file_832_port, QN => 
                           n_1287);
   IF_Regsxreg_file_regx6xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468384, Q => IF_Regsxreg_file_800_port, QN => 
                           n_1288);
   IF_Regsxreg_file_regx7xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468379, Q => IF_Regsxreg_file_768_port, QN => 
                           n_1289);
   IF_Regsxreg_file_regx8xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468374, Q => IF_Regsxreg_file_736_port, QN => 
                           n_1290);
   IF_Regsxreg_file_regx9xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468369, Q => IF_Regsxreg_file_704_port, QN => 
                           n_1291);
   IF_Regsxreg_file_regx10xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468364, Q => IF_Regsxreg_file_672_port, QN => 
                           n_1292);
   IF_Regsxreg_file_regx11xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468359, Q => IF_Regsxreg_file_640_port, QN => 
                           n_1293);
   IF_Regsxreg_file_regx12xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468354, Q => IF_Regsxreg_file_608_port, QN => 
                           n_1294);
   IF_Regsxreg_file_regx13xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468349, Q => IF_Regsxreg_file_576_port, QN => 
                           n_1295);
   IF_Regsxreg_file_regx14xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468344, Q => IF_Regsxreg_file_544_port, QN => 
                           n_1296);
   IF_Regsxreg_file_regx15xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468339, Q => IF_Regsxreg_file_512_port, QN => 
                           n_1297);
   IF_Regsxreg_file_regx16xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468334, Q => IF_Regsxreg_file_480_port, QN => 
                           n_1298);
   IF_Regsxreg_file_regx17xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468329, Q => IF_Regsxreg_file_448_port, QN => 
                           n_1299);
   IF_Regsxreg_file_regx18xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468324, Q => IF_Regsxreg_file_416_port, QN => 
                           n_1300);
   IF_Regsxreg_file_regx19xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468319, Q => IF_Regsxreg_file_384_port, QN => 
                           n_1301);
   IF_Regsxreg_file_regx20xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468314, Q => IF_Regsxreg_file_352_port, QN => 
                           n_1302);
   IF_Regsxreg_file_regx21xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468309, Q => IF_Regsxreg_file_320_port, QN => 
                           n_1303);
   IF_Regsxreg_file_regx22xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468304, Q => IF_Regsxreg_file_288_port, QN => 
                           n_1304);
   IF_Regsxreg_file_regx23xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468299, Q => IF_Regsxreg_file_256_port, QN => 
                           n_1305);
   IF_Regsxreg_file_regx24xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468294, Q => IF_Regsxreg_file_224_port, QN => 
                           n_1306);
   IF_Regsxreg_file_regx25xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468289, Q => IF_Regsxreg_file_192_port, QN => 
                           n_1307);
   IF_Regsxreg_file_regx26xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468284, Q => IF_Regsxreg_file_160_port, QN => 
                           n_1308);
   IF_Regsxreg_file_regx27xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468279, Q => IF_Regsxreg_file_128_port, QN => 
                           n_1309);
   IF_Regsxreg_file_regx28xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468274, Q => IF_Regsxreg_file_96_port, QN => 
                           n_1310);
   IF_Regsxreg_file_regx29xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468269, Q => IF_Regsxreg_file_64_port, QN => 
                           n_1311);
   IF_Regsxreg_file_regx30xx0x : DFF_X1 port map( D => IF_RegsxN660, CK => 
                           net2468264, Q => IF_Regsxreg_file_32_port, QN => 
                           n_1312);
   IF_RegsxRegsToCtl_port_contents2_regx0x : DFF_X1 port map( D => IF_RegsxN627
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents2_0_port, QN => n_1313);
   IF_CPathxRegsToCtl_data_signal_contents2_regx0x : DFF_X1 port map( D => 
                           IF_CPathxN2124, CK => net2468199, Q => n_1314, QN =>
                           n6287);
   IF_CPathxCtlToMem_port_dataIn_regx0x : DFF_X1 port map( D => n6496, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(0), QN => 
                           n_1315);
   IF_CPathxCtlToALU_port_reg2_contents_regx0x : DFF_X1 port map( D => n6641, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_0_port, QN => n_1316);
   IF_RegsxRegsToCtl_port_contents1_regx0x : DFF_X1 port map( D => IF_RegsxN595
                           , CK => net2468414, Q => n_1317, QN => n6373);
   IF_CPathxRegsToCtl_data_signal_contents1_regx0x : DFF_X1 port map( D => 
                           IF_CPathxN2090, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_0_port, QN 
                           => n6340);
   IF_CPathxCtlToALU_port_reg1_contents_regx0x : DFF_X1 port map( D => n6640, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_0_port, QN => n_1318);
   IF_ALUxALUtoCtl_port_regx16x : DFF_X1 port map( D => IF_ALUxN954, CK => 
                           net2468144, Q => ALUtoCtl_port_16_port, QN => n6278)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx16x : DFF_X1 port map( D => IF_CPathxN1876
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_16_port, QN => n_1319)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx16x : DFF_X1 port map( D => n6495, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(16), QN => 
                           n_1320);
   IF_CPathxCtlToRegs_port_dst_data_regx16x : DFF_X1 port map( D => n6577, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_16_port,
                           QN => n_1321);
   IF_Regsxreg_file_regx31xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468259, Q => IF_Regsxreg_file_16_port, QN => 
                           n_1322);
   IF_Regsxreg_file_regx1xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468409, Q => IF_Regsxreg_file_976_port, QN => 
                           n_1323);
   IF_Regsxreg_file_regx2xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468404, Q => IF_Regsxreg_file_944_port, QN => 
                           n_1324);
   IF_Regsxreg_file_regx3xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468399, Q => IF_Regsxreg_file_912_port, QN => 
                           n_1325);
   IF_Regsxreg_file_regx4xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468394, Q => IF_Regsxreg_file_880_port, QN => 
                           n_1326);
   IF_Regsxreg_file_regx5xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468389, Q => IF_Regsxreg_file_848_port, QN => 
                           n_1327);
   IF_Regsxreg_file_regx6xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468384, Q => IF_Regsxreg_file_816_port, QN => 
                           n_1328);
   IF_Regsxreg_file_regx7xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468379, Q => IF_Regsxreg_file_784_port, QN => 
                           n_1329);
   IF_Regsxreg_file_regx8xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468374, Q => IF_Regsxreg_file_752_port, QN => 
                           n_1330);
   IF_Regsxreg_file_regx9xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468369, Q => IF_Regsxreg_file_720_port, QN => 
                           n_1331);
   IF_Regsxreg_file_regx10xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468364, Q => IF_Regsxreg_file_688_port, QN => 
                           n_1332);
   IF_Regsxreg_file_regx11xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468359, Q => IF_Regsxreg_file_656_port, QN => 
                           n_1333);
   IF_Regsxreg_file_regx12xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468354, Q => IF_Regsxreg_file_624_port, QN => 
                           n_1334);
   IF_Regsxreg_file_regx13xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468349, Q => IF_Regsxreg_file_592_port, QN => 
                           n_1335);
   IF_Regsxreg_file_regx14xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468344, Q => IF_Regsxreg_file_560_port, QN => 
                           n_1336);
   IF_Regsxreg_file_regx15xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468339, Q => IF_Regsxreg_file_528_port, QN => 
                           n_1337);
   IF_Regsxreg_file_regx16xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468334, Q => IF_Regsxreg_file_496_port, QN => 
                           n_1338);
   IF_Regsxreg_file_regx17xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468329, Q => IF_Regsxreg_file_464_port, QN => 
                           n_1339);
   IF_Regsxreg_file_regx18xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468324, Q => IF_Regsxreg_file_432_port, QN => 
                           n_1340);
   IF_Regsxreg_file_regx19xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468319, Q => IF_Regsxreg_file_400_port, QN => 
                           n_1341);
   IF_Regsxreg_file_regx20xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468314, Q => IF_Regsxreg_file_368_port, QN => 
                           n_1342);
   IF_Regsxreg_file_regx21xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468309, Q => IF_Regsxreg_file_336_port, QN => 
                           n_1343);
   IF_Regsxreg_file_regx22xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468304, Q => IF_Regsxreg_file_304_port, QN => 
                           n_1344);
   IF_Regsxreg_file_regx23xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468299, Q => IF_Regsxreg_file_272_port, QN => 
                           n_1345);
   IF_Regsxreg_file_regx24xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468294, Q => IF_Regsxreg_file_240_port, QN => 
                           n_1346);
   IF_Regsxreg_file_regx25xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468289, Q => IF_Regsxreg_file_208_port, QN => 
                           n_1347);
   IF_Regsxreg_file_regx26xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468284, Q => IF_Regsxreg_file_176_port, QN => 
                           n_1348);
   IF_Regsxreg_file_regx27xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468279, Q => IF_Regsxreg_file_144_port, QN => 
                           n_1349);
   IF_Regsxreg_file_regx28xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468274, Q => IF_Regsxreg_file_112_port, QN => 
                           n_1350);
   IF_Regsxreg_file_regx29xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468269, Q => IF_Regsxreg_file_80_port, QN => 
                           n_1351);
   IF_Regsxreg_file_regx30xx16x : DFF_X1 port map( D => IF_RegsxN676, CK => 
                           net2468264, Q => IF_Regsxreg_file_48_port, QN => 
                           n_1352);
   IF_RegsxRegsToCtl_port_contents2_regx16x : DFF_X1 port map( D => 
                           IF_RegsxN643, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_16_port, QN => n_1353);
   IF_CPathxRegsToCtl_data_signal_contents2_regx16x : DFF_X1 port map( D => 
                           IF_CPathxN2140, CK => net2468199, Q => n_1354, QN =>
                           n6288);
   IF_CPathxCtlToMem_port_dataIn_regx16x : DFF_X1 port map( D => n6494, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(16), QN => 
                           n_1355);
   IF_CPathxCtlToALU_port_reg2_contents_regx16x : DFF_X1 port map( D => n6639, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_16_port, QN => n_1356);
   IF_RegsxRegsToCtl_port_contents1_regx16x : DFF_X1 port map( D => 
                           IF_RegsxN611, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_16_port, QN => n_1357);
   IF_CPathxRegsToCtl_data_signal_contents1_regx16x : DFF_X1 port map( D => 
                           n6390, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_16_port, QN
                           => n6365);
   IF_CPathxCtlToALU_port_reg1_contents_regx16x : DFF_X1 port map( D => n6638, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_16_port, QN => n_1358);
   IF_ALUxALUtoCtl_port_regx24x : DFF_X1 port map( D => IF_ALUxN962, CK => 
                           net2468144, Q => ALUtoCtl_port_24_port, QN => n_1359
                           );
   IF_CPathxALUtoCtl_data_signal_regx24x : DFF_X1 port map( D => IF_CPathxN1884
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_24_port, QN => n_1360)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx24x : DFF_X1 port map( D => n6493, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(24), QN => 
                           n_1361);
   IF_CPathxCtlToRegs_port_dst_data_regx24x : DFF_X1 port map( D => n6576, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_24_port,
                           QN => n_1362);
   IF_Regsxreg_file_regx31xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468259, Q => IF_Regsxreg_file_24_port, QN => 
                           n_1363);
   IF_Regsxreg_file_regx1xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468409, Q => IF_Regsxreg_file_984_port, QN => 
                           n_1364);
   IF_Regsxreg_file_regx2xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468404, Q => IF_Regsxreg_file_952_port, QN => 
                           n_1365);
   IF_Regsxreg_file_regx3xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468399, Q => IF_Regsxreg_file_920_port, QN => 
                           n_1366);
   IF_Regsxreg_file_regx4xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468394, Q => IF_Regsxreg_file_888_port, QN => 
                           n_1367);
   IF_Regsxreg_file_regx5xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468389, Q => IF_Regsxreg_file_856_port, QN => 
                           n_1368);
   IF_Regsxreg_file_regx6xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468384, Q => IF_Regsxreg_file_824_port, QN => 
                           n_1369);
   IF_Regsxreg_file_regx7xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468379, Q => IF_Regsxreg_file_792_port, QN => 
                           n_1370);
   IF_Regsxreg_file_regx8xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468374, Q => IF_Regsxreg_file_760_port, QN => 
                           n_1371);
   IF_Regsxreg_file_regx9xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468369, Q => IF_Regsxreg_file_728_port, QN => 
                           n_1372);
   IF_Regsxreg_file_regx10xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468364, Q => IF_Regsxreg_file_696_port, QN => 
                           n_1373);
   IF_Regsxreg_file_regx11xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468359, Q => IF_Regsxreg_file_664_port, QN => 
                           n_1374);
   IF_Regsxreg_file_regx12xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468354, Q => IF_Regsxreg_file_632_port, QN => 
                           n_1375);
   IF_Regsxreg_file_regx13xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468349, Q => IF_Regsxreg_file_600_port, QN => 
                           n_1376);
   IF_Regsxreg_file_regx14xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468344, Q => IF_Regsxreg_file_568_port, QN => 
                           n_1377);
   IF_Regsxreg_file_regx15xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468339, Q => IF_Regsxreg_file_536_port, QN => 
                           n_1378);
   IF_Regsxreg_file_regx16xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468334, Q => IF_Regsxreg_file_504_port, QN => 
                           n_1379);
   IF_Regsxreg_file_regx17xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468329, Q => IF_Regsxreg_file_472_port, QN => 
                           n_1380);
   IF_Regsxreg_file_regx18xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468324, Q => IF_Regsxreg_file_440_port, QN => 
                           n_1381);
   IF_Regsxreg_file_regx19xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468319, Q => IF_Regsxreg_file_408_port, QN => 
                           n_1382);
   IF_Regsxreg_file_regx20xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468314, Q => IF_Regsxreg_file_376_port, QN => 
                           n_1383);
   IF_Regsxreg_file_regx21xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468309, Q => IF_Regsxreg_file_344_port, QN => 
                           n_1384);
   IF_Regsxreg_file_regx22xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468304, Q => IF_Regsxreg_file_312_port, QN => 
                           n_1385);
   IF_Regsxreg_file_regx23xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468299, Q => IF_Regsxreg_file_280_port, QN => 
                           n_1386);
   IF_Regsxreg_file_regx24xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468294, Q => IF_Regsxreg_file_248_port, QN => 
                           n_1387);
   IF_Regsxreg_file_regx25xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468289, Q => IF_Regsxreg_file_216_port, QN => 
                           n_1388);
   IF_Regsxreg_file_regx26xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468284, Q => IF_Regsxreg_file_184_port, QN => 
                           n_1389);
   IF_Regsxreg_file_regx27xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468279, Q => IF_Regsxreg_file_152_port, QN => 
                           n_1390);
   IF_Regsxreg_file_regx28xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468274, Q => IF_Regsxreg_file_120_port, QN => 
                           n_1391);
   IF_Regsxreg_file_regx29xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468269, Q => IF_Regsxreg_file_88_port, QN => 
                           n_1392);
   IF_Regsxreg_file_regx30xx24x : DFF_X1 port map( D => IF_RegsxN684, CK => 
                           net2468264, Q => IF_Regsxreg_file_56_port, QN => 
                           n_1393);
   IF_RegsxRegsToCtl_port_contents2_regx24x : DFF_X1 port map( D => 
                           IF_RegsxN651, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_24_port, QN => n_1394);
   IF_CPathxRegsToCtl_data_signal_contents2_regx24x : DFF_X1 port map( D => 
                           IF_CPathxN2148, CK => net2468199, Q => n_1395, QN =>
                           n6289);
   IF_CPathxCtlToMem_port_dataIn_regx24x : DFF_X1 port map( D => n6492, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(24), QN => 
                           n_1396);
   IF_CPathxCtlToALU_port_reg2_contents_regx24x : DFF_X1 port map( D => n6637, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_24_port, QN => n_1397);
   IF_RegsxRegsToCtl_port_contents1_regx24x : DFF_X1 port map( D => 
                           IF_RegsxN619, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_24_port, QN => n_1398);
   IF_CPathxRegsToCtl_data_signal_contents1_regx24x : DFF_X1 port map( D => 
                           n6398, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_24_port, QN
                           => n6353);
   IF_CPathxCtlToALU_port_reg1_contents_regx24x : DFF_X1 port map( D => n6636, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_24_port, QN => n_1399);
   IF_ALUxALUtoCtl_port_regx28x : DFF_X1 port map( D => IF_ALUxN966, CK => 
                           net2468144, Q => ALUtoCtl_port_28_port, QN => n6284)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx28x : DFF_X1 port map( D => IF_CPathxN1888
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_28_port, QN => n_1400)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx28x : DFF_X1 port map( D => n6491, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(28), QN => 
                           n_1401);
   IF_CPathxCtlToRegs_port_dst_data_regx28x : DFF_X1 port map( D => n6575, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_28_port,
                           QN => n_1402);
   IF_Regsxreg_file_regx31xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468259, Q => IF_Regsxreg_file_28_port, QN => 
                           n_1403);
   IF_Regsxreg_file_regx1xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468409, Q => IF_Regsxreg_file_988_port, QN => 
                           n_1404);
   IF_Regsxreg_file_regx2xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468404, Q => IF_Regsxreg_file_956_port, QN => 
                           n_1405);
   IF_Regsxreg_file_regx3xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468399, Q => IF_Regsxreg_file_924_port, QN => 
                           n_1406);
   IF_Regsxreg_file_regx4xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468394, Q => IF_Regsxreg_file_892_port, QN => 
                           n_1407);
   IF_Regsxreg_file_regx5xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468389, Q => IF_Regsxreg_file_860_port, QN => 
                           n_1408);
   IF_Regsxreg_file_regx6xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468384, Q => IF_Regsxreg_file_828_port, QN => 
                           n_1409);
   IF_Regsxreg_file_regx7xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468379, Q => IF_Regsxreg_file_796_port, QN => 
                           n_1410);
   IF_Regsxreg_file_regx8xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468374, Q => IF_Regsxreg_file_764_port, QN => 
                           n_1411);
   IF_Regsxreg_file_regx9xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468369, Q => IF_Regsxreg_file_732_port, QN => 
                           n_1412);
   IF_Regsxreg_file_regx10xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468364, Q => IF_Regsxreg_file_700_port, QN => 
                           n_1413);
   IF_Regsxreg_file_regx11xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468359, Q => IF_Regsxreg_file_668_port, QN => 
                           n_1414);
   IF_Regsxreg_file_regx12xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468354, Q => IF_Regsxreg_file_636_port, QN => 
                           n_1415);
   IF_Regsxreg_file_regx13xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468349, Q => IF_Regsxreg_file_604_port, QN => 
                           n_1416);
   IF_Regsxreg_file_regx14xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468344, Q => IF_Regsxreg_file_572_port, QN => 
                           n_1417);
   IF_Regsxreg_file_regx15xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468339, Q => IF_Regsxreg_file_540_port, QN => 
                           n_1418);
   IF_Regsxreg_file_regx16xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468334, Q => IF_Regsxreg_file_508_port, QN => 
                           n_1419);
   IF_Regsxreg_file_regx17xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468329, Q => IF_Regsxreg_file_476_port, QN => 
                           n_1420);
   IF_Regsxreg_file_regx18xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468324, Q => IF_Regsxreg_file_444_port, QN => 
                           n_1421);
   IF_Regsxreg_file_regx19xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468319, Q => IF_Regsxreg_file_412_port, QN => 
                           n_1422);
   IF_Regsxreg_file_regx20xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468314, Q => IF_Regsxreg_file_380_port, QN => 
                           n_1423);
   IF_Regsxreg_file_regx21xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468309, Q => IF_Regsxreg_file_348_port, QN => 
                           n_1424);
   IF_Regsxreg_file_regx22xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468304, Q => IF_Regsxreg_file_316_port, QN => 
                           n_1425);
   IF_Regsxreg_file_regx23xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468299, Q => IF_Regsxreg_file_284_port, QN => 
                           n_1426);
   IF_Regsxreg_file_regx24xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468294, Q => IF_Regsxreg_file_252_port, QN => 
                           n_1427);
   IF_Regsxreg_file_regx25xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468289, Q => IF_Regsxreg_file_220_port, QN => 
                           n_1428);
   IF_Regsxreg_file_regx26xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468284, Q => IF_Regsxreg_file_188_port, QN => 
                           n_1429);
   IF_Regsxreg_file_regx27xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468279, Q => IF_Regsxreg_file_156_port, QN => 
                           n_1430);
   IF_Regsxreg_file_regx28xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468274, Q => IF_Regsxreg_file_124_port, QN => 
                           n_1431);
   IF_Regsxreg_file_regx29xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468269, Q => IF_Regsxreg_file_92_port, QN => 
                           n_1432);
   IF_Regsxreg_file_regx30xx28x : DFF_X1 port map( D => IF_RegsxN688, CK => 
                           net2468264, Q => IF_Regsxreg_file_60_port, QN => 
                           n_1433);
   IF_RegsxRegsToCtl_port_contents2_regx28x : DFF_X1 port map( D => 
                           IF_RegsxN655, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_28_port, QN => n_1434);
   IF_CPathxRegsToCtl_data_signal_contents2_regx28x : DFF_X1 port map( D => 
                           IF_CPathxN2152, CK => net2468199, Q => n_1435, QN =>
                           n6290);
   IF_CPathxCtlToMem_port_dataIn_regx28x : DFF_X1 port map( D => n6490, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(28), QN => 
                           n_1436);
   IF_CPathxCtlToALU_port_reg2_contents_regx28x : DFF_X1 port map( D => n6635, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_28_port, QN => n_1437);
   IF_RegsxRegsToCtl_port_contents1_regx28x : DFF_X1 port map( D => 
                           IF_RegsxN623, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_28_port, QN => n_1438);
   IF_CPathxRegsToCtl_data_signal_contents1_regx28x : DFF_X1 port map( D => 
                           n6402, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_28_port, QN
                           => n6370);
   IF_CPathxCtlToALU_port_reg1_contents_regx28x : DFF_X1 port map( D => n6634, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_28_port, QN => n_1439);
   IF_ALUxALUtoCtl_port_regx29x : DFF_X1 port map( D => IF_ALUxN967, CK => 
                           net2468144, Q => ALUtoCtl_port_29_port, QN => n6285)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx29x : DFF_X1 port map( D => IF_CPathxN1889
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_29_port, QN => n_1440)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx29x : DFF_X1 port map( D => n6489, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(29), QN => 
                           n_1441);
   IF_CPathxCtlToRegs_port_dst_data_regx29x : DFF_X1 port map( D => n6574, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_29_port,
                           QN => n_1442);
   IF_Regsxreg_file_regx31xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468259, Q => IF_Regsxreg_file_29_port, QN => 
                           n_1443);
   IF_Regsxreg_file_regx1xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468409, Q => IF_Regsxreg_file_989_port, QN => 
                           n_1444);
   IF_Regsxreg_file_regx2xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468404, Q => IF_Regsxreg_file_957_port, QN => 
                           n_1445);
   IF_Regsxreg_file_regx3xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468399, Q => IF_Regsxreg_file_925_port, QN => 
                           n_1446);
   IF_Regsxreg_file_regx4xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468394, Q => IF_Regsxreg_file_893_port, QN => 
                           n_1447);
   IF_Regsxreg_file_regx5xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468389, Q => IF_Regsxreg_file_861_port, QN => 
                           n_1448);
   IF_Regsxreg_file_regx6xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468384, Q => IF_Regsxreg_file_829_port, QN => 
                           n_1449);
   IF_Regsxreg_file_regx7xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468379, Q => IF_Regsxreg_file_797_port, QN => 
                           n_1450);
   IF_Regsxreg_file_regx8xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468374, Q => IF_Regsxreg_file_765_port, QN => 
                           n_1451);
   IF_Regsxreg_file_regx9xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468369, Q => IF_Regsxreg_file_733_port, QN => 
                           n_1452);
   IF_Regsxreg_file_regx10xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468364, Q => IF_Regsxreg_file_701_port, QN => 
                           n_1453);
   IF_Regsxreg_file_regx11xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468359, Q => IF_Regsxreg_file_669_port, QN => 
                           n_1454);
   IF_Regsxreg_file_regx12xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468354, Q => IF_Regsxreg_file_637_port, QN => 
                           n_1455);
   IF_Regsxreg_file_regx13xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468349, Q => IF_Regsxreg_file_605_port, QN => 
                           n_1456);
   IF_Regsxreg_file_regx14xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468344, Q => IF_Regsxreg_file_573_port, QN => 
                           n_1457);
   IF_Regsxreg_file_regx15xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468339, Q => IF_Regsxreg_file_541_port, QN => 
                           n_1458);
   IF_Regsxreg_file_regx16xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468334, Q => IF_Regsxreg_file_509_port, QN => 
                           n_1459);
   IF_Regsxreg_file_regx17xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468329, Q => IF_Regsxreg_file_477_port, QN => 
                           n_1460);
   IF_Regsxreg_file_regx18xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468324, Q => IF_Regsxreg_file_445_port, QN => 
                           n_1461);
   IF_Regsxreg_file_regx19xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468319, Q => IF_Regsxreg_file_413_port, QN => 
                           n_1462);
   IF_Regsxreg_file_regx20xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468314, Q => IF_Regsxreg_file_381_port, QN => 
                           n_1463);
   IF_Regsxreg_file_regx21xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468309, Q => IF_Regsxreg_file_349_port, QN => 
                           n_1464);
   IF_Regsxreg_file_regx22xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468304, Q => IF_Regsxreg_file_317_port, QN => 
                           n_1465);
   IF_Regsxreg_file_regx23xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468299, Q => IF_Regsxreg_file_285_port, QN => 
                           n_1466);
   IF_Regsxreg_file_regx24xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468294, Q => IF_Regsxreg_file_253_port, QN => 
                           n_1467);
   IF_Regsxreg_file_regx25xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468289, Q => IF_Regsxreg_file_221_port, QN => 
                           n_1468);
   IF_Regsxreg_file_regx26xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468284, Q => IF_Regsxreg_file_189_port, QN => 
                           n_1469);
   IF_Regsxreg_file_regx27xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468279, Q => IF_Regsxreg_file_157_port, QN => 
                           n_1470);
   IF_Regsxreg_file_regx28xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468274, Q => IF_Regsxreg_file_125_port, QN => 
                           n_1471);
   IF_Regsxreg_file_regx29xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468269, Q => IF_Regsxreg_file_93_port, QN => 
                           n_1472);
   IF_Regsxreg_file_regx30xx29x : DFF_X1 port map( D => IF_RegsxN689, CK => 
                           net2468264, Q => IF_Regsxreg_file_61_port, QN => 
                           n_1473);
   IF_RegsxRegsToCtl_port_contents2_regx29x : DFF_X1 port map( D => 
                           IF_RegsxN656, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_29_port, QN => n_1474);
   IF_CPathxRegsToCtl_data_signal_contents2_regx29x : DFF_X1 port map( D => 
                           IF_CPathxN2153, CK => net2468199, Q => n_1475, QN =>
                           n6291);
   IF_CPathxCtlToMem_port_dataIn_regx29x : DFF_X1 port map( D => n6488, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(29), QN => 
                           n_1476);
   IF_CPathxCtlToALU_port_reg2_contents_regx29x : DFF_X1 port map( D => n6633, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_29_port, QN => n_1477);
   IF_RegsxRegsToCtl_port_contents1_regx29x : DFF_X1 port map( D => 
                           IF_RegsxN624, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_29_port, QN => n_1478);
   IF_CPathxRegsToCtl_data_signal_contents1_regx29x : DFF_X1 port map( D => 
                           n6403, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_29_port, QN
                           => n6371);
   IF_CPathxCtlToALU_port_reg1_contents_regx29x : DFF_X1 port map( D => n6632, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_29_port, QN => n_1479);
   IF_ALUxALUtoCtl_port_regx10x : DFF_X1 port map( D => IF_ALUxN948, CK => 
                           net2468144, Q => ALUtoCtl_port_10_port, QN => n6275)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx10x : DFF_X1 port map( D => IF_CPathxN1870
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_10_port, QN => n_1480)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx10x : DFF_X1 port map( D => n6487, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(10), QN => 
                           n_1481);
   IF_CPathxCtlToRegs_port_dst_data_regx10x : DFF_X1 port map( D => n6573, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_10_port,
                           QN => n_1482);
   IF_Regsxreg_file_regx31xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468259, Q => IF_Regsxreg_file_10_port, QN => 
                           n_1483);
   IF_Regsxreg_file_regx1xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468409, Q => IF_Regsxreg_file_970_port, QN => 
                           n_1484);
   IF_Regsxreg_file_regx2xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468404, Q => IF_Regsxreg_file_938_port, QN => 
                           n_1485);
   IF_Regsxreg_file_regx3xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468399, Q => IF_Regsxreg_file_906_port, QN => 
                           n_1486);
   IF_Regsxreg_file_regx4xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468394, Q => IF_Regsxreg_file_874_port, QN => 
                           n_1487);
   IF_Regsxreg_file_regx5xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468389, Q => IF_Regsxreg_file_842_port, QN => 
                           n_1488);
   IF_Regsxreg_file_regx6xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468384, Q => IF_Regsxreg_file_810_port, QN => 
                           n_1489);
   IF_Regsxreg_file_regx7xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468379, Q => IF_Regsxreg_file_778_port, QN => 
                           n_1490);
   IF_Regsxreg_file_regx8xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468374, Q => IF_Regsxreg_file_746_port, QN => 
                           n_1491);
   IF_Regsxreg_file_regx9xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468369, Q => IF_Regsxreg_file_714_port, QN => 
                           n_1492);
   IF_Regsxreg_file_regx10xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468364, Q => IF_Regsxreg_file_682_port, QN => 
                           n_1493);
   IF_Regsxreg_file_regx11xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468359, Q => IF_Regsxreg_file_650_port, QN => 
                           n_1494);
   IF_Regsxreg_file_regx12xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468354, Q => IF_Regsxreg_file_618_port, QN => 
                           n_1495);
   IF_Regsxreg_file_regx13xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468349, Q => IF_Regsxreg_file_586_port, QN => 
                           n_1496);
   IF_Regsxreg_file_regx14xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468344, Q => IF_Regsxreg_file_554_port, QN => 
                           n_1497);
   IF_Regsxreg_file_regx15xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468339, Q => IF_Regsxreg_file_522_port, QN => 
                           n_1498);
   IF_Regsxreg_file_regx16xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468334, Q => IF_Regsxreg_file_490_port, QN => 
                           n_1499);
   IF_Regsxreg_file_regx17xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468329, Q => IF_Regsxreg_file_458_port, QN => 
                           n_1500);
   IF_Regsxreg_file_regx18xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468324, Q => IF_Regsxreg_file_426_port, QN => 
                           n_1501);
   IF_Regsxreg_file_regx19xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468319, Q => IF_Regsxreg_file_394_port, QN => 
                           n_1502);
   IF_Regsxreg_file_regx20xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468314, Q => IF_Regsxreg_file_362_port, QN => 
                           n_1503);
   IF_Regsxreg_file_regx21xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468309, Q => IF_Regsxreg_file_330_port, QN => 
                           n_1504);
   IF_Regsxreg_file_regx22xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468304, Q => IF_Regsxreg_file_298_port, QN => 
                           n_1505);
   IF_Regsxreg_file_regx23xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468299, Q => IF_Regsxreg_file_266_port, QN => 
                           n_1506);
   IF_Regsxreg_file_regx24xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468294, Q => IF_Regsxreg_file_234_port, QN => 
                           n_1507);
   IF_Regsxreg_file_regx25xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468289, Q => IF_Regsxreg_file_202_port, QN => 
                           n_1508);
   IF_Regsxreg_file_regx26xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468284, Q => IF_Regsxreg_file_170_port, QN => 
                           n_1509);
   IF_Regsxreg_file_regx27xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468279, Q => IF_Regsxreg_file_138_port, QN => 
                           n_1510);
   IF_Regsxreg_file_regx28xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468274, Q => IF_Regsxreg_file_106_port, QN => 
                           n_1511);
   IF_Regsxreg_file_regx29xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468269, Q => IF_Regsxreg_file_74_port, QN => 
                           n_1512);
   IF_Regsxreg_file_regx30xx10x : DFF_X1 port map( D => IF_RegsxN670, CK => 
                           net2468264, Q => IF_Regsxreg_file_42_port, QN => 
                           n_1513);
   IF_RegsxRegsToCtl_port_contents2_regx10x : DFF_X1 port map( D => 
                           IF_RegsxN637, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_10_port, QN => n_1514);
   IF_CPathxRegsToCtl_data_signal_contents2_regx10x : DFF_X1 port map( D => 
                           IF_CPathxN2134, CK => net2468199, Q => n_1515, QN =>
                           n6292);
   IF_CPathxCtlToMem_port_dataIn_regx10x : DFF_X1 port map( D => n6486, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(10), QN => 
                           n_1516);
   IF_CPathxCtlToALU_port_reg2_contents_regx10x : DFF_X1 port map( D => n6631, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_10_port, QN => n_1517);
   IF_RegsxRegsToCtl_port_contents1_regx10x : DFF_X1 port map( D => 
                           IF_RegsxN605, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_10_port, QN => n_1518);
   IF_CPathxRegsToCtl_data_signal_contents1_regx10x : DFF_X1 port map( D => 
                           n6384, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_10_port, QN
                           => n6364);
   IF_CPathxCtlToALU_port_reg1_contents_regx10x : DFF_X1 port map( D => n6630, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_10_port, QN => n_1519);
   IF_ALUxALUtoCtl_port_regx26x : DFF_X1 port map( D => IF_ALUxN964, CK => 
                           net2468144, Q => ALUtoCtl_port_26_port, QN => n_1520
                           );
   IF_CPathxALUtoCtl_data_signal_regx26x : DFF_X1 port map( D => IF_CPathxN1886
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_26_port, QN => n_1521)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx26x : DFF_X1 port map( D => n6485, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(26), QN => 
                           n_1522);
   IF_CPathxCtlToRegs_port_dst_data_regx26x : DFF_X1 port map( D => n6572, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_26_port,
                           QN => n_1523);
   IF_Regsxreg_file_regx31xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468259, Q => IF_Regsxreg_file_26_port, QN => 
                           n_1524);
   IF_Regsxreg_file_regx1xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468409, Q => IF_Regsxreg_file_986_port, QN => 
                           n_1525);
   IF_Regsxreg_file_regx2xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468404, Q => IF_Regsxreg_file_954_port, QN => 
                           n_1526);
   IF_Regsxreg_file_regx3xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468399, Q => IF_Regsxreg_file_922_port, QN => 
                           n_1527);
   IF_Regsxreg_file_regx4xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468394, Q => IF_Regsxreg_file_890_port, QN => 
                           n_1528);
   IF_Regsxreg_file_regx5xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468389, Q => IF_Regsxreg_file_858_port, QN => 
                           n_1529);
   IF_Regsxreg_file_regx6xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468384, Q => IF_Regsxreg_file_826_port, QN => 
                           n_1530);
   IF_Regsxreg_file_regx7xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468379, Q => IF_Regsxreg_file_794_port, QN => 
                           n_1531);
   IF_Regsxreg_file_regx8xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468374, Q => IF_Regsxreg_file_762_port, QN => 
                           n_1532);
   IF_Regsxreg_file_regx9xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468369, Q => IF_Regsxreg_file_730_port, QN => 
                           n_1533);
   IF_Regsxreg_file_regx10xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468364, Q => IF_Regsxreg_file_698_port, QN => 
                           n_1534);
   IF_Regsxreg_file_regx11xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468359, Q => IF_Regsxreg_file_666_port, QN => 
                           n_1535);
   IF_Regsxreg_file_regx12xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468354, Q => IF_Regsxreg_file_634_port, QN => 
                           n_1536);
   IF_Regsxreg_file_regx13xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468349, Q => IF_Regsxreg_file_602_port, QN => 
                           n_1537);
   IF_Regsxreg_file_regx14xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468344, Q => IF_Regsxreg_file_570_port, QN => 
                           n_1538);
   IF_Regsxreg_file_regx15xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468339, Q => IF_Regsxreg_file_538_port, QN => 
                           n_1539);
   IF_Regsxreg_file_regx16xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468334, Q => IF_Regsxreg_file_506_port, QN => 
                           n_1540);
   IF_Regsxreg_file_regx17xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468329, Q => IF_Regsxreg_file_474_port, QN => 
                           n_1541);
   IF_Regsxreg_file_regx18xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468324, Q => IF_Regsxreg_file_442_port, QN => 
                           n_1542);
   IF_Regsxreg_file_regx19xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468319, Q => IF_Regsxreg_file_410_port, QN => 
                           n_1543);
   IF_Regsxreg_file_regx20xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468314, Q => IF_Regsxreg_file_378_port, QN => 
                           n_1544);
   IF_Regsxreg_file_regx21xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468309, Q => IF_Regsxreg_file_346_port, QN => 
                           n_1545);
   IF_Regsxreg_file_regx22xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468304, Q => IF_Regsxreg_file_314_port, QN => 
                           n_1546);
   IF_Regsxreg_file_regx23xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468299, Q => IF_Regsxreg_file_282_port, QN => 
                           n_1547);
   IF_Regsxreg_file_regx24xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468294, Q => IF_Regsxreg_file_250_port, QN => 
                           n_1548);
   IF_Regsxreg_file_regx25xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468289, Q => IF_Regsxreg_file_218_port, QN => 
                           n_1549);
   IF_Regsxreg_file_regx26xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468284, Q => IF_Regsxreg_file_186_port, QN => 
                           n_1550);
   IF_Regsxreg_file_regx27xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468279, Q => IF_Regsxreg_file_154_port, QN => 
                           n_1551);
   IF_Regsxreg_file_regx28xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468274, Q => IF_Regsxreg_file_122_port, QN => 
                           n_1552);
   IF_Regsxreg_file_regx29xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468269, Q => IF_Regsxreg_file_90_port, QN => 
                           n_1553);
   IF_Regsxreg_file_regx30xx26x : DFF_X1 port map( D => IF_RegsxN686, CK => 
                           net2468264, Q => IF_Regsxreg_file_58_port, QN => 
                           n_1554);
   IF_RegsxRegsToCtl_port_contents2_regx26x : DFF_X1 port map( D => 
                           IF_RegsxN653, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_26_port, QN => n_1555);
   IF_CPathxRegsToCtl_data_signal_contents2_regx26x : DFF_X1 port map( D => 
                           IF_CPathxN2150, CK => net2468199, Q => n_1556, QN =>
                           n6293);
   IF_CPathxCtlToMem_port_dataIn_regx26x : DFF_X1 port map( D => n6484, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(26), QN => 
                           n_1557);
   IF_CPathxCtlToALU_port_reg2_contents_regx26x : DFF_X1 port map( D => n6629, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_26_port, QN => n_1558);
   IF_RegsxRegsToCtl_port_contents1_regx26x : DFF_X1 port map( D => 
                           IF_RegsxN621, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_26_port, QN => n_1559);
   IF_CPathxRegsToCtl_data_signal_contents1_regx26x : DFF_X1 port map( D => 
                           n6400, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_26_port, QN
                           => n6348);
   IF_CPathxCtlToALU_port_reg1_contents_regx26x : DFF_X1 port map( D => n6628, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_26_port, QN => n_1560);
   IF_ALUxALUtoCtl_port_regx27x : DFF_X1 port map( D => IF_ALUxN965, CK => 
                           net2468144, Q => ALUtoCtl_port_27_port, QN => n6283)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx27x : DFF_X1 port map( D => IF_CPathxN1887
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_27_port, QN => n_1561)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx27x : DFF_X1 port map( D => n6483, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(27), QN => 
                           n_1562);
   IF_CPathxCtlToRegs_port_dst_data_regx27x : DFF_X1 port map( D => n6571, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_27_port,
                           QN => n_1563);
   IF_Regsxreg_file_regx31xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468259, Q => IF_Regsxreg_file_27_port, QN => 
                           n_1564);
   IF_Regsxreg_file_regx1xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468409, Q => IF_Regsxreg_file_987_port, QN => 
                           n_1565);
   IF_Regsxreg_file_regx2xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468404, Q => IF_Regsxreg_file_955_port, QN => 
                           n_1566);
   IF_Regsxreg_file_regx3xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468399, Q => IF_Regsxreg_file_923_port, QN => 
                           n_1567);
   IF_Regsxreg_file_regx4xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468394, Q => IF_Regsxreg_file_891_port, QN => 
                           n_1568);
   IF_Regsxreg_file_regx5xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468389, Q => IF_Regsxreg_file_859_port, QN => 
                           n_1569);
   IF_Regsxreg_file_regx6xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468384, Q => IF_Regsxreg_file_827_port, QN => 
                           n_1570);
   IF_Regsxreg_file_regx7xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468379, Q => IF_Regsxreg_file_795_port, QN => 
                           n_1571);
   IF_Regsxreg_file_regx8xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468374, Q => IF_Regsxreg_file_763_port, QN => 
                           n_1572);
   IF_Regsxreg_file_regx9xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468369, Q => IF_Regsxreg_file_731_port, QN => 
                           n_1573);
   IF_Regsxreg_file_regx10xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468364, Q => IF_Regsxreg_file_699_port, QN => 
                           n_1574);
   IF_Regsxreg_file_regx11xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468359, Q => IF_Regsxreg_file_667_port, QN => 
                           n_1575);
   IF_Regsxreg_file_regx12xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468354, Q => IF_Regsxreg_file_635_port, QN => 
                           n_1576);
   IF_Regsxreg_file_regx13xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468349, Q => IF_Regsxreg_file_603_port, QN => 
                           n_1577);
   IF_Regsxreg_file_regx14xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468344, Q => IF_Regsxreg_file_571_port, QN => 
                           n_1578);
   IF_Regsxreg_file_regx15xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468339, Q => IF_Regsxreg_file_539_port, QN => 
                           n_1579);
   IF_Regsxreg_file_regx16xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468334, Q => IF_Regsxreg_file_507_port, QN => 
                           n_1580);
   IF_Regsxreg_file_regx17xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468329, Q => IF_Regsxreg_file_475_port, QN => 
                           n_1581);
   IF_Regsxreg_file_regx18xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468324, Q => IF_Regsxreg_file_443_port, QN => 
                           n_1582);
   IF_Regsxreg_file_regx19xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468319, Q => IF_Regsxreg_file_411_port, QN => 
                           n_1583);
   IF_Regsxreg_file_regx20xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468314, Q => IF_Regsxreg_file_379_port, QN => 
                           n_1584);
   IF_Regsxreg_file_regx21xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468309, Q => IF_Regsxreg_file_347_port, QN => 
                           n_1585);
   IF_Regsxreg_file_regx22xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468304, Q => IF_Regsxreg_file_315_port, QN => 
                           n_1586);
   IF_Regsxreg_file_regx23xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468299, Q => IF_Regsxreg_file_283_port, QN => 
                           n_1587);
   IF_Regsxreg_file_regx24xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468294, Q => IF_Regsxreg_file_251_port, QN => 
                           n_1588);
   IF_Regsxreg_file_regx25xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468289, Q => IF_Regsxreg_file_219_port, QN => 
                           n_1589);
   IF_Regsxreg_file_regx26xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468284, Q => IF_Regsxreg_file_187_port, QN => 
                           n_1590);
   IF_Regsxreg_file_regx27xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468279, Q => IF_Regsxreg_file_155_port, QN => 
                           n_1591);
   IF_Regsxreg_file_regx28xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468274, Q => IF_Regsxreg_file_123_port, QN => 
                           n_1592);
   IF_Regsxreg_file_regx29xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468269, Q => IF_Regsxreg_file_91_port, QN => 
                           n_1593);
   IF_Regsxreg_file_regx30xx27x : DFF_X1 port map( D => IF_RegsxN687, CK => 
                           net2468264, Q => IF_Regsxreg_file_59_port, QN => 
                           n_1594);
   IF_RegsxRegsToCtl_port_contents2_regx27x : DFF_X1 port map( D => 
                           IF_RegsxN654, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_27_port, QN => n_1595);
   IF_CPathxRegsToCtl_data_signal_contents2_regx27x : DFF_X1 port map( D => 
                           IF_CPathxN2151, CK => net2468199, Q => n_1596, QN =>
                           n6294);
   IF_CPathxCtlToMem_port_dataIn_regx27x : DFF_X1 port map( D => n6482, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(27), QN => 
                           n_1597);
   IF_CPathxCtlToALU_port_reg2_contents_regx27x : DFF_X1 port map( D => n6627, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_27_port, QN => n_1598);
   IF_RegsxRegsToCtl_port_contents1_regx27x : DFF_X1 port map( D => 
                           IF_RegsxN622, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_27_port, QN => n_1599);
   IF_CPathxRegsToCtl_data_signal_contents1_regx27x : DFF_X1 port map( D => 
                           n6401, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_27_port, QN
                           => n6347);
   IF_CPathxCtlToALU_port_reg1_contents_regx27x : DFF_X1 port map( D => n6626, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_27_port, QN => n_1600);
   IF_ALUxALUtoCtl_port_regx12x : DFF_X1 port map( D => IF_ALUxN950, CK => 
                           net2468144, Q => ALUtoCtl_port_12_port, QN => n_1601
                           );
   IF_CPathxALUtoCtl_data_signal_regx12x : DFF_X1 port map( D => IF_CPathxN1872
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_12_port, QN => n_1602)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx12x : DFF_X1 port map( D => n6481, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(12), QN => 
                           n_1603);
   IF_CPathxCtlToRegs_port_dst_data_regx12x : DFF_X1 port map( D => n6570, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_12_port,
                           QN => n_1604);
   IF_Regsxreg_file_regx31xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468259, Q => IF_Regsxreg_file_12_port, QN => 
                           n_1605);
   IF_Regsxreg_file_regx1xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468409, Q => IF_Regsxreg_file_972_port, QN => 
                           n_1606);
   IF_Regsxreg_file_regx2xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468404, Q => IF_Regsxreg_file_940_port, QN => 
                           n_1607);
   IF_Regsxreg_file_regx3xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468399, Q => IF_Regsxreg_file_908_port, QN => 
                           n_1608);
   IF_Regsxreg_file_regx4xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468394, Q => IF_Regsxreg_file_876_port, QN => 
                           n_1609);
   IF_Regsxreg_file_regx5xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468389, Q => IF_Regsxreg_file_844_port, QN => 
                           n_1610);
   IF_Regsxreg_file_regx6xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468384, Q => IF_Regsxreg_file_812_port, QN => 
                           n_1611);
   IF_Regsxreg_file_regx7xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468379, Q => IF_Regsxreg_file_780_port, QN => 
                           n_1612);
   IF_Regsxreg_file_regx8xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468374, Q => IF_Regsxreg_file_748_port, QN => 
                           n_1613);
   IF_Regsxreg_file_regx9xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468369, Q => IF_Regsxreg_file_716_port, QN => 
                           n_1614);
   IF_Regsxreg_file_regx10xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468364, Q => IF_Regsxreg_file_684_port, QN => 
                           n_1615);
   IF_Regsxreg_file_regx11xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468359, Q => IF_Regsxreg_file_652_port, QN => 
                           n_1616);
   IF_Regsxreg_file_regx12xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468354, Q => IF_Regsxreg_file_620_port, QN => 
                           n_1617);
   IF_Regsxreg_file_regx13xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468349, Q => IF_Regsxreg_file_588_port, QN => 
                           n_1618);
   IF_Regsxreg_file_regx14xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468344, Q => IF_Regsxreg_file_556_port, QN => 
                           n_1619);
   IF_Regsxreg_file_regx15xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468339, Q => IF_Regsxreg_file_524_port, QN => 
                           n_1620);
   IF_Regsxreg_file_regx16xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468334, Q => IF_Regsxreg_file_492_port, QN => 
                           n_1621);
   IF_Regsxreg_file_regx17xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468329, Q => IF_Regsxreg_file_460_port, QN => 
                           n_1622);
   IF_Regsxreg_file_regx18xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468324, Q => IF_Regsxreg_file_428_port, QN => 
                           n_1623);
   IF_Regsxreg_file_regx19xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468319, Q => IF_Regsxreg_file_396_port, QN => 
                           n_1624);
   IF_Regsxreg_file_regx20xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468314, Q => IF_Regsxreg_file_364_port, QN => 
                           n_1625);
   IF_Regsxreg_file_regx21xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468309, Q => IF_Regsxreg_file_332_port, QN => 
                           n_1626);
   IF_Regsxreg_file_regx22xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468304, Q => IF_Regsxreg_file_300_port, QN => 
                           n_1627);
   IF_Regsxreg_file_regx23xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468299, Q => IF_Regsxreg_file_268_port, QN => 
                           n_1628);
   IF_Regsxreg_file_regx24xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468294, Q => IF_Regsxreg_file_236_port, QN => 
                           n_1629);
   IF_Regsxreg_file_regx25xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468289, Q => IF_Regsxreg_file_204_port, QN => 
                           n_1630);
   IF_Regsxreg_file_regx26xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468284, Q => IF_Regsxreg_file_172_port, QN => 
                           n_1631);
   IF_Regsxreg_file_regx27xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468279, Q => IF_Regsxreg_file_140_port, QN => 
                           n_1632);
   IF_Regsxreg_file_regx28xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468274, Q => IF_Regsxreg_file_108_port, QN => 
                           n_1633);
   IF_Regsxreg_file_regx29xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468269, Q => IF_Regsxreg_file_76_port, QN => 
                           n_1634);
   IF_Regsxreg_file_regx30xx12x : DFF_X1 port map( D => IF_RegsxN672, CK => 
                           net2468264, Q => IF_Regsxreg_file_44_port, QN => 
                           n_1635);
   IF_RegsxRegsToCtl_port_contents2_regx12x : DFF_X1 port map( D => 
                           IF_RegsxN639, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_12_port, QN => n_1636);
   IF_CPathxRegsToCtl_data_signal_contents2_regx12x : DFF_X1 port map( D => 
                           IF_CPathxN2136, CK => net2468199, Q => n_1637, QN =>
                           n6295);
   IF_CPathxCtlToMem_port_dataIn_regx12x : DFF_X1 port map( D => n6480, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(12), QN => 
                           n_1638);
   IF_CPathxCtlToALU_port_reg2_contents_regx12x : DFF_X1 port map( D => n6625, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_12_port, QN => n_1639);
   IF_RegsxRegsToCtl_port_contents1_regx12x : DFF_X1 port map( D => 
                           IF_RegsxN607, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_12_port, QN => n_1640);
   IF_CPathxRegsToCtl_data_signal_contents1_regx12x : DFF_X1 port map( D => 
                           n6386, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_12_port, QN
                           => n6357);
   IF_CPathxCtlToALU_port_reg1_contents_regx12x : DFF_X1 port map( D => n6624, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_12_port, QN => n_1641);
   IF_ALUxALUtoCtl_port_regx20x : DFF_X1 port map( D => IF_ALUxN958, CK => 
                           net2468144, Q => ALUtoCtl_port_20_port, QN => n_1642
                           );
   IF_CPathxALUtoCtl_data_signal_regx20x : DFF_X1 port map( D => IF_CPathxN1880
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_20_port, QN => n_1643)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx20x : DFF_X1 port map( D => n6479, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(20), QN => 
                           n_1644);
   IF_CPathxCtlToRegs_port_dst_data_regx20x : DFF_X1 port map( D => n6569, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_20_port,
                           QN => n_1645);
   IF_Regsxreg_file_regx31xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468259, Q => IF_Regsxreg_file_20_port, QN => 
                           n_1646);
   IF_Regsxreg_file_regx1xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468409, Q => IF_Regsxreg_file_980_port, QN => 
                           n_1647);
   IF_Regsxreg_file_regx2xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468404, Q => IF_Regsxreg_file_948_port, QN => 
                           n_1648);
   IF_Regsxreg_file_regx3xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468399, Q => IF_Regsxreg_file_916_port, QN => 
                           n_1649);
   IF_Regsxreg_file_regx4xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468394, Q => IF_Regsxreg_file_884_port, QN => 
                           n_1650);
   IF_Regsxreg_file_regx5xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468389, Q => IF_Regsxreg_file_852_port, QN => 
                           n_1651);
   IF_Regsxreg_file_regx6xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468384, Q => IF_Regsxreg_file_820_port, QN => 
                           n_1652);
   IF_Regsxreg_file_regx7xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468379, Q => IF_Regsxreg_file_788_port, QN => 
                           n_1653);
   IF_Regsxreg_file_regx8xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468374, Q => IF_Regsxreg_file_756_port, QN => 
                           n_1654);
   IF_Regsxreg_file_regx9xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468369, Q => IF_Regsxreg_file_724_port, QN => 
                           n_1655);
   IF_Regsxreg_file_regx10xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468364, Q => IF_Regsxreg_file_692_port, QN => 
                           n_1656);
   IF_Regsxreg_file_regx11xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468359, Q => IF_Regsxreg_file_660_port, QN => 
                           n_1657);
   IF_Regsxreg_file_regx12xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468354, Q => IF_Regsxreg_file_628_port, QN => 
                           n_1658);
   IF_Regsxreg_file_regx13xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468349, Q => IF_Regsxreg_file_596_port, QN => 
                           n_1659);
   IF_Regsxreg_file_regx14xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468344, Q => IF_Regsxreg_file_564_port, QN => 
                           n_1660);
   IF_Regsxreg_file_regx15xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468339, Q => IF_Regsxreg_file_532_port, QN => 
                           n_1661);
   IF_Regsxreg_file_regx16xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468334, Q => IF_Regsxreg_file_500_port, QN => 
                           n_1662);
   IF_Regsxreg_file_regx17xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468329, Q => IF_Regsxreg_file_468_port, QN => 
                           n_1663);
   IF_Regsxreg_file_regx18xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468324, Q => IF_Regsxreg_file_436_port, QN => 
                           n_1664);
   IF_Regsxreg_file_regx19xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468319, Q => IF_Regsxreg_file_404_port, QN => 
                           n_1665);
   IF_Regsxreg_file_regx20xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468314, Q => IF_Regsxreg_file_372_port, QN => 
                           n_1666);
   IF_Regsxreg_file_regx21xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468309, Q => IF_Regsxreg_file_340_port, QN => 
                           n_1667);
   IF_Regsxreg_file_regx22xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468304, Q => IF_Regsxreg_file_308_port, QN => 
                           n_1668);
   IF_Regsxreg_file_regx23xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468299, Q => IF_Regsxreg_file_276_port, QN => 
                           n_1669);
   IF_Regsxreg_file_regx24xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468294, Q => IF_Regsxreg_file_244_port, QN => 
                           n_1670);
   IF_Regsxreg_file_regx25xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468289, Q => IF_Regsxreg_file_212_port, QN => 
                           n_1671);
   IF_Regsxreg_file_regx26xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468284, Q => IF_Regsxreg_file_180_port, QN => 
                           n_1672);
   IF_Regsxreg_file_regx27xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468279, Q => IF_Regsxreg_file_148_port, QN => 
                           n_1673);
   IF_Regsxreg_file_regx28xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468274, Q => IF_Regsxreg_file_116_port, QN => 
                           n_1674);
   IF_Regsxreg_file_regx29xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468269, Q => IF_Regsxreg_file_84_port, QN => 
                           n_1675);
   IF_Regsxreg_file_regx30xx20x : DFF_X1 port map( D => IF_RegsxN680, CK => 
                           net2468264, Q => IF_Regsxreg_file_52_port, QN => 
                           n_1676);
   IF_RegsxRegsToCtl_port_contents2_regx20x : DFF_X1 port map( D => 
                           IF_RegsxN647, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_20_port, QN => n_1677);
   IF_CPathxRegsToCtl_data_signal_contents2_regx20x : DFF_X1 port map( D => 
                           IF_CPathxN2144, CK => net2468199, Q => n_1678, QN =>
                           n6296);
   IF_CPathxCtlToMem_port_dataIn_regx20x : DFF_X1 port map( D => n6478, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(20), QN => 
                           n_1679);
   IF_CPathxCtlToALU_port_reg2_contents_regx20x : DFF_X1 port map( D => n6623, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_20_port, QN => n_1680);
   IF_RegsxRegsToCtl_port_contents1_regx20x : DFF_X1 port map( D => 
                           IF_RegsxN615, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_20_port, QN => n_1681);
   IF_CPathxRegsToCtl_data_signal_contents1_regx20x : DFF_X1 port map( D => 
                           n6394, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_20_port, QN
                           => n6369);
   IF_CPathxCtlToALU_port_reg1_contents_regx20x : DFF_X1 port map( D => n6622, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_20_port, QN => n_1682);
   IF_ALUxALUtoCtl_port_regx22x : DFF_X1 port map( D => IF_ALUxN960, CK => 
                           net2468144, Q => ALUtoCtl_port_22_port, QN => n6276)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx22x : DFF_X1 port map( D => IF_CPathxN1882
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_22_port, QN => n_1683)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx22x : DFF_X1 port map( D => n6477, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(22), QN => 
                           n_1684);
   IF_CPathxCtlToRegs_port_dst_data_regx22x : DFF_X1 port map( D => n6568, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_22_port,
                           QN => n_1685);
   IF_Regsxreg_file_regx31xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468259, Q => IF_Regsxreg_file_22_port, QN => 
                           n_1686);
   IF_Regsxreg_file_regx1xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468409, Q => IF_Regsxreg_file_982_port, QN => 
                           n_1687);
   IF_Regsxreg_file_regx2xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468404, Q => IF_Regsxreg_file_950_port, QN => 
                           n_1688);
   IF_Regsxreg_file_regx3xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468399, Q => IF_Regsxreg_file_918_port, QN => 
                           n_1689);
   IF_Regsxreg_file_regx4xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468394, Q => IF_Regsxreg_file_886_port, QN => 
                           n_1690);
   IF_Regsxreg_file_regx5xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468389, Q => IF_Regsxreg_file_854_port, QN => 
                           n_1691);
   IF_Regsxreg_file_regx6xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468384, Q => IF_Regsxreg_file_822_port, QN => 
                           n_1692);
   IF_Regsxreg_file_regx7xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468379, Q => IF_Regsxreg_file_790_port, QN => 
                           n_1693);
   IF_Regsxreg_file_regx8xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468374, Q => IF_Regsxreg_file_758_port, QN => 
                           n_1694);
   IF_Regsxreg_file_regx9xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468369, Q => IF_Regsxreg_file_726_port, QN => 
                           n_1695);
   IF_Regsxreg_file_regx10xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468364, Q => IF_Regsxreg_file_694_port, QN => 
                           n_1696);
   IF_Regsxreg_file_regx11xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468359, Q => IF_Regsxreg_file_662_port, QN => 
                           n_1697);
   IF_Regsxreg_file_regx12xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468354, Q => IF_Regsxreg_file_630_port, QN => 
                           n_1698);
   IF_Regsxreg_file_regx13xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468349, Q => IF_Regsxreg_file_598_port, QN => 
                           n_1699);
   IF_Regsxreg_file_regx14xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468344, Q => IF_Regsxreg_file_566_port, QN => 
                           n_1700);
   IF_Regsxreg_file_regx15xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468339, Q => IF_Regsxreg_file_534_port, QN => 
                           n_1701);
   IF_Regsxreg_file_regx16xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468334, Q => IF_Regsxreg_file_502_port, QN => 
                           n_1702);
   IF_Regsxreg_file_regx17xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468329, Q => IF_Regsxreg_file_470_port, QN => 
                           n_1703);
   IF_Regsxreg_file_regx18xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468324, Q => IF_Regsxreg_file_438_port, QN => 
                           n_1704);
   IF_Regsxreg_file_regx19xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468319, Q => IF_Regsxreg_file_406_port, QN => 
                           n_1705);
   IF_Regsxreg_file_regx20xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468314, Q => IF_Regsxreg_file_374_port, QN => 
                           n_1706);
   IF_Regsxreg_file_regx21xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468309, Q => IF_Regsxreg_file_342_port, QN => 
                           n_1707);
   IF_Regsxreg_file_regx22xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468304, Q => IF_Regsxreg_file_310_port, QN => 
                           n_1708);
   IF_Regsxreg_file_regx23xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468299, Q => IF_Regsxreg_file_278_port, QN => 
                           n_1709);
   IF_Regsxreg_file_regx24xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468294, Q => IF_Regsxreg_file_246_port, QN => 
                           n_1710);
   IF_Regsxreg_file_regx25xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468289, Q => IF_Regsxreg_file_214_port, QN => 
                           n_1711);
   IF_Regsxreg_file_regx26xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468284, Q => IF_Regsxreg_file_182_port, QN => 
                           n_1712);
   IF_Regsxreg_file_regx27xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468279, Q => IF_Regsxreg_file_150_port, QN => 
                           n_1713);
   IF_Regsxreg_file_regx28xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468274, Q => IF_Regsxreg_file_118_port, QN => 
                           n_1714);
   IF_Regsxreg_file_regx29xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468269, Q => IF_Regsxreg_file_86_port, QN => 
                           n_1715);
   IF_Regsxreg_file_regx30xx22x : DFF_X1 port map( D => IF_RegsxN682, CK => 
                           net2468264, Q => IF_Regsxreg_file_54_port, QN => 
                           n_1716);
   IF_RegsxRegsToCtl_port_contents2_regx22x : DFF_X1 port map( D => 
                           IF_RegsxN649, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_22_port, QN => n_1717);
   IF_CPathxRegsToCtl_data_signal_contents2_regx22x : DFF_X1 port map( D => 
                           IF_CPathxN2146, CK => net2468199, Q => n_1718, QN =>
                           n6297);
   IF_CPathxCtlToMem_port_dataIn_regx22x : DFF_X1 port map( D => n6476, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(22), QN => 
                           n_1719);
   IF_CPathxCtlToALU_port_reg2_contents_regx22x : DFF_X1 port map( D => n6621, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_22_port, QN => n_1720);
   IF_RegsxRegsToCtl_port_contents1_regx22x : DFF_X1 port map( D => 
                           IF_RegsxN617, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_22_port, QN => n_1721);
   IF_CPathxRegsToCtl_data_signal_contents1_regx22x : DFF_X1 port map( D => 
                           n6396, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_22_port, QN
                           => n6351);
   IF_CPathxCtlToALU_port_reg1_contents_regx22x : DFF_X1 port map( D => n6620, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_22_port, QN => n_1722);
   IF_ALUxALUtoCtl_port_regx23x : DFF_X1 port map( D => IF_ALUxN961, CK => 
                           net2468144, Q => ALUtoCtl_port_23_port, QN => n_1723
                           );
   IF_CPathxALUtoCtl_data_signal_regx23x : DFF_X1 port map( D => IF_CPathxN1883
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_23_port, QN => n_1724)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx23x : DFF_X1 port map( D => n6475, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(23), QN => 
                           n_1725);
   IF_CPathxCtlToRegs_port_dst_data_regx23x : DFF_X1 port map( D => n6567, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_23_port,
                           QN => n_1726);
   IF_Regsxreg_file_regx31xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468259, Q => IF_Regsxreg_file_23_port, QN => 
                           n_1727);
   IF_Regsxreg_file_regx1xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468409, Q => IF_Regsxreg_file_983_port, QN => 
                           n_1728);
   IF_Regsxreg_file_regx2xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468404, Q => IF_Regsxreg_file_951_port, QN => 
                           n_1729);
   IF_Regsxreg_file_regx3xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468399, Q => IF_Regsxreg_file_919_port, QN => 
                           n_1730);
   IF_Regsxreg_file_regx4xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468394, Q => IF_Regsxreg_file_887_port, QN => 
                           n_1731);
   IF_Regsxreg_file_regx5xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468389, Q => IF_Regsxreg_file_855_port, QN => 
                           n_1732);
   IF_Regsxreg_file_regx6xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468384, Q => IF_Regsxreg_file_823_port, QN => 
                           n_1733);
   IF_Regsxreg_file_regx7xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468379, Q => IF_Regsxreg_file_791_port, QN => 
                           n_1734);
   IF_Regsxreg_file_regx8xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468374, Q => IF_Regsxreg_file_759_port, QN => 
                           n_1735);
   IF_Regsxreg_file_regx9xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468369, Q => IF_Regsxreg_file_727_port, QN => 
                           n_1736);
   IF_Regsxreg_file_regx10xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468364, Q => IF_Regsxreg_file_695_port, QN => 
                           n_1737);
   IF_Regsxreg_file_regx11xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468359, Q => IF_Regsxreg_file_663_port, QN => 
                           n_1738);
   IF_Regsxreg_file_regx12xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468354, Q => IF_Regsxreg_file_631_port, QN => 
                           n_1739);
   IF_Regsxreg_file_regx13xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468349, Q => IF_Regsxreg_file_599_port, QN => 
                           n_1740);
   IF_Regsxreg_file_regx14xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468344, Q => IF_Regsxreg_file_567_port, QN => 
                           n_1741);
   IF_Regsxreg_file_regx15xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468339, Q => IF_Regsxreg_file_535_port, QN => 
                           n_1742);
   IF_Regsxreg_file_regx16xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468334, Q => IF_Regsxreg_file_503_port, QN => 
                           n_1743);
   IF_Regsxreg_file_regx17xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468329, Q => IF_Regsxreg_file_471_port, QN => 
                           n_1744);
   IF_Regsxreg_file_regx18xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468324, Q => IF_Regsxreg_file_439_port, QN => 
                           n_1745);
   IF_Regsxreg_file_regx19xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468319, Q => IF_Regsxreg_file_407_port, QN => 
                           n_1746);
   IF_Regsxreg_file_regx20xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468314, Q => IF_Regsxreg_file_375_port, QN => 
                           n_1747);
   IF_Regsxreg_file_regx21xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468309, Q => IF_Regsxreg_file_343_port, QN => 
                           n_1748);
   IF_Regsxreg_file_regx22xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468304, Q => IF_Regsxreg_file_311_port, QN => 
                           n_1749);
   IF_Regsxreg_file_regx23xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468299, Q => IF_Regsxreg_file_279_port, QN => 
                           n_1750);
   IF_Regsxreg_file_regx24xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468294, Q => IF_Regsxreg_file_247_port, QN => 
                           n_1751);
   IF_Regsxreg_file_regx25xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468289, Q => IF_Regsxreg_file_215_port, QN => 
                           n_1752);
   IF_Regsxreg_file_regx26xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468284, Q => IF_Regsxreg_file_183_port, QN => 
                           n_1753);
   IF_Regsxreg_file_regx27xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468279, Q => IF_Regsxreg_file_151_port, QN => 
                           n_1754);
   IF_Regsxreg_file_regx28xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468274, Q => IF_Regsxreg_file_119_port, QN => 
                           n_1755);
   IF_Regsxreg_file_regx29xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468269, Q => IF_Regsxreg_file_87_port, QN => 
                           n_1756);
   IF_Regsxreg_file_regx30xx23x : DFF_X1 port map( D => IF_RegsxN683, CK => 
                           net2468264, Q => IF_Regsxreg_file_55_port, QN => 
                           n_1757);
   IF_RegsxRegsToCtl_port_contents2_regx23x : DFF_X1 port map( D => 
                           IF_RegsxN650, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_23_port, QN => n_1758);
   IF_CPathxRegsToCtl_data_signal_contents2_regx23x : DFF_X1 port map( D => 
                           IF_CPathxN2147, CK => net2468199, Q => n_1759, QN =>
                           n6298);
   IF_CPathxCtlToMem_port_dataIn_regx23x : DFF_X1 port map( D => n6474, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(23), QN => 
                           n_1760);
   IF_CPathxCtlToALU_port_reg2_contents_regx23x : DFF_X1 port map( D => n6619, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_23_port, QN => n_1761);
   IF_RegsxRegsToCtl_port_contents1_regx23x : DFF_X1 port map( D => 
                           IF_RegsxN618, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_23_port, QN => n_1762);
   IF_CPathxRegsToCtl_data_signal_contents1_regx23x : DFF_X1 port map( D => 
                           n6397, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_23_port, QN
                           => n6350);
   IF_CPathxCtlToALU_port_reg1_contents_regx23x : DFF_X1 port map( D => n6618, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_23_port, QN => n_1763);
   IF_ALUxALUtoCtl_port_regx8x : DFF_X1 port map( D => IF_ALUxN946, CK => 
                           net2468144, Q => ALUtoCtl_port_8_port, QN => n_1764)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx8x : DFF_X1 port map( D => IF_CPathxN1868,
                           CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_8_port, QN => n_1765);
   IF_CPathxCtlToMem_port_addrIn_regx8x : DFF_X1 port map( D => n6473, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(8), QN => 
                           n_1766);
   IF_CPathxCtlToRegs_port_dst_data_regx8x : DFF_X1 port map( D => n6566, CK =>
                           net2468214, Q => CtlToRegs_port_dst_data_8_port, QN 
                           => n_1767);
   IF_Regsxreg_file_regx31xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468259, Q => IF_Regsxreg_file_8_port, QN => 
                           n_1768);
   IF_Regsxreg_file_regx1xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468409, Q => IF_Regsxreg_file_968_port, QN => 
                           n_1769);
   IF_Regsxreg_file_regx2xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468404, Q => IF_Regsxreg_file_936_port, QN => 
                           n_1770);
   IF_Regsxreg_file_regx3xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468399, Q => IF_Regsxreg_file_904_port, QN => 
                           n_1771);
   IF_Regsxreg_file_regx4xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468394, Q => IF_Regsxreg_file_872_port, QN => 
                           n_1772);
   IF_Regsxreg_file_regx5xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468389, Q => IF_Regsxreg_file_840_port, QN => 
                           n_1773);
   IF_Regsxreg_file_regx6xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468384, Q => IF_Regsxreg_file_808_port, QN => 
                           n_1774);
   IF_Regsxreg_file_regx7xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468379, Q => IF_Regsxreg_file_776_port, QN => 
                           n_1775);
   IF_Regsxreg_file_regx8xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468374, Q => IF_Regsxreg_file_744_port, QN => 
                           n_1776);
   IF_Regsxreg_file_regx9xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468369, Q => IF_Regsxreg_file_712_port, QN => 
                           n_1777);
   IF_Regsxreg_file_regx10xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468364, Q => IF_Regsxreg_file_680_port, QN => 
                           n_1778);
   IF_Regsxreg_file_regx11xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468359, Q => IF_Regsxreg_file_648_port, QN => 
                           n_1779);
   IF_Regsxreg_file_regx12xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468354, Q => IF_Regsxreg_file_616_port, QN => 
                           n_1780);
   IF_Regsxreg_file_regx13xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468349, Q => IF_Regsxreg_file_584_port, QN => 
                           n_1781);
   IF_Regsxreg_file_regx14xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468344, Q => IF_Regsxreg_file_552_port, QN => 
                           n_1782);
   IF_Regsxreg_file_regx15xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468339, Q => IF_Regsxreg_file_520_port, QN => 
                           n_1783);
   IF_Regsxreg_file_regx16xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468334, Q => IF_Regsxreg_file_488_port, QN => 
                           n_1784);
   IF_Regsxreg_file_regx17xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468329, Q => IF_Regsxreg_file_456_port, QN => 
                           n_1785);
   IF_Regsxreg_file_regx18xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468324, Q => IF_Regsxreg_file_424_port, QN => 
                           n_1786);
   IF_Regsxreg_file_regx19xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468319, Q => IF_Regsxreg_file_392_port, QN => 
                           n_1787);
   IF_Regsxreg_file_regx20xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468314, Q => IF_Regsxreg_file_360_port, QN => 
                           n_1788);
   IF_Regsxreg_file_regx21xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468309, Q => IF_Regsxreg_file_328_port, QN => 
                           n_1789);
   IF_Regsxreg_file_regx22xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468304, Q => IF_Regsxreg_file_296_port, QN => 
                           n_1790);
   IF_Regsxreg_file_regx23xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468299, Q => IF_Regsxreg_file_264_port, QN => 
                           n_1791);
   IF_Regsxreg_file_regx24xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468294, Q => IF_Regsxreg_file_232_port, QN => 
                           n_1792);
   IF_Regsxreg_file_regx25xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468289, Q => IF_Regsxreg_file_200_port, QN => 
                           n_1793);
   IF_Regsxreg_file_regx26xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468284, Q => IF_Regsxreg_file_168_port, QN => 
                           n_1794);
   IF_Regsxreg_file_regx27xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468279, Q => IF_Regsxreg_file_136_port, QN => 
                           n_1795);
   IF_Regsxreg_file_regx28xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468274, Q => IF_Regsxreg_file_104_port, QN => 
                           n_1796);
   IF_Regsxreg_file_regx29xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468269, Q => IF_Regsxreg_file_72_port, QN => 
                           n_1797);
   IF_Regsxreg_file_regx30xx8x : DFF_X1 port map( D => IF_RegsxN668, CK => 
                           net2468264, Q => IF_Regsxreg_file_40_port, QN => 
                           n_1798);
   IF_RegsxRegsToCtl_port_contents2_regx8x : DFF_X1 port map( D => IF_RegsxN635
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents2_8_port, QN => n_1799);
   IF_CPathxRegsToCtl_data_signal_contents2_regx8x : DFF_X1 port map( D => 
                           IF_CPathxN2132, CK => net2468199, Q => n_1800, QN =>
                           n6299);
   IF_CPathxCtlToMem_port_dataIn_regx8x : DFF_X1 port map( D => n6472, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(8), QN => 
                           n_1801);
   IF_CPathxCtlToALU_port_reg2_contents_regx8x : DFF_X1 port map( D => n6617, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_8_port, QN => n_1802);
   IF_RegsxRegsToCtl_port_contents1_regx8x : DFF_X1 port map( D => IF_RegsxN603
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents1_8_port, QN => n_1803);
   IF_CPathxRegsToCtl_data_signal_contents1_regx8x : DFF_X1 port map( D => 
                           n6382, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_8_port, QN 
                           => n6358);
   IF_CPathxCtlToALU_port_reg1_contents_regx8x : DFF_X1 port map( D => n6616, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_8_port, QN => n_1804);
   IF_ALUxALUtoCtl_port_regx11x : DFF_X1 port map( D => IF_ALUxN949, CK => 
                           net2468144, Q => ALUtoCtl_port_11_port, QN => n_1805
                           );
   IF_CPathxALUtoCtl_data_signal_regx11x : DFF_X1 port map( D => IF_CPathxN1871
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_11_port, QN => n_1806)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx11x : DFF_X1 port map( D => n6471, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(11), QN => 
                           n_1807);
   IF_CPathxCtlToRegs_port_dst_data_regx11x : DFF_X1 port map( D => n6565, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_11_port,
                           QN => n_1808);
   IF_Regsxreg_file_regx31xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468259, Q => IF_Regsxreg_file_11_port, QN => 
                           n_1809);
   IF_Regsxreg_file_regx1xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468409, Q => IF_Regsxreg_file_971_port, QN => 
                           n_1810);
   IF_Regsxreg_file_regx2xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468404, Q => IF_Regsxreg_file_939_port, QN => 
                           n_1811);
   IF_Regsxreg_file_regx3xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468399, Q => IF_Regsxreg_file_907_port, QN => 
                           n_1812);
   IF_Regsxreg_file_regx4xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468394, Q => IF_Regsxreg_file_875_port, QN => 
                           n_1813);
   IF_Regsxreg_file_regx5xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468389, Q => IF_Regsxreg_file_843_port, QN => 
                           n_1814);
   IF_Regsxreg_file_regx6xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468384, Q => IF_Regsxreg_file_811_port, QN => 
                           n_1815);
   IF_Regsxreg_file_regx7xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468379, Q => IF_Regsxreg_file_779_port, QN => 
                           n_1816);
   IF_Regsxreg_file_regx8xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468374, Q => IF_Regsxreg_file_747_port, QN => 
                           n_1817);
   IF_Regsxreg_file_regx9xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468369, Q => IF_Regsxreg_file_715_port, QN => 
                           n_1818);
   IF_Regsxreg_file_regx10xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468364, Q => IF_Regsxreg_file_683_port, QN => 
                           n_1819);
   IF_Regsxreg_file_regx11xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468359, Q => IF_Regsxreg_file_651_port, QN => 
                           n_1820);
   IF_Regsxreg_file_regx12xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468354, Q => IF_Regsxreg_file_619_port, QN => 
                           n_1821);
   IF_Regsxreg_file_regx13xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468349, Q => IF_Regsxreg_file_587_port, QN => 
                           n_1822);
   IF_Regsxreg_file_regx14xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468344, Q => IF_Regsxreg_file_555_port, QN => 
                           n_1823);
   IF_Regsxreg_file_regx15xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468339, Q => IF_Regsxreg_file_523_port, QN => 
                           n_1824);
   IF_Regsxreg_file_regx16xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468334, Q => IF_Regsxreg_file_491_port, QN => 
                           n_1825);
   IF_Regsxreg_file_regx17xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468329, Q => IF_Regsxreg_file_459_port, QN => 
                           n_1826);
   IF_Regsxreg_file_regx18xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468324, Q => IF_Regsxreg_file_427_port, QN => 
                           n_1827);
   IF_Regsxreg_file_regx19xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468319, Q => IF_Regsxreg_file_395_port, QN => 
                           n_1828);
   IF_Regsxreg_file_regx20xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468314, Q => IF_Regsxreg_file_363_port, QN => 
                           n_1829);
   IF_Regsxreg_file_regx21xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468309, Q => IF_Regsxreg_file_331_port, QN => 
                           n_1830);
   IF_Regsxreg_file_regx22xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468304, Q => IF_Regsxreg_file_299_port, QN => 
                           n_1831);
   IF_Regsxreg_file_regx23xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468299, Q => IF_Regsxreg_file_267_port, QN => 
                           n_1832);
   IF_Regsxreg_file_regx24xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468294, Q => IF_Regsxreg_file_235_port, QN => 
                           n_1833);
   IF_Regsxreg_file_regx25xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468289, Q => IF_Regsxreg_file_203_port, QN => 
                           n_1834);
   IF_Regsxreg_file_regx26xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468284, Q => IF_Regsxreg_file_171_port, QN => 
                           n_1835);
   IF_Regsxreg_file_regx27xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468279, Q => IF_Regsxreg_file_139_port, QN => 
                           n_1836);
   IF_Regsxreg_file_regx28xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468274, Q => IF_Regsxreg_file_107_port, QN => 
                           n_1837);
   IF_Regsxreg_file_regx29xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468269, Q => IF_Regsxreg_file_75_port, QN => 
                           n_1838);
   IF_Regsxreg_file_regx30xx11x : DFF_X1 port map( D => IF_RegsxN671, CK => 
                           net2468264, Q => IF_Regsxreg_file_43_port, QN => 
                           n_1839);
   IF_RegsxRegsToCtl_port_contents2_regx11x : DFF_X1 port map( D => 
                           IF_RegsxN638, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_11_port, QN => n_1840);
   IF_CPathxRegsToCtl_data_signal_contents2_regx11x : DFF_X1 port map( D => 
                           IF_CPathxN2135, CK => net2468199, Q => n_1841, QN =>
                           n6300);
   IF_CPathxCtlToMem_port_dataIn_regx11x : DFF_X1 port map( D => n6470, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(11), QN => 
                           n_1842);
   IF_CPathxCtlToALU_port_reg2_contents_regx11x : DFF_X1 port map( D => n6615, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_11_port, QN => n_1843);
   IF_RegsxRegsToCtl_port_contents1_regx11x : DFF_X1 port map( D => 
                           IF_RegsxN606, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_11_port, QN => n_1844);
   IF_CPathxRegsToCtl_data_signal_contents1_regx11x : DFF_X1 port map( D => 
                           n6385, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_11_port, QN
                           => n6363);
   IF_CPathxCtlToALU_port_reg1_contents_regx11x : DFF_X1 port map( D => n6614, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_11_port, QN => n_1845);
   IF_ALUxALUtoCtl_port_regx13x : DFF_X1 port map( D => IF_ALUxN951, CK => 
                           net2468144, Q => ALUtoCtl_port_13_port, QN => n6282)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx13x : DFF_X1 port map( D => IF_CPathxN1873
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_13_port, QN => n_1846)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx13x : DFF_X1 port map( D => n6469, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(13), QN => 
                           n_1847);
   IF_CPathxCtlToRegs_port_dst_data_regx13x : DFF_X1 port map( D => n6564, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_13_port,
                           QN => n_1848);
   IF_Regsxreg_file_regx31xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468259, Q => IF_Regsxreg_file_13_port, QN => 
                           n_1849);
   IF_Regsxreg_file_regx1xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468409, Q => IF_Regsxreg_file_973_port, QN => 
                           n_1850);
   IF_Regsxreg_file_regx2xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468404, Q => IF_Regsxreg_file_941_port, QN => 
                           n_1851);
   IF_Regsxreg_file_regx3xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468399, Q => IF_Regsxreg_file_909_port, QN => 
                           n_1852);
   IF_Regsxreg_file_regx4xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468394, Q => IF_Regsxreg_file_877_port, QN => 
                           n_1853);
   IF_Regsxreg_file_regx5xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468389, Q => IF_Regsxreg_file_845_port, QN => 
                           n_1854);
   IF_Regsxreg_file_regx6xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468384, Q => IF_Regsxreg_file_813_port, QN => 
                           n_1855);
   IF_Regsxreg_file_regx7xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468379, Q => IF_Regsxreg_file_781_port, QN => 
                           n_1856);
   IF_Regsxreg_file_regx8xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468374, Q => IF_Regsxreg_file_749_port, QN => 
                           n_1857);
   IF_Regsxreg_file_regx9xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468369, Q => IF_Regsxreg_file_717_port, QN => 
                           n_1858);
   IF_Regsxreg_file_regx10xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468364, Q => IF_Regsxreg_file_685_port, QN => 
                           n_1859);
   IF_Regsxreg_file_regx11xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468359, Q => IF_Regsxreg_file_653_port, QN => 
                           n_1860);
   IF_Regsxreg_file_regx12xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468354, Q => IF_Regsxreg_file_621_port, QN => 
                           n_1861);
   IF_Regsxreg_file_regx13xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468349, Q => IF_Regsxreg_file_589_port, QN => 
                           n_1862);
   IF_Regsxreg_file_regx14xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468344, Q => IF_Regsxreg_file_557_port, QN => 
                           n_1863);
   IF_Regsxreg_file_regx15xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468339, Q => IF_Regsxreg_file_525_port, QN => 
                           n_1864);
   IF_Regsxreg_file_regx16xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468334, Q => IF_Regsxreg_file_493_port, QN => 
                           n_1865);
   IF_Regsxreg_file_regx17xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468329, Q => IF_Regsxreg_file_461_port, QN => 
                           n_1866);
   IF_Regsxreg_file_regx18xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468324, Q => IF_Regsxreg_file_429_port, QN => 
                           n_1867);
   IF_Regsxreg_file_regx19xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468319, Q => IF_Regsxreg_file_397_port, QN => 
                           n_1868);
   IF_Regsxreg_file_regx20xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468314, Q => IF_Regsxreg_file_365_port, QN => 
                           n_1869);
   IF_Regsxreg_file_regx21xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468309, Q => IF_Regsxreg_file_333_port, QN => 
                           n_1870);
   IF_Regsxreg_file_regx22xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468304, Q => IF_Regsxreg_file_301_port, QN => 
                           n_1871);
   IF_Regsxreg_file_regx23xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468299, Q => IF_Regsxreg_file_269_port, QN => 
                           n_1872);
   IF_Regsxreg_file_regx24xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468294, Q => IF_Regsxreg_file_237_port, QN => 
                           n_1873);
   IF_Regsxreg_file_regx25xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468289, Q => IF_Regsxreg_file_205_port, QN => 
                           n_1874);
   IF_Regsxreg_file_regx26xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468284, Q => IF_Regsxreg_file_173_port, QN => 
                           n_1875);
   IF_Regsxreg_file_regx27xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468279, Q => IF_Regsxreg_file_141_port, QN => 
                           n_1876);
   IF_Regsxreg_file_regx28xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468274, Q => IF_Regsxreg_file_109_port, QN => 
                           n_1877);
   IF_Regsxreg_file_regx29xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468269, Q => IF_Regsxreg_file_77_port, QN => 
                           n_1878);
   IF_Regsxreg_file_regx30xx13x : DFF_X1 port map( D => IF_RegsxN673, CK => 
                           net2468264, Q => IF_Regsxreg_file_45_port, QN => 
                           n_1879);
   IF_RegsxRegsToCtl_port_contents2_regx13x : DFF_X1 port map( D => 
                           IF_RegsxN640, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_13_port, QN => n_1880);
   IF_CPathxRegsToCtl_data_signal_contents2_regx13x : DFF_X1 port map( D => 
                           IF_CPathxN2137, CK => net2468199, Q => n_1881, QN =>
                           n6301);
   IF_CPathxCtlToMem_port_dataIn_regx13x : DFF_X1 port map( D => n6468, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(13), QN => 
                           n_1882);
   IF_CPathxCtlToALU_port_reg2_contents_regx13x : DFF_X1 port map( D => n6613, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_13_port, QN => n_1883);
   IF_RegsxRegsToCtl_port_contents1_regx13x : DFF_X1 port map( D => 
                           IF_RegsxN608, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_13_port, QN => n_1884);
   IF_CPathxRegsToCtl_data_signal_contents1_regx13x : DFF_X1 port map( D => 
                           n6387, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_13_port, QN
                           => n6356);
   IF_CPathxCtlToALU_port_reg1_contents_regx13x : DFF_X1 port map( D => n6612, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_13_port, QN => n_1885);
   IF_ALUxALUtoCtl_port_regx15x : DFF_X1 port map( D => IF_ALUxN953, CK => 
                           net2468144, Q => ALUtoCtl_port_15_port, QN => n_1886
                           );
   IF_CPathxALUtoCtl_data_signal_regx15x : DFF_X1 port map( D => IF_CPathxN1875
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_15_port, QN => n_1887)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx15x : DFF_X1 port map( D => n6467, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(15), QN => 
                           n_1888);
   IF_CPathxCtlToRegs_port_dst_data_regx15x : DFF_X1 port map( D => n6563, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_15_port,
                           QN => n_1889);
   IF_Regsxreg_file_regx31xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468259, Q => IF_Regsxreg_file_15_port, QN => 
                           n_1890);
   IF_Regsxreg_file_regx1xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468409, Q => IF_Regsxreg_file_975_port, QN => 
                           n_1891);
   IF_Regsxreg_file_regx2xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468404, Q => IF_Regsxreg_file_943_port, QN => 
                           n_1892);
   IF_Regsxreg_file_regx3xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468399, Q => IF_Regsxreg_file_911_port, QN => 
                           n_1893);
   IF_Regsxreg_file_regx4xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468394, Q => IF_Regsxreg_file_879_port, QN => 
                           n_1894);
   IF_Regsxreg_file_regx5xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468389, Q => IF_Regsxreg_file_847_port, QN => 
                           n_1895);
   IF_Regsxreg_file_regx6xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468384, Q => IF_Regsxreg_file_815_port, QN => 
                           n_1896);
   IF_Regsxreg_file_regx7xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468379, Q => IF_Regsxreg_file_783_port, QN => 
                           n_1897);
   IF_Regsxreg_file_regx8xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468374, Q => IF_Regsxreg_file_751_port, QN => 
                           n_1898);
   IF_Regsxreg_file_regx9xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468369, Q => IF_Regsxreg_file_719_port, QN => 
                           n_1899);
   IF_Regsxreg_file_regx10xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468364, Q => IF_Regsxreg_file_687_port, QN => 
                           n_1900);
   IF_Regsxreg_file_regx11xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468359, Q => IF_Regsxreg_file_655_port, QN => 
                           n_1901);
   IF_Regsxreg_file_regx12xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468354, Q => IF_Regsxreg_file_623_port, QN => 
                           n_1902);
   IF_Regsxreg_file_regx13xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468349, Q => IF_Regsxreg_file_591_port, QN => 
                           n_1903);
   IF_Regsxreg_file_regx14xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468344, Q => IF_Regsxreg_file_559_port, QN => 
                           n_1904);
   IF_Regsxreg_file_regx15xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468339, Q => IF_Regsxreg_file_527_port, QN => 
                           n_1905);
   IF_Regsxreg_file_regx16xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468334, Q => IF_Regsxreg_file_495_port, QN => 
                           n_1906);
   IF_Regsxreg_file_regx17xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468329, Q => IF_Regsxreg_file_463_port, QN => 
                           n_1907);
   IF_Regsxreg_file_regx18xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468324, Q => IF_Regsxreg_file_431_port, QN => 
                           n_1908);
   IF_Regsxreg_file_regx19xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468319, Q => IF_Regsxreg_file_399_port, QN => 
                           n_1909);
   IF_Regsxreg_file_regx20xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468314, Q => IF_Regsxreg_file_367_port, QN => 
                           n_1910);
   IF_Regsxreg_file_regx21xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468309, Q => IF_Regsxreg_file_335_port, QN => 
                           n_1911);
   IF_Regsxreg_file_regx22xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468304, Q => IF_Regsxreg_file_303_port, QN => 
                           n_1912);
   IF_Regsxreg_file_regx23xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468299, Q => IF_Regsxreg_file_271_port, QN => 
                           n_1913);
   IF_Regsxreg_file_regx24xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468294, Q => IF_Regsxreg_file_239_port, QN => 
                           n_1914);
   IF_Regsxreg_file_regx25xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468289, Q => IF_Regsxreg_file_207_port, QN => 
                           n_1915);
   IF_Regsxreg_file_regx26xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468284, Q => IF_Regsxreg_file_175_port, QN => 
                           n_1916);
   IF_Regsxreg_file_regx27xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468279, Q => IF_Regsxreg_file_143_port, QN => 
                           n_1917);
   IF_Regsxreg_file_regx28xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468274, Q => IF_Regsxreg_file_111_port, QN => 
                           n_1918);
   IF_Regsxreg_file_regx29xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468269, Q => IF_Regsxreg_file_79_port, QN => 
                           n_1919);
   IF_Regsxreg_file_regx30xx15x : DFF_X1 port map( D => IF_RegsxN675, CK => 
                           net2468264, Q => IF_Regsxreg_file_47_port, QN => 
                           n_1920);
   IF_RegsxRegsToCtl_port_contents2_regx15x : DFF_X1 port map( D => 
                           IF_RegsxN642, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_15_port, QN => n_1921);
   IF_CPathxRegsToCtl_data_signal_contents2_regx15x : DFF_X1 port map( D => 
                           IF_CPathxN2139, CK => net2468199, Q => n_1922, QN =>
                           n6302);
   IF_CPathxCtlToMem_port_dataIn_regx15x : DFF_X1 port map( D => n6466, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(15), QN => 
                           n_1923);
   IF_CPathxCtlToALU_port_reg2_contents_regx15x : DFF_X1 port map( D => n6611, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_15_port, QN => n_1924);
   IF_RegsxRegsToCtl_port_contents1_regx15x : DFF_X1 port map( D => 
                           IF_RegsxN610, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_15_port, QN => n_1925);
   IF_CPathxRegsToCtl_data_signal_contents1_regx15x : DFF_X1 port map( D => 
                           n6389, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_15_port, QN
                           => n6354);
   IF_CPathxCtlToALU_port_reg1_contents_regx15x : DFF_X1 port map( D => n6610, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_15_port, QN => n_1926);
   IF_ALUxALUtoCtl_port_regx17x : DFF_X1 port map( D => IF_ALUxN955, CK => 
                           net2468144, Q => ALUtoCtl_port_17_port, QN => n_1927
                           );
   IF_CPathxALUtoCtl_data_signal_regx17x : DFF_X1 port map( D => IF_CPathxN1877
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_17_port, QN => n_1928)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx17x : DFF_X1 port map( D => n6465, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(17), QN => 
                           n_1929);
   IF_CPathxCtlToRegs_port_dst_data_regx17x : DFF_X1 port map( D => n6562, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_17_port,
                           QN => n_1930);
   IF_Regsxreg_file_regx31xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468259, Q => IF_Regsxreg_file_17_port, QN => 
                           n_1931);
   IF_Regsxreg_file_regx1xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468409, Q => IF_Regsxreg_file_977_port, QN => 
                           n_1932);
   IF_Regsxreg_file_regx2xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468404, Q => IF_Regsxreg_file_945_port, QN => 
                           n_1933);
   IF_Regsxreg_file_regx3xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468399, Q => IF_Regsxreg_file_913_port, QN => 
                           n_1934);
   IF_Regsxreg_file_regx4xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468394, Q => IF_Regsxreg_file_881_port, QN => 
                           n_1935);
   IF_Regsxreg_file_regx5xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468389, Q => IF_Regsxreg_file_849_port, QN => 
                           n_1936);
   IF_Regsxreg_file_regx6xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468384, Q => IF_Regsxreg_file_817_port, QN => 
                           n_1937);
   IF_Regsxreg_file_regx7xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468379, Q => IF_Regsxreg_file_785_port, QN => 
                           n_1938);
   IF_Regsxreg_file_regx8xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468374, Q => IF_Regsxreg_file_753_port, QN => 
                           n_1939);
   IF_Regsxreg_file_regx9xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468369, Q => IF_Regsxreg_file_721_port, QN => 
                           n_1940);
   IF_Regsxreg_file_regx10xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468364, Q => IF_Regsxreg_file_689_port, QN => 
                           n_1941);
   IF_Regsxreg_file_regx11xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468359, Q => IF_Regsxreg_file_657_port, QN => 
                           n_1942);
   IF_Regsxreg_file_regx12xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468354, Q => IF_Regsxreg_file_625_port, QN => 
                           n_1943);
   IF_Regsxreg_file_regx13xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468349, Q => IF_Regsxreg_file_593_port, QN => 
                           n_1944);
   IF_Regsxreg_file_regx14xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468344, Q => IF_Regsxreg_file_561_port, QN => 
                           n_1945);
   IF_Regsxreg_file_regx15xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468339, Q => IF_Regsxreg_file_529_port, QN => 
                           n_1946);
   IF_Regsxreg_file_regx16xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468334, Q => IF_Regsxreg_file_497_port, QN => 
                           n_1947);
   IF_Regsxreg_file_regx17xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468329, Q => IF_Regsxreg_file_465_port, QN => 
                           n_1948);
   IF_Regsxreg_file_regx18xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468324, Q => IF_Regsxreg_file_433_port, QN => 
                           n_1949);
   IF_Regsxreg_file_regx19xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468319, Q => IF_Regsxreg_file_401_port, QN => 
                           n_1950);
   IF_Regsxreg_file_regx20xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468314, Q => IF_Regsxreg_file_369_port, QN => 
                           n_1951);
   IF_Regsxreg_file_regx21xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468309, Q => IF_Regsxreg_file_337_port, QN => 
                           n_1952);
   IF_Regsxreg_file_regx22xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468304, Q => IF_Regsxreg_file_305_port, QN => 
                           n_1953);
   IF_Regsxreg_file_regx23xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468299, Q => IF_Regsxreg_file_273_port, QN => 
                           n_1954);
   IF_Regsxreg_file_regx24xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468294, Q => IF_Regsxreg_file_241_port, QN => 
                           n_1955);
   IF_Regsxreg_file_regx25xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468289, Q => IF_Regsxreg_file_209_port, QN => 
                           n_1956);
   IF_Regsxreg_file_regx26xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468284, Q => IF_Regsxreg_file_177_port, QN => 
                           n_1957);
   IF_Regsxreg_file_regx27xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468279, Q => IF_Regsxreg_file_145_port, QN => 
                           n_1958);
   IF_Regsxreg_file_regx28xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468274, Q => IF_Regsxreg_file_113_port, QN => 
                           n_1959);
   IF_Regsxreg_file_regx29xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468269, Q => IF_Regsxreg_file_81_port, QN => 
                           n_1960);
   IF_Regsxreg_file_regx30xx17x : DFF_X1 port map( D => IF_RegsxN677, CK => 
                           net2468264, Q => IF_Regsxreg_file_49_port, QN => 
                           n_1961);
   IF_RegsxRegsToCtl_port_contents2_regx17x : DFF_X1 port map( D => 
                           IF_RegsxN644, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_17_port, QN => n_1962);
   IF_CPathxRegsToCtl_data_signal_contents2_regx17x : DFF_X1 port map( D => 
                           IF_CPathxN2141, CK => net2468199, Q => n_1963, QN =>
                           n6303);
   IF_CPathxCtlToMem_port_dataIn_regx17x : DFF_X1 port map( D => n6464, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(17), QN => 
                           n_1964);
   IF_CPathxCtlToALU_port_reg2_contents_regx17x : DFF_X1 port map( D => n6609, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_17_port, QN => n_1965);
   IF_RegsxRegsToCtl_port_contents1_regx17x : DFF_X1 port map( D => 
                           IF_RegsxN612, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_17_port, QN => n_1966);
   IF_CPathxRegsToCtl_data_signal_contents1_regx17x : DFF_X1 port map( D => 
                           n6391, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_17_port, QN
                           => n6366);
   IF_CPathxCtlToALU_port_reg1_contents_regx17x : DFF_X1 port map( D => n6608, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_17_port, QN => n_1967);
   IF_ALUxALUtoCtl_port_regx19x : DFF_X1 port map( D => IF_ALUxN957, CK => 
                           net2468144, Q => ALUtoCtl_port_19_port, QN => n_1968
                           );
   IF_CPathxALUtoCtl_data_signal_regx19x : DFF_X1 port map( D => IF_CPathxN1879
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_19_port, QN => n_1969)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx19x : DFF_X1 port map( D => n6463, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(19), QN => 
                           n_1970);
   IF_CPathxCtlToRegs_port_dst_data_regx19x : DFF_X1 port map( D => n6561, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_19_port,
                           QN => n_1971);
   IF_Regsxreg_file_regx31xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468259, Q => IF_Regsxreg_file_19_port, QN => 
                           n_1972);
   IF_Regsxreg_file_regx1xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468409, Q => IF_Regsxreg_file_979_port, QN => 
                           n_1973);
   IF_Regsxreg_file_regx2xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468404, Q => IF_Regsxreg_file_947_port, QN => 
                           n_1974);
   IF_Regsxreg_file_regx3xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468399, Q => IF_Regsxreg_file_915_port, QN => 
                           n_1975);
   IF_Regsxreg_file_regx4xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468394, Q => IF_Regsxreg_file_883_port, QN => 
                           n_1976);
   IF_Regsxreg_file_regx5xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468389, Q => IF_Regsxreg_file_851_port, QN => 
                           n_1977);
   IF_Regsxreg_file_regx6xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468384, Q => IF_Regsxreg_file_819_port, QN => 
                           n_1978);
   IF_Regsxreg_file_regx7xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468379, Q => IF_Regsxreg_file_787_port, QN => 
                           n_1979);
   IF_Regsxreg_file_regx8xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468374, Q => IF_Regsxreg_file_755_port, QN => 
                           n_1980);
   IF_Regsxreg_file_regx9xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468369, Q => IF_Regsxreg_file_723_port, QN => 
                           n_1981);
   IF_Regsxreg_file_regx10xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468364, Q => IF_Regsxreg_file_691_port, QN => 
                           n_1982);
   IF_Regsxreg_file_regx11xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468359, Q => IF_Regsxreg_file_659_port, QN => 
                           n_1983);
   IF_Regsxreg_file_regx12xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468354, Q => IF_Regsxreg_file_627_port, QN => 
                           n_1984);
   IF_Regsxreg_file_regx13xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468349, Q => IF_Regsxreg_file_595_port, QN => 
                           n_1985);
   IF_Regsxreg_file_regx14xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468344, Q => IF_Regsxreg_file_563_port, QN => 
                           n_1986);
   IF_Regsxreg_file_regx15xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468339, Q => IF_Regsxreg_file_531_port, QN => 
                           n_1987);
   IF_Regsxreg_file_regx16xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468334, Q => IF_Regsxreg_file_499_port, QN => 
                           n_1988);
   IF_Regsxreg_file_regx17xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468329, Q => IF_Regsxreg_file_467_port, QN => 
                           n_1989);
   IF_Regsxreg_file_regx18xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468324, Q => IF_Regsxreg_file_435_port, QN => 
                           n_1990);
   IF_Regsxreg_file_regx19xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468319, Q => IF_Regsxreg_file_403_port, QN => 
                           n_1991);
   IF_Regsxreg_file_regx20xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468314, Q => IF_Regsxreg_file_371_port, QN => 
                           n_1992);
   IF_Regsxreg_file_regx21xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468309, Q => IF_Regsxreg_file_339_port, QN => 
                           n_1993);
   IF_Regsxreg_file_regx22xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468304, Q => IF_Regsxreg_file_307_port, QN => 
                           n_1994);
   IF_Regsxreg_file_regx23xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468299, Q => IF_Regsxreg_file_275_port, QN => 
                           n_1995);
   IF_Regsxreg_file_regx24xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468294, Q => IF_Regsxreg_file_243_port, QN => 
                           n_1996);
   IF_Regsxreg_file_regx25xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468289, Q => IF_Regsxreg_file_211_port, QN => 
                           n_1997);
   IF_Regsxreg_file_regx26xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468284, Q => IF_Regsxreg_file_179_port, QN => 
                           n_1998);
   IF_Regsxreg_file_regx27xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468279, Q => IF_Regsxreg_file_147_port, QN => 
                           n_1999);
   IF_Regsxreg_file_regx28xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468274, Q => IF_Regsxreg_file_115_port, QN => 
                           n_2000);
   IF_Regsxreg_file_regx29xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468269, Q => IF_Regsxreg_file_83_port, QN => 
                           n_2001);
   IF_Regsxreg_file_regx30xx19x : DFF_X1 port map( D => IF_RegsxN679, CK => 
                           net2468264, Q => IF_Regsxreg_file_51_port, QN => 
                           n_2002);
   IF_RegsxRegsToCtl_port_contents2_regx19x : DFF_X1 port map( D => 
                           IF_RegsxN646, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_19_port, QN => n_2003);
   IF_CPathxRegsToCtl_data_signal_contents2_regx19x : DFF_X1 port map( D => 
                           IF_CPathxN2143, CK => net2468199, Q => n_2004, QN =>
                           n6304);
   IF_CPathxCtlToMem_port_dataIn_regx19x : DFF_X1 port map( D => n6462, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(19), QN => 
                           n_2005);
   IF_CPathxCtlToALU_port_reg2_contents_regx19x : DFF_X1 port map( D => n6607, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_19_port, QN => n_2006);
   IF_RegsxRegsToCtl_port_contents1_regx19x : DFF_X1 port map( D => 
                           IF_RegsxN614, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_19_port, QN => n_2007);
   IF_CPathxRegsToCtl_data_signal_contents1_regx19x : DFF_X1 port map( D => 
                           n6393, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_19_port, QN
                           => n6367);
   IF_CPathxCtlToALU_port_reg1_contents_regx19x : DFF_X1 port map( D => n6606, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_19_port, QN => n_2008);
   IF_ALUxALUtoCtl_port_regx21x : DFF_X1 port map( D => IF_ALUxN959, CK => 
                           net2468144, Q => ALUtoCtl_port_21_port, QN => n_2009
                           );
   IF_CPathxALUtoCtl_data_signal_regx21x : DFF_X1 port map( D => IF_CPathxN1881
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_21_port, QN => n_2010)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx21x : DFF_X1 port map( D => n6461, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(21), QN => 
                           n_2011);
   IF_CPathxCtlToRegs_port_dst_data_regx21x : DFF_X1 port map( D => n6560, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_21_port,
                           QN => n_2012);
   IF_Regsxreg_file_regx31xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468259, Q => IF_Regsxreg_file_21_port, QN => 
                           n_2013);
   IF_Regsxreg_file_regx1xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468409, Q => IF_Regsxreg_file_981_port, QN => 
                           n_2014);
   IF_Regsxreg_file_regx2xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468404, Q => IF_Regsxreg_file_949_port, QN => 
                           n_2015);
   IF_Regsxreg_file_regx3xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468399, Q => IF_Regsxreg_file_917_port, QN => 
                           n_2016);
   IF_Regsxreg_file_regx4xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468394, Q => IF_Regsxreg_file_885_port, QN => 
                           n_2017);
   IF_Regsxreg_file_regx5xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468389, Q => IF_Regsxreg_file_853_port, QN => 
                           n_2018);
   IF_Regsxreg_file_regx6xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468384, Q => IF_Regsxreg_file_821_port, QN => 
                           n_2019);
   IF_Regsxreg_file_regx7xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468379, Q => IF_Regsxreg_file_789_port, QN => 
                           n_2020);
   IF_Regsxreg_file_regx8xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468374, Q => IF_Regsxreg_file_757_port, QN => 
                           n_2021);
   IF_Regsxreg_file_regx9xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468369, Q => IF_Regsxreg_file_725_port, QN => 
                           n_2022);
   IF_Regsxreg_file_regx10xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468364, Q => IF_Regsxreg_file_693_port, QN => 
                           n_2023);
   IF_Regsxreg_file_regx11xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468359, Q => IF_Regsxreg_file_661_port, QN => 
                           n_2024);
   IF_Regsxreg_file_regx12xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468354, Q => IF_Regsxreg_file_629_port, QN => 
                           n_2025);
   IF_Regsxreg_file_regx13xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468349, Q => IF_Regsxreg_file_597_port, QN => 
                           n_2026);
   IF_Regsxreg_file_regx14xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468344, Q => IF_Regsxreg_file_565_port, QN => 
                           n_2027);
   IF_Regsxreg_file_regx15xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468339, Q => IF_Regsxreg_file_533_port, QN => 
                           n_2028);
   IF_Regsxreg_file_regx16xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468334, Q => IF_Regsxreg_file_501_port, QN => 
                           n_2029);
   IF_Regsxreg_file_regx17xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468329, Q => IF_Regsxreg_file_469_port, QN => 
                           n_2030);
   IF_Regsxreg_file_regx18xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468324, Q => IF_Regsxreg_file_437_port, QN => 
                           n_2031);
   IF_Regsxreg_file_regx19xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468319, Q => IF_Regsxreg_file_405_port, QN => 
                           n_2032);
   IF_Regsxreg_file_regx20xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468314, Q => IF_Regsxreg_file_373_port, QN => 
                           n_2033);
   IF_Regsxreg_file_regx21xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468309, Q => IF_Regsxreg_file_341_port, QN => 
                           n_2034);
   IF_Regsxreg_file_regx22xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468304, Q => IF_Regsxreg_file_309_port, QN => 
                           n_2035);
   IF_Regsxreg_file_regx23xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468299, Q => IF_Regsxreg_file_277_port, QN => 
                           n_2036);
   IF_Regsxreg_file_regx24xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468294, Q => IF_Regsxreg_file_245_port, QN => 
                           n_2037);
   IF_Regsxreg_file_regx25xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468289, Q => IF_Regsxreg_file_213_port, QN => 
                           n_2038);
   IF_Regsxreg_file_regx26xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468284, Q => IF_Regsxreg_file_181_port, QN => 
                           n_2039);
   IF_Regsxreg_file_regx27xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468279, Q => IF_Regsxreg_file_149_port, QN => 
                           n_2040);
   IF_Regsxreg_file_regx28xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468274, Q => IF_Regsxreg_file_117_port, QN => 
                           n_2041);
   IF_Regsxreg_file_regx29xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468269, Q => IF_Regsxreg_file_85_port, QN => 
                           n_2042);
   IF_Regsxreg_file_regx30xx21x : DFF_X1 port map( D => IF_RegsxN681, CK => 
                           net2468264, Q => IF_Regsxreg_file_53_port, QN => 
                           n_2043);
   IF_RegsxRegsToCtl_port_contents2_regx21x : DFF_X1 port map( D => 
                           IF_RegsxN648, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_21_port, QN => n_2044);
   IF_CPathxRegsToCtl_data_signal_contents2_regx21x : DFF_X1 port map( D => 
                           IF_CPathxN2145, CK => net2468199, Q => n_2045, QN =>
                           n6305);
   IF_CPathxCtlToMem_port_dataIn_regx21x : DFF_X1 port map( D => n6460, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(21), QN => 
                           n_2046);
   IF_CPathxCtlToALU_port_reg2_contents_regx21x : DFF_X1 port map( D => n6605, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_21_port, QN => n_2047);
   IF_RegsxRegsToCtl_port_contents1_regx21x : DFF_X1 port map( D => 
                           IF_RegsxN616, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_21_port, QN => n_2048);
   IF_CPathxRegsToCtl_data_signal_contents1_regx21x : DFF_X1 port map( D => 
                           n6395, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_21_port, QN
                           => n6352);
   IF_CPathxCtlToALU_port_reg1_contents_regx21x : DFF_X1 port map( D => n6604, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_21_port, QN => n_2049);
   IF_ALUxALUtoCtl_port_regx18x : DFF_X1 port map( D => IF_ALUxN956, CK => 
                           net2468144, Q => ALUtoCtl_port_18_port, QN => n_2050
                           );
   IF_CPathxALUtoCtl_data_signal_regx18x : DFF_X1 port map( D => IF_CPathxN1878
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_18_port, QN => n_2051)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx18x : DFF_X1 port map( D => n6459, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(18), QN => 
                           n_2052);
   IF_CPathxCtlToRegs_port_dst_data_regx18x : DFF_X1 port map( D => n6559, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_18_port,
                           QN => n_2053);
   IF_Regsxreg_file_regx31xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468259, Q => IF_Regsxreg_file_18_port, QN => 
                           n_2054);
   IF_Regsxreg_file_regx1xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468409, Q => IF_Regsxreg_file_978_port, QN => 
                           n_2055);
   IF_Regsxreg_file_regx2xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468404, Q => IF_Regsxreg_file_946_port, QN => 
                           n_2056);
   IF_Regsxreg_file_regx3xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468399, Q => IF_Regsxreg_file_914_port, QN => 
                           n_2057);
   IF_Regsxreg_file_regx4xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468394, Q => IF_Regsxreg_file_882_port, QN => 
                           n_2058);
   IF_Regsxreg_file_regx5xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468389, Q => IF_Regsxreg_file_850_port, QN => 
                           n_2059);
   IF_Regsxreg_file_regx6xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468384, Q => IF_Regsxreg_file_818_port, QN => 
                           n_2060);
   IF_Regsxreg_file_regx7xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468379, Q => IF_Regsxreg_file_786_port, QN => 
                           n_2061);
   IF_Regsxreg_file_regx8xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468374, Q => IF_Regsxreg_file_754_port, QN => 
                           n_2062);
   IF_Regsxreg_file_regx9xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468369, Q => IF_Regsxreg_file_722_port, QN => 
                           n_2063);
   IF_Regsxreg_file_regx10xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468364, Q => IF_Regsxreg_file_690_port, QN => 
                           n_2064);
   IF_Regsxreg_file_regx11xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468359, Q => IF_Regsxreg_file_658_port, QN => 
                           n_2065);
   IF_Regsxreg_file_regx12xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468354, Q => IF_Regsxreg_file_626_port, QN => 
                           n_2066);
   IF_Regsxreg_file_regx13xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468349, Q => IF_Regsxreg_file_594_port, QN => 
                           n_2067);
   IF_Regsxreg_file_regx14xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468344, Q => IF_Regsxreg_file_562_port, QN => 
                           n_2068);
   IF_Regsxreg_file_regx15xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468339, Q => IF_Regsxreg_file_530_port, QN => 
                           n_2069);
   IF_Regsxreg_file_regx16xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468334, Q => IF_Regsxreg_file_498_port, QN => 
                           n_2070);
   IF_Regsxreg_file_regx17xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468329, Q => IF_Regsxreg_file_466_port, QN => 
                           n_2071);
   IF_Regsxreg_file_regx18xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468324, Q => IF_Regsxreg_file_434_port, QN => 
                           n_2072);
   IF_Regsxreg_file_regx19xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468319, Q => IF_Regsxreg_file_402_port, QN => 
                           n_2073);
   IF_Regsxreg_file_regx20xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468314, Q => IF_Regsxreg_file_370_port, QN => 
                           n_2074);
   IF_Regsxreg_file_regx21xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468309, Q => IF_Regsxreg_file_338_port, QN => 
                           n_2075);
   IF_Regsxreg_file_regx22xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468304, Q => IF_Regsxreg_file_306_port, QN => 
                           n_2076);
   IF_Regsxreg_file_regx23xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468299, Q => IF_Regsxreg_file_274_port, QN => 
                           n_2077);
   IF_Regsxreg_file_regx24xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468294, Q => IF_Regsxreg_file_242_port, QN => 
                           n_2078);
   IF_Regsxreg_file_regx25xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468289, Q => IF_Regsxreg_file_210_port, QN => 
                           n_2079);
   IF_Regsxreg_file_regx26xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468284, Q => IF_Regsxreg_file_178_port, QN => 
                           n_2080);
   IF_Regsxreg_file_regx27xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468279, Q => IF_Regsxreg_file_146_port, QN => 
                           n_2081);
   IF_Regsxreg_file_regx28xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468274, Q => IF_Regsxreg_file_114_port, QN => 
                           n_2082);
   IF_Regsxreg_file_regx29xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468269, Q => IF_Regsxreg_file_82_port, QN => 
                           n_2083);
   IF_Regsxreg_file_regx30xx18x : DFF_X1 port map( D => IF_RegsxN678, CK => 
                           net2468264, Q => IF_Regsxreg_file_50_port, QN => 
                           n_2084);
   IF_RegsxRegsToCtl_port_contents2_regx18x : DFF_X1 port map( D => 
                           IF_RegsxN645, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_18_port, QN => n_2085);
   IF_CPathxRegsToCtl_data_signal_contents2_regx18x : DFF_X1 port map( D => 
                           IF_CPathxN2142, CK => net2468199, Q => n_2086, QN =>
                           n6306);
   IF_CPathxCtlToMem_port_dataIn_regx18x : DFF_X1 port map( D => n6458, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(18), QN => 
                           n_2087);
   IF_CPathxCtlToALU_port_reg2_contents_regx18x : DFF_X1 port map( D => n6603, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_18_port, QN => n_2088);
   IF_RegsxRegsToCtl_port_contents1_regx18x : DFF_X1 port map( D => 
                           IF_RegsxN613, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_18_port, QN => n_2089);
   IF_CPathxRegsToCtl_data_signal_contents1_regx18x : DFF_X1 port map( D => 
                           n6392, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_18_port, QN
                           => n6368);
   IF_CPathxCtlToALU_port_reg1_contents_regx18x : DFF_X1 port map( D => n6602, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_18_port, QN => n_2090);
   IF_ALUxALUtoCtl_port_regx4x : DFF_X1 port map( D => IF_ALUxN942, CK => 
                           net2468144, Q => ALUtoCtl_port_4_port, QN => n_2091)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx4x : DFF_X1 port map( D => IF_CPathxN1864,
                           CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_4_port, QN => n_2092);
   IF_CPathxCtlToMem_port_addrIn_regx4x : DFF_X1 port map( D => n6457, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(4), QN => 
                           n_2093);
   IF_CPathxCtlToRegs_port_dst_data_regx4x : DFF_X1 port map( D => n6558, CK =>
                           net2468214, Q => CtlToRegs_port_dst_data_4_port, QN 
                           => n_2094);
   IF_Regsxreg_file_regx31xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468259, Q => IF_Regsxreg_file_4_port, QN => 
                           n_2095);
   IF_Regsxreg_file_regx1xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468409, Q => IF_Regsxreg_file_964_port, QN => 
                           n_2096);
   IF_Regsxreg_file_regx2xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468404, Q => IF_Regsxreg_file_932_port, QN => 
                           n_2097);
   IF_Regsxreg_file_regx3xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468399, Q => IF_Regsxreg_file_900_port, QN => 
                           n_2098);
   IF_Regsxreg_file_regx4xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468394, Q => IF_Regsxreg_file_868_port, QN => 
                           n_2099);
   IF_Regsxreg_file_regx5xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468389, Q => IF_Regsxreg_file_836_port, QN => 
                           n_2100);
   IF_Regsxreg_file_regx6xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468384, Q => IF_Regsxreg_file_804_port, QN => 
                           n_2101);
   IF_Regsxreg_file_regx7xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468379, Q => IF_Regsxreg_file_772_port, QN => 
                           n_2102);
   IF_Regsxreg_file_regx8xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468374, Q => IF_Regsxreg_file_740_port, QN => 
                           n_2103);
   IF_Regsxreg_file_regx9xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468369, Q => IF_Regsxreg_file_708_port, QN => 
                           n_2104);
   IF_Regsxreg_file_regx10xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468364, Q => IF_Regsxreg_file_676_port, QN => 
                           n_2105);
   IF_Regsxreg_file_regx11xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468359, Q => IF_Regsxreg_file_644_port, QN => 
                           n_2106);
   IF_Regsxreg_file_regx12xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468354, Q => IF_Regsxreg_file_612_port, QN => 
                           n_2107);
   IF_Regsxreg_file_regx13xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468349, Q => IF_Regsxreg_file_580_port, QN => 
                           n_2108);
   IF_Regsxreg_file_regx14xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468344, Q => IF_Regsxreg_file_548_port, QN => 
                           n_2109);
   IF_Regsxreg_file_regx15xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468339, Q => IF_Regsxreg_file_516_port, QN => 
                           n_2110);
   IF_Regsxreg_file_regx16xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468334, Q => IF_Regsxreg_file_484_port, QN => 
                           n_2111);
   IF_Regsxreg_file_regx17xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468329, Q => IF_Regsxreg_file_452_port, QN => 
                           n_2112);
   IF_Regsxreg_file_regx18xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468324, Q => IF_Regsxreg_file_420_port, QN => 
                           n_2113);
   IF_Regsxreg_file_regx19xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468319, Q => IF_Regsxreg_file_388_port, QN => 
                           n_2114);
   IF_Regsxreg_file_regx20xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468314, Q => IF_Regsxreg_file_356_port, QN => 
                           n_2115);
   IF_Regsxreg_file_regx21xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468309, Q => IF_Regsxreg_file_324_port, QN => 
                           n_2116);
   IF_Regsxreg_file_regx22xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468304, Q => IF_Regsxreg_file_292_port, QN => 
                           n_2117);
   IF_Regsxreg_file_regx23xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468299, Q => IF_Regsxreg_file_260_port, QN => 
                           n_2118);
   IF_Regsxreg_file_regx24xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468294, Q => IF_Regsxreg_file_228_port, QN => 
                           n_2119);
   IF_Regsxreg_file_regx25xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468289, Q => IF_Regsxreg_file_196_port, QN => 
                           n_2120);
   IF_Regsxreg_file_regx26xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468284, Q => IF_Regsxreg_file_164_port, QN => 
                           n_2121);
   IF_Regsxreg_file_regx27xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468279, Q => IF_Regsxreg_file_132_port, QN => 
                           n_2122);
   IF_Regsxreg_file_regx28xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468274, Q => IF_Regsxreg_file_100_port, QN => 
                           n_2123);
   IF_Regsxreg_file_regx29xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468269, Q => IF_Regsxreg_file_68_port, QN => 
                           n_2124);
   IF_Regsxreg_file_regx30xx4x : DFF_X1 port map( D => IF_RegsxN664, CK => 
                           net2468264, Q => IF_Regsxreg_file_36_port, QN => 
                           n_2125);
   IF_RegsxRegsToCtl_port_contents2_regx4x : DFF_X1 port map( D => IF_RegsxN631
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents2_4_port, QN => n_2126);
   IF_CPathxRegsToCtl_data_signal_contents2_regx4x : DFF_X1 port map( D => 
                           IF_CPathxN2128, CK => net2468199, Q => n_2127, QN =>
                           n6307);
   IF_CPathxCtlToMem_port_dataIn_regx4x : DFF_X1 port map( D => n6456, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(4), QN => 
                           n_2128);
   IF_CPathxCtlToALU_port_reg2_contents_regx4x : DFF_X1 port map( D => n6601, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_4_port, QN => n_2129);
   IF_RegsxRegsToCtl_port_contents1_regx4x : DFF_X1 port map( D => IF_RegsxN599
                           , CK => net2468414, Q => n_2130, QN => n6374);
   IF_CPathxRegsToCtl_data_signal_contents1_regx4x : DFF_X1 port map( D => 
                           IF_CPathxN2096, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_4_port, QN 
                           => n6341);
   IF_CPathxCtlToALU_port_reg1_contents_regx4x : DFF_X1 port map( D => n6600, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_4_port, QN => n_2131);
   IF_ALUxALUtoCtl_port_regx14x : DFF_X1 port map( D => IF_ALUxN952, CK => 
                           net2468144, Q => ALUtoCtl_port_14_port, QN => n_2132
                           );
   IF_CPathxALUtoCtl_data_signal_regx14x : DFF_X1 port map( D => IF_CPathxN1874
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_14_port, QN => n_2133)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx14x : DFF_X1 port map( D => n6455, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(14), QN => 
                           n_2134);
   IF_CPathxCtlToRegs_port_dst_data_regx14x : DFF_X1 port map( D => n6557, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_14_port,
                           QN => n_2135);
   IF_Regsxreg_file_regx31xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468259, Q => IF_Regsxreg_file_14_port, QN => 
                           n_2136);
   IF_Regsxreg_file_regx1xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468409, Q => IF_Regsxreg_file_974_port, QN => 
                           n_2137);
   IF_Regsxreg_file_regx2xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468404, Q => IF_Regsxreg_file_942_port, QN => 
                           n_2138);
   IF_Regsxreg_file_regx3xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468399, Q => IF_Regsxreg_file_910_port, QN => 
                           n_2139);
   IF_Regsxreg_file_regx4xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468394, Q => IF_Regsxreg_file_878_port, QN => 
                           n_2140);
   IF_Regsxreg_file_regx5xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468389, Q => IF_Regsxreg_file_846_port, QN => 
                           n_2141);
   IF_Regsxreg_file_regx6xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468384, Q => IF_Regsxreg_file_814_port, QN => 
                           n_2142);
   IF_Regsxreg_file_regx7xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468379, Q => IF_Regsxreg_file_782_port, QN => 
                           n_2143);
   IF_Regsxreg_file_regx8xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468374, Q => IF_Regsxreg_file_750_port, QN => 
                           n_2144);
   IF_Regsxreg_file_regx9xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468369, Q => IF_Regsxreg_file_718_port, QN => 
                           n_2145);
   IF_Regsxreg_file_regx10xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468364, Q => IF_Regsxreg_file_686_port, QN => 
                           n_2146);
   IF_Regsxreg_file_regx11xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468359, Q => IF_Regsxreg_file_654_port, QN => 
                           n_2147);
   IF_Regsxreg_file_regx12xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468354, Q => IF_Regsxreg_file_622_port, QN => 
                           n_2148);
   IF_Regsxreg_file_regx13xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468349, Q => IF_Regsxreg_file_590_port, QN => 
                           n_2149);
   IF_Regsxreg_file_regx14xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468344, Q => IF_Regsxreg_file_558_port, QN => 
                           n_2150);
   IF_Regsxreg_file_regx15xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468339, Q => IF_Regsxreg_file_526_port, QN => 
                           n_2151);
   IF_Regsxreg_file_regx16xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468334, Q => IF_Regsxreg_file_494_port, QN => 
                           n_2152);
   IF_Regsxreg_file_regx17xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468329, Q => IF_Regsxreg_file_462_port, QN => 
                           n_2153);
   IF_Regsxreg_file_regx18xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468324, Q => IF_Regsxreg_file_430_port, QN => 
                           n_2154);
   IF_Regsxreg_file_regx19xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468319, Q => IF_Regsxreg_file_398_port, QN => 
                           n_2155);
   IF_Regsxreg_file_regx20xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468314, Q => IF_Regsxreg_file_366_port, QN => 
                           n_2156);
   IF_Regsxreg_file_regx21xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468309, Q => IF_Regsxreg_file_334_port, QN => 
                           n_2157);
   IF_Regsxreg_file_regx22xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468304, Q => IF_Regsxreg_file_302_port, QN => 
                           n_2158);
   IF_Regsxreg_file_regx23xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468299, Q => IF_Regsxreg_file_270_port, QN => 
                           n_2159);
   IF_Regsxreg_file_regx24xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468294, Q => IF_Regsxreg_file_238_port, QN => 
                           n_2160);
   IF_Regsxreg_file_regx25xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468289, Q => IF_Regsxreg_file_206_port, QN => 
                           n_2161);
   IF_Regsxreg_file_regx26xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468284, Q => IF_Regsxreg_file_174_port, QN => 
                           n_2162);
   IF_Regsxreg_file_regx27xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468279, Q => IF_Regsxreg_file_142_port, QN => 
                           n_2163);
   IF_Regsxreg_file_regx28xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468274, Q => IF_Regsxreg_file_110_port, QN => 
                           n_2164);
   IF_Regsxreg_file_regx29xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468269, Q => IF_Regsxreg_file_78_port, QN => 
                           n_2165);
   IF_Regsxreg_file_regx30xx14x : DFF_X1 port map( D => IF_RegsxN674, CK => 
                           net2468264, Q => IF_Regsxreg_file_46_port, QN => 
                           n_2166);
   IF_RegsxRegsToCtl_port_contents2_regx14x : DFF_X1 port map( D => 
                           IF_RegsxN641, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_14_port, QN => n_2167);
   IF_CPathxRegsToCtl_data_signal_contents2_regx14x : DFF_X1 port map( D => 
                           IF_CPathxN2138, CK => net2468199, Q => n_2168, QN =>
                           n6308);
   IF_CPathxCtlToMem_port_dataIn_regx14x : DFF_X1 port map( D => n6454, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(14), QN => 
                           n_2169);
   IF_CPathxCtlToALU_port_reg2_contents_regx14x : DFF_X1 port map( D => n6599, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_14_port, QN => n_2170);
   IF_RegsxRegsToCtl_port_contents1_regx14x : DFF_X1 port map( D => 
                           IF_RegsxN609, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_14_port, QN => n_2171);
   IF_CPathxRegsToCtl_data_signal_contents1_regx14x : DFF_X1 port map( D => 
                           n6388, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_14_port, QN
                           => n6355);
   IF_CPathxCtlToALU_port_reg1_contents_regx14x : DFF_X1 port map( D => n6598, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_14_port, QN => n_2172);
   IF_ALUxALUtoCtl_port_regx2x : DFF_X1 port map( D => IF_ALUxN940, CK => 
                           net2468144, Q => ALUtoCtl_port_2_port, QN => n_2173)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx2x : DFF_X1 port map( D => IF_CPathxN1862,
                           CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_2_port, QN => n_2174);
   IF_CPathxCtlToMem_port_addrIn_regx2x : DFF_X1 port map( D => n6453, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(2), QN => 
                           n_2175);
   IF_CPathxCtlToRegs_port_dst_data_regx2x : DFF_X1 port map( D => n6556, CK =>
                           net2468214, Q => CtlToRegs_port_dst_data_2_port, QN 
                           => n_2176);
   IF_Regsxreg_file_regx31xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468259, Q => IF_Regsxreg_file_2_port, QN => 
                           n_2177);
   IF_Regsxreg_file_regx1xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468409, Q => IF_Regsxreg_file_962_port, QN => 
                           n_2178);
   IF_Regsxreg_file_regx2xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468404, Q => IF_Regsxreg_file_930_port, QN => 
                           n_2179);
   IF_Regsxreg_file_regx3xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468399, Q => IF_Regsxreg_file_898_port, QN => 
                           n_2180);
   IF_Regsxreg_file_regx4xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468394, Q => IF_Regsxreg_file_866_port, QN => 
                           n_2181);
   IF_Regsxreg_file_regx5xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468389, Q => IF_Regsxreg_file_834_port, QN => 
                           n_2182);
   IF_Regsxreg_file_regx6xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468384, Q => IF_Regsxreg_file_802_port, QN => 
                           n_2183);
   IF_Regsxreg_file_regx7xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468379, Q => IF_Regsxreg_file_770_port, QN => 
                           n_2184);
   IF_Regsxreg_file_regx8xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468374, Q => IF_Regsxreg_file_738_port, QN => 
                           n_2185);
   IF_Regsxreg_file_regx9xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468369, Q => IF_Regsxreg_file_706_port, QN => 
                           n_2186);
   IF_Regsxreg_file_regx10xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468364, Q => IF_Regsxreg_file_674_port, QN => 
                           n_2187);
   IF_Regsxreg_file_regx11xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468359, Q => IF_Regsxreg_file_642_port, QN => 
                           n_2188);
   IF_Regsxreg_file_regx12xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468354, Q => IF_Regsxreg_file_610_port, QN => 
                           n_2189);
   IF_Regsxreg_file_regx13xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468349, Q => IF_Regsxreg_file_578_port, QN => 
                           n_2190);
   IF_Regsxreg_file_regx14xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468344, Q => IF_Regsxreg_file_546_port, QN => 
                           n_2191);
   IF_Regsxreg_file_regx15xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468339, Q => IF_Regsxreg_file_514_port, QN => 
                           n_2192);
   IF_Regsxreg_file_regx16xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468334, Q => IF_Regsxreg_file_482_port, QN => 
                           n_2193);
   IF_Regsxreg_file_regx17xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468329, Q => IF_Regsxreg_file_450_port, QN => 
                           n_2194);
   IF_Regsxreg_file_regx18xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468324, Q => IF_Regsxreg_file_418_port, QN => 
                           n_2195);
   IF_Regsxreg_file_regx19xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468319, Q => IF_Regsxreg_file_386_port, QN => 
                           n_2196);
   IF_Regsxreg_file_regx20xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468314, Q => IF_Regsxreg_file_354_port, QN => 
                           n_2197);
   IF_Regsxreg_file_regx21xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468309, Q => IF_Regsxreg_file_322_port, QN => 
                           n_2198);
   IF_Regsxreg_file_regx22xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468304, Q => IF_Regsxreg_file_290_port, QN => 
                           n_2199);
   IF_Regsxreg_file_regx23xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468299, Q => IF_Regsxreg_file_258_port, QN => 
                           n_2200);
   IF_Regsxreg_file_regx24xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468294, Q => IF_Regsxreg_file_226_port, QN => 
                           n_2201);
   IF_Regsxreg_file_regx25xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468289, Q => IF_Regsxreg_file_194_port, QN => 
                           n_2202);
   IF_Regsxreg_file_regx26xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468284, Q => IF_Regsxreg_file_162_port, QN => 
                           n_2203);
   IF_Regsxreg_file_regx27xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468279, Q => IF_Regsxreg_file_130_port, QN => 
                           n_2204);
   IF_Regsxreg_file_regx28xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468274, Q => IF_Regsxreg_file_98_port, QN => 
                           n_2205);
   IF_Regsxreg_file_regx29xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468269, Q => IF_Regsxreg_file_66_port, QN => 
                           n_2206);
   IF_Regsxreg_file_regx30xx2x : DFF_X1 port map( D => IF_RegsxN662, CK => 
                           net2468264, Q => IF_Regsxreg_file_34_port, QN => 
                           n_2207);
   IF_RegsxRegsToCtl_port_contents2_regx2x : DFF_X1 port map( D => IF_RegsxN629
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents2_2_port, QN => n_2208);
   IF_CPathxRegsToCtl_data_signal_contents2_regx2x : DFF_X1 port map( D => 
                           IF_CPathxN2126, CK => net2468199, Q => n_2209, QN =>
                           n6309);
   IF_CPathxCtlToMem_port_dataIn_regx2x : DFF_X1 port map( D => n6452, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(2), QN => 
                           n_2210);
   IF_CPathxCtlToALU_port_reg2_contents_regx2x : DFF_X1 port map( D => n6597, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_2_port, QN => n_2211);
   IF_RegsxRegsToCtl_port_contents1_regx2x : DFF_X1 port map( D => IF_RegsxN597
                           , CK => net2468414, Q => n_2212, QN => n6375);
   IF_CPathxRegsToCtl_data_signal_contents1_regx2x : DFF_X1 port map( D => 
                           IF_CPathxN2094, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_2_port, QN 
                           => n6342);
   IF_CPathxCtlToALU_port_reg1_contents_regx2x : DFF_X1 port map( D => n6596, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_2_port, QN => n_2213);
   IF_ALUxALUtoCtl_port_regx3x : DFF_X1 port map( D => IF_ALUxN941, CK => 
                           net2468144, Q => ALUtoCtl_port_3_port, QN => n6277);
   IF_CPathxALUtoCtl_data_signal_regx3x : DFF_X1 port map( D => IF_CPathxN1863,
                           CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_3_port, QN => n_2214);
   IF_CPathxCtlToMem_port_addrIn_regx3x : DFF_X1 port map( D => n6451, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(3), QN => 
                           n_2215);
   IF_CPathxCtlToRegs_port_dst_data_regx3x : DFF_X1 port map( D => n6555, CK =>
                           net2468214, Q => CtlToRegs_port_dst_data_3_port, QN 
                           => n_2216);
   IF_Regsxreg_file_regx31xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468259, Q => IF_Regsxreg_file_3_port, QN => 
                           n_2217);
   IF_Regsxreg_file_regx1xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468409, Q => IF_Regsxreg_file_963_port, QN => 
                           n_2218);
   IF_Regsxreg_file_regx2xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468404, Q => IF_Regsxreg_file_931_port, QN => 
                           n_2219);
   IF_Regsxreg_file_regx3xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468399, Q => IF_Regsxreg_file_899_port, QN => 
                           n_2220);
   IF_Regsxreg_file_regx4xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468394, Q => IF_Regsxreg_file_867_port, QN => 
                           n_2221);
   IF_Regsxreg_file_regx5xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468389, Q => IF_Regsxreg_file_835_port, QN => 
                           n_2222);
   IF_Regsxreg_file_regx6xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468384, Q => IF_Regsxreg_file_803_port, QN => 
                           n_2223);
   IF_Regsxreg_file_regx7xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468379, Q => IF_Regsxreg_file_771_port, QN => 
                           n_2224);
   IF_Regsxreg_file_regx8xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468374, Q => IF_Regsxreg_file_739_port, QN => 
                           n_2225);
   IF_Regsxreg_file_regx9xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468369, Q => IF_Regsxreg_file_707_port, QN => 
                           n_2226);
   IF_Regsxreg_file_regx10xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468364, Q => IF_Regsxreg_file_675_port, QN => 
                           n_2227);
   IF_Regsxreg_file_regx11xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468359, Q => IF_Regsxreg_file_643_port, QN => 
                           n_2228);
   IF_Regsxreg_file_regx12xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468354, Q => IF_Regsxreg_file_611_port, QN => 
                           n_2229);
   IF_Regsxreg_file_regx13xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468349, Q => IF_Regsxreg_file_579_port, QN => 
                           n_2230);
   IF_Regsxreg_file_regx14xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468344, Q => IF_Regsxreg_file_547_port, QN => 
                           n_2231);
   IF_Regsxreg_file_regx15xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468339, Q => IF_Regsxreg_file_515_port, QN => 
                           n_2232);
   IF_Regsxreg_file_regx16xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468334, Q => IF_Regsxreg_file_483_port, QN => 
                           n_2233);
   IF_Regsxreg_file_regx17xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468329, Q => IF_Regsxreg_file_451_port, QN => 
                           n_2234);
   IF_Regsxreg_file_regx18xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468324, Q => IF_Regsxreg_file_419_port, QN => 
                           n_2235);
   IF_Regsxreg_file_regx19xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468319, Q => IF_Regsxreg_file_387_port, QN => 
                           n_2236);
   IF_Regsxreg_file_regx20xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468314, Q => IF_Regsxreg_file_355_port, QN => 
                           n_2237);
   IF_Regsxreg_file_regx21xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468309, Q => IF_Regsxreg_file_323_port, QN => 
                           n_2238);
   IF_Regsxreg_file_regx22xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468304, Q => IF_Regsxreg_file_291_port, QN => 
                           n_2239);
   IF_Regsxreg_file_regx23xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468299, Q => IF_Regsxreg_file_259_port, QN => 
                           n_2240);
   IF_Regsxreg_file_regx24xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468294, Q => IF_Regsxreg_file_227_port, QN => 
                           n_2241);
   IF_Regsxreg_file_regx25xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468289, Q => IF_Regsxreg_file_195_port, QN => 
                           n_2242);
   IF_Regsxreg_file_regx26xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468284, Q => IF_Regsxreg_file_163_port, QN => 
                           n_2243);
   IF_Regsxreg_file_regx27xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468279, Q => IF_Regsxreg_file_131_port, QN => 
                           n_2244);
   IF_Regsxreg_file_regx28xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468274, Q => IF_Regsxreg_file_99_port, QN => 
                           n_2245);
   IF_Regsxreg_file_regx29xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468269, Q => IF_Regsxreg_file_67_port, QN => 
                           n_2246);
   IF_Regsxreg_file_regx30xx3x : DFF_X1 port map( D => IF_RegsxN663, CK => 
                           net2468264, Q => IF_Regsxreg_file_35_port, QN => 
                           n_2247);
   IF_RegsxRegsToCtl_port_contents2_regx3x : DFF_X1 port map( D => IF_RegsxN630
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents2_3_port, QN => n_2248);
   IF_CPathxRegsToCtl_data_signal_contents2_regx3x : DFF_X1 port map( D => 
                           IF_CPathxN2127, CK => net2468199, Q => n_2249, QN =>
                           n6310);
   IF_CPathxCtlToMem_port_dataIn_regx3x : DFF_X1 port map( D => n6450, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(3), QN => 
                           n_2250);
   IF_CPathxCtlToALU_port_reg2_contents_regx3x : DFF_X1 port map( D => n6595, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_3_port, QN => n_2251);
   IF_RegsxRegsToCtl_port_contents1_regx3x : DFF_X1 port map( D => IF_RegsxN598
                           , CK => net2468414, Q => n_2252, QN => n6376);
   IF_CPathxRegsToCtl_data_signal_contents1_regx3x : DFF_X1 port map( D => 
                           IF_CPathxN2095, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_3_port, QN 
                           => n6343);
   IF_CPathxCtlToALU_port_reg1_contents_regx3x : DFF_X1 port map( D => n6594, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_3_port, QN => n_2253);
   IF_ALUxALUtoCtl_port_regx1x : DFF_X1 port map( D => IF_ALUxN939, CK => 
                           net2468144, Q => ALUtoCtl_port_1_port, QN => n_2254)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx1x : DFF_X1 port map( D => IF_CPathxN1861,
                           CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_1_port, QN => n_2255);
   IF_CPathxCtlToMem_port_addrIn_regx1x : DFF_X1 port map( D => n6449, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(1), QN => 
                           n_2256);
   IF_CPathxCtlToRegs_port_dst_data_regx1x : DFF_X1 port map( D => n6554, CK =>
                           net2468214, Q => CtlToRegs_port_dst_data_1_port, QN 
                           => n_2257);
   IF_Regsxreg_file_regx31xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468259, Q => IF_Regsxreg_file_1_port, QN => 
                           n_2258);
   IF_Regsxreg_file_regx1xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468409, Q => IF_Regsxreg_file_961_port, QN => 
                           n_2259);
   IF_Regsxreg_file_regx2xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468404, Q => IF_Regsxreg_file_929_port, QN => 
                           n_2260);
   IF_Regsxreg_file_regx3xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468399, Q => IF_Regsxreg_file_897_port, QN => 
                           n_2261);
   IF_Regsxreg_file_regx4xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468394, Q => IF_Regsxreg_file_865_port, QN => 
                           n_2262);
   IF_Regsxreg_file_regx5xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468389, Q => IF_Regsxreg_file_833_port, QN => 
                           n_2263);
   IF_Regsxreg_file_regx6xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468384, Q => IF_Regsxreg_file_801_port, QN => 
                           n_2264);
   IF_Regsxreg_file_regx7xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468379, Q => IF_Regsxreg_file_769_port, QN => 
                           n_2265);
   IF_Regsxreg_file_regx8xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468374, Q => IF_Regsxreg_file_737_port, QN => 
                           n_2266);
   IF_Regsxreg_file_regx9xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468369, Q => IF_Regsxreg_file_705_port, QN => 
                           n_2267);
   IF_Regsxreg_file_regx10xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468364, Q => IF_Regsxreg_file_673_port, QN => 
                           n_2268);
   IF_Regsxreg_file_regx11xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468359, Q => IF_Regsxreg_file_641_port, QN => 
                           n_2269);
   IF_Regsxreg_file_regx12xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468354, Q => IF_Regsxreg_file_609_port, QN => 
                           n_2270);
   IF_Regsxreg_file_regx13xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468349, Q => IF_Regsxreg_file_577_port, QN => 
                           n_2271);
   IF_Regsxreg_file_regx14xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468344, Q => IF_Regsxreg_file_545_port, QN => 
                           n_2272);
   IF_Regsxreg_file_regx15xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468339, Q => IF_Regsxreg_file_513_port, QN => 
                           n_2273);
   IF_Regsxreg_file_regx16xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468334, Q => IF_Regsxreg_file_481_port, QN => 
                           n_2274);
   IF_Regsxreg_file_regx17xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468329, Q => IF_Regsxreg_file_449_port, QN => 
                           n_2275);
   IF_Regsxreg_file_regx18xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468324, Q => IF_Regsxreg_file_417_port, QN => 
                           n_2276);
   IF_Regsxreg_file_regx19xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468319, Q => IF_Regsxreg_file_385_port, QN => 
                           n_2277);
   IF_Regsxreg_file_regx20xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468314, Q => IF_Regsxreg_file_353_port, QN => 
                           n_2278);
   IF_Regsxreg_file_regx21xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468309, Q => IF_Regsxreg_file_321_port, QN => 
                           n_2279);
   IF_Regsxreg_file_regx22xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468304, Q => IF_Regsxreg_file_289_port, QN => 
                           n_2280);
   IF_Regsxreg_file_regx23xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468299, Q => IF_Regsxreg_file_257_port, QN => 
                           n_2281);
   IF_Regsxreg_file_regx24xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468294, Q => IF_Regsxreg_file_225_port, QN => 
                           n_2282);
   IF_Regsxreg_file_regx25xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468289, Q => IF_Regsxreg_file_193_port, QN => 
                           n_2283);
   IF_Regsxreg_file_regx26xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468284, Q => IF_Regsxreg_file_161_port, QN => 
                           n_2284);
   IF_Regsxreg_file_regx27xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468279, Q => IF_Regsxreg_file_129_port, QN => 
                           n_2285);
   IF_Regsxreg_file_regx28xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468274, Q => IF_Regsxreg_file_97_port, QN => 
                           n_2286);
   IF_Regsxreg_file_regx29xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468269, Q => IF_Regsxreg_file_65_port, QN => 
                           n_2287);
   IF_Regsxreg_file_regx30xx1x : DFF_X1 port map( D => IF_RegsxN661, CK => 
                           net2468264, Q => IF_Regsxreg_file_33_port, QN => 
                           n_2288);
   IF_RegsxRegsToCtl_port_contents2_regx1x : DFF_X1 port map( D => IF_RegsxN628
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents2_1_port, QN => n_2289);
   IF_CPathxRegsToCtl_data_signal_contents2_regx1x : DFF_X1 port map( D => 
                           IF_CPathxN2125, CK => net2468199, Q => n_2290, QN =>
                           n6311);
   IF_CPathxCtlToMem_port_dataIn_regx1x : DFF_X1 port map( D => n6448, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(1), QN => 
                           n_2291);
   IF_CPathxCtlToALU_port_reg2_contents_regx1x : DFF_X1 port map( D => n6593, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_1_port, QN => n_2292);
   IF_RegsxRegsToCtl_port_contents1_regx1x : DFF_X1 port map( D => IF_RegsxN596
                           , CK => net2468414, Q => n_2293, QN => n6377);
   IF_CPathxRegsToCtl_data_signal_contents1_regx1x : DFF_X1 port map( D => 
                           IF_CPathxN2092, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_1_port, QN 
                           => n6344);
   IF_CPathxCtlToALU_port_reg1_contents_regx1x : DFF_X1 port map( D => n6592, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_1_port, QN => n_2294);
   IF_ALUxALUtoCtl_port_regx5x : DFF_X1 port map( D => IF_ALUxN943, CK => 
                           net2468144, Q => ALUtoCtl_port_5_port, QN => n6280);
   IF_CPathxALUtoCtl_data_signal_regx5x : DFF_X1 port map( D => IF_CPathxN1865,
                           CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_5_port, QN => n_2295);
   IF_CPathxCtlToMem_port_addrIn_regx5x : DFF_X1 port map( D => n6447, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(5), QN => 
                           n_2296);
   IF_CPathxCtlToRegs_port_dst_data_regx5x : DFF_X1 port map( D => n6553, CK =>
                           net2468214, Q => CtlToRegs_port_dst_data_5_port, QN 
                           => n_2297);
   IF_Regsxreg_file_regx31xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468259, Q => IF_Regsxreg_file_5_port, QN => 
                           n_2298);
   IF_Regsxreg_file_regx1xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468409, Q => IF_Regsxreg_file_965_port, QN => 
                           n_2299);
   IF_Regsxreg_file_regx2xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468404, Q => IF_Regsxreg_file_933_port, QN => 
                           n_2300);
   IF_Regsxreg_file_regx3xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468399, Q => IF_Regsxreg_file_901_port, QN => 
                           n_2301);
   IF_Regsxreg_file_regx4xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468394, Q => IF_Regsxreg_file_869_port, QN => 
                           n_2302);
   IF_Regsxreg_file_regx5xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468389, Q => IF_Regsxreg_file_837_port, QN => 
                           n_2303);
   IF_Regsxreg_file_regx6xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468384, Q => IF_Regsxreg_file_805_port, QN => 
                           n_2304);
   IF_Regsxreg_file_regx7xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468379, Q => IF_Regsxreg_file_773_port, QN => 
                           n_2305);
   IF_Regsxreg_file_regx8xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468374, Q => IF_Regsxreg_file_741_port, QN => 
                           n_2306);
   IF_Regsxreg_file_regx9xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468369, Q => IF_Regsxreg_file_709_port, QN => 
                           n_2307);
   IF_Regsxreg_file_regx10xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468364, Q => IF_Regsxreg_file_677_port, QN => 
                           n_2308);
   IF_Regsxreg_file_regx11xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468359, Q => IF_Regsxreg_file_645_port, QN => 
                           n_2309);
   IF_Regsxreg_file_regx12xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468354, Q => IF_Regsxreg_file_613_port, QN => 
                           n_2310);
   IF_Regsxreg_file_regx13xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468349, Q => IF_Regsxreg_file_581_port, QN => 
                           n_2311);
   IF_Regsxreg_file_regx14xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468344, Q => IF_Regsxreg_file_549_port, QN => 
                           n_2312);
   IF_Regsxreg_file_regx15xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468339, Q => IF_Regsxreg_file_517_port, QN => 
                           n_2313);
   IF_Regsxreg_file_regx16xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468334, Q => IF_Regsxreg_file_485_port, QN => 
                           n_2314);
   IF_Regsxreg_file_regx17xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468329, Q => IF_Regsxreg_file_453_port, QN => 
                           n_2315);
   IF_Regsxreg_file_regx18xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468324, Q => IF_Regsxreg_file_421_port, QN => 
                           n_2316);
   IF_Regsxreg_file_regx19xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468319, Q => IF_Regsxreg_file_389_port, QN => 
                           n_2317);
   IF_Regsxreg_file_regx20xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468314, Q => IF_Regsxreg_file_357_port, QN => 
                           n_2318);
   IF_Regsxreg_file_regx21xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468309, Q => IF_Regsxreg_file_325_port, QN => 
                           n_2319);
   IF_Regsxreg_file_regx22xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468304, Q => IF_Regsxreg_file_293_port, QN => 
                           n_2320);
   IF_Regsxreg_file_regx23xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468299, Q => IF_Regsxreg_file_261_port, QN => 
                           n_2321);
   IF_Regsxreg_file_regx24xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468294, Q => IF_Regsxreg_file_229_port, QN => 
                           n_2322);
   IF_Regsxreg_file_regx25xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468289, Q => IF_Regsxreg_file_197_port, QN => 
                           n_2323);
   IF_Regsxreg_file_regx26xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468284, Q => IF_Regsxreg_file_165_port, QN => 
                           n_2324);
   IF_Regsxreg_file_regx27xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468279, Q => IF_Regsxreg_file_133_port, QN => 
                           n_2325);
   IF_Regsxreg_file_regx28xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468274, Q => IF_Regsxreg_file_101_port, QN => 
                           n_2326);
   IF_Regsxreg_file_regx29xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468269, Q => IF_Regsxreg_file_69_port, QN => 
                           n_2327);
   IF_Regsxreg_file_regx30xx5x : DFF_X1 port map( D => IF_RegsxN665, CK => 
                           net2468264, Q => IF_Regsxreg_file_37_port, QN => 
                           n_2328);
   IF_RegsxRegsToCtl_port_contents2_regx5x : DFF_X1 port map( D => IF_RegsxN632
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents2_5_port, QN => n_2329);
   IF_CPathxRegsToCtl_data_signal_contents2_regx5x : DFF_X1 port map( D => 
                           IF_CPathxN2129, CK => net2468199, Q => n_2330, QN =>
                           n6312);
   IF_CPathxCtlToMem_port_dataIn_regx5x : DFF_X1 port map( D => n6446, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(5), QN => 
                           n_2331);
   IF_CPathxCtlToALU_port_reg2_contents_regx5x : DFF_X1 port map( D => n6591, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_5_port, QN => n_2332);
   IF_RegsxRegsToCtl_port_contents1_regx5x : DFF_X1 port map( D => IF_RegsxN600
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents1_5_port, QN => n_2333);
   IF_CPathxRegsToCtl_data_signal_contents1_regx5x : DFF_X1 port map( D => 
                           n6379, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_5_port, QN 
                           => n6360);
   IF_CPathxCtlToALU_port_reg1_contents_regx5x : DFF_X1 port map( D => n6590, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_5_port, QN => n_2334);
   IF_ALUxALUtoCtl_port_regx7x : DFF_X1 port map( D => IF_ALUxN945, CK => 
                           net2468144, Q => ALUtoCtl_port_7_port, QN => n_2335)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx7x : DFF_X1 port map( D => IF_CPathxN1867,
                           CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_7_port, QN => n_2336);
   IF_CPathxCtlToMem_port_addrIn_regx7x : DFF_X1 port map( D => n6445, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(7), QN => 
                           n_2337);
   IF_CPathxCtlToRegs_port_dst_data_regx7x : DFF_X1 port map( D => n6552, CK =>
                           net2468214, Q => CtlToRegs_port_dst_data_7_port, QN 
                           => n_2338);
   IF_Regsxreg_file_regx31xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468259, Q => IF_Regsxreg_file_7_port, QN => 
                           n_2339);
   IF_Regsxreg_file_regx1xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468409, Q => IF_Regsxreg_file_967_port, QN => 
                           n_2340);
   IF_Regsxreg_file_regx2xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468404, Q => IF_Regsxreg_file_935_port, QN => 
                           n_2341);
   IF_Regsxreg_file_regx3xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468399, Q => IF_Regsxreg_file_903_port, QN => 
                           n_2342);
   IF_Regsxreg_file_regx4xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468394, Q => IF_Regsxreg_file_871_port, QN => 
                           n_2343);
   IF_Regsxreg_file_regx5xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468389, Q => IF_Regsxreg_file_839_port, QN => 
                           n_2344);
   IF_Regsxreg_file_regx6xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468384, Q => IF_Regsxreg_file_807_port, QN => 
                           n_2345);
   IF_Regsxreg_file_regx7xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468379, Q => IF_Regsxreg_file_775_port, QN => 
                           n_2346);
   IF_Regsxreg_file_regx8xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468374, Q => IF_Regsxreg_file_743_port, QN => 
                           n_2347);
   IF_Regsxreg_file_regx9xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468369, Q => IF_Regsxreg_file_711_port, QN => 
                           n_2348);
   IF_Regsxreg_file_regx10xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468364, Q => IF_Regsxreg_file_679_port, QN => 
                           n_2349);
   IF_Regsxreg_file_regx11xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468359, Q => IF_Regsxreg_file_647_port, QN => 
                           n_2350);
   IF_Regsxreg_file_regx12xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468354, Q => IF_Regsxreg_file_615_port, QN => 
                           n_2351);
   IF_Regsxreg_file_regx13xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468349, Q => IF_Regsxreg_file_583_port, QN => 
                           n_2352);
   IF_Regsxreg_file_regx14xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468344, Q => IF_Regsxreg_file_551_port, QN => 
                           n_2353);
   IF_Regsxreg_file_regx15xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468339, Q => IF_Regsxreg_file_519_port, QN => 
                           n_2354);
   IF_Regsxreg_file_regx16xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468334, Q => IF_Regsxreg_file_487_port, QN => 
                           n_2355);
   IF_Regsxreg_file_regx17xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468329, Q => IF_Regsxreg_file_455_port, QN => 
                           n_2356);
   IF_Regsxreg_file_regx18xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468324, Q => IF_Regsxreg_file_423_port, QN => 
                           n_2357);
   IF_Regsxreg_file_regx19xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468319, Q => IF_Regsxreg_file_391_port, QN => 
                           n_2358);
   IF_Regsxreg_file_regx20xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468314, Q => IF_Regsxreg_file_359_port, QN => 
                           n_2359);
   IF_Regsxreg_file_regx21xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468309, Q => IF_Regsxreg_file_327_port, QN => 
                           n_2360);
   IF_Regsxreg_file_regx22xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468304, Q => IF_Regsxreg_file_295_port, QN => 
                           n_2361);
   IF_Regsxreg_file_regx23xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468299, Q => IF_Regsxreg_file_263_port, QN => 
                           n_2362);
   IF_Regsxreg_file_regx24xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468294, Q => IF_Regsxreg_file_231_port, QN => 
                           n_2363);
   IF_Regsxreg_file_regx25xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468289, Q => IF_Regsxreg_file_199_port, QN => 
                           n_2364);
   IF_Regsxreg_file_regx26xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468284, Q => IF_Regsxreg_file_167_port, QN => 
                           n_2365);
   IF_Regsxreg_file_regx27xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468279, Q => IF_Regsxreg_file_135_port, QN => 
                           n_2366);
   IF_Regsxreg_file_regx28xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468274, Q => IF_Regsxreg_file_103_port, QN => 
                           n_2367);
   IF_Regsxreg_file_regx29xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468269, Q => IF_Regsxreg_file_71_port, QN => 
                           n_2368);
   IF_Regsxreg_file_regx30xx7x : DFF_X1 port map( D => IF_RegsxN667, CK => 
                           net2468264, Q => IF_Regsxreg_file_39_port, QN => 
                           n_2369);
   IF_RegsxRegsToCtl_port_contents2_regx7x : DFF_X1 port map( D => IF_RegsxN634
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents2_7_port, QN => n_2370);
   IF_CPathxRegsToCtl_data_signal_contents2_regx7x : DFF_X1 port map( D => 
                           IF_CPathxN2131, CK => net2468199, Q => n_2371, QN =>
                           n6313);
   IF_CPathxCtlToMem_port_dataIn_regx7x : DFF_X1 port map( D => n6444, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(7), QN => 
                           n_2372);
   IF_CPathxCtlToALU_port_reg2_contents_regx7x : DFF_X1 port map( D => n6589, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_7_port, QN => n_2373);
   IF_RegsxRegsToCtl_port_contents1_regx7x : DFF_X1 port map( D => IF_RegsxN602
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents1_7_port, QN => n_2374);
   IF_CPathxRegsToCtl_data_signal_contents1_regx7x : DFF_X1 port map( D => 
                           n6381, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_7_port, QN 
                           => n6362);
   IF_CPathxCtlToALU_port_reg1_contents_regx7x : DFF_X1 port map( D => n6588, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_7_port, QN => n_2375);
   IF_ALUxALUtoCtl_port_regx25x : DFF_X1 port map( D => IF_ALUxN963, CK => 
                           net2468144, Q => ALUtoCtl_port_25_port, QN => n_2376
                           );
   IF_CPathxALUtoCtl_data_signal_regx25x : DFF_X1 port map( D => IF_CPathxN1885
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_25_port, QN => n_2377)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx25x : DFF_X1 port map( D => n6443, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(25), QN => 
                           n_2378);
   IF_CPathxCtlToRegs_port_dst_data_regx25x : DFF_X1 port map( D => n6551, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_25_port,
                           QN => n_2379);
   IF_Regsxreg_file_regx31xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468259, Q => IF_Regsxreg_file_25_port, QN => 
                           n_2380);
   IF_Regsxreg_file_regx1xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468409, Q => IF_Regsxreg_file_985_port, QN => 
                           n_2381);
   IF_Regsxreg_file_regx2xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468404, Q => IF_Regsxreg_file_953_port, QN => 
                           n_2382);
   IF_Regsxreg_file_regx3xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468399, Q => IF_Regsxreg_file_921_port, QN => 
                           n_2383);
   IF_Regsxreg_file_regx4xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468394, Q => IF_Regsxreg_file_889_port, QN => 
                           n_2384);
   IF_Regsxreg_file_regx5xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468389, Q => IF_Regsxreg_file_857_port, QN => 
                           n_2385);
   IF_Regsxreg_file_regx6xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468384, Q => IF_Regsxreg_file_825_port, QN => 
                           n_2386);
   IF_Regsxreg_file_regx7xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468379, Q => IF_Regsxreg_file_793_port, QN => 
                           n_2387);
   IF_Regsxreg_file_regx8xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468374, Q => IF_Regsxreg_file_761_port, QN => 
                           n_2388);
   IF_Regsxreg_file_regx9xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468369, Q => IF_Regsxreg_file_729_port, QN => 
                           n_2389);
   IF_Regsxreg_file_regx10xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468364, Q => IF_Regsxreg_file_697_port, QN => 
                           n_2390);
   IF_Regsxreg_file_regx11xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468359, Q => IF_Regsxreg_file_665_port, QN => 
                           n_2391);
   IF_Regsxreg_file_regx12xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468354, Q => IF_Regsxreg_file_633_port, QN => 
                           n_2392);
   IF_Regsxreg_file_regx13xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468349, Q => IF_Regsxreg_file_601_port, QN => 
                           n_2393);
   IF_Regsxreg_file_regx14xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468344, Q => IF_Regsxreg_file_569_port, QN => 
                           n_2394);
   IF_Regsxreg_file_regx15xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468339, Q => IF_Regsxreg_file_537_port, QN => 
                           n_2395);
   IF_Regsxreg_file_regx16xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468334, Q => IF_Regsxreg_file_505_port, QN => 
                           n_2396);
   IF_Regsxreg_file_regx17xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468329, Q => IF_Regsxreg_file_473_port, QN => 
                           n_2397);
   IF_Regsxreg_file_regx18xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468324, Q => IF_Regsxreg_file_441_port, QN => 
                           n_2398);
   IF_Regsxreg_file_regx19xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468319, Q => IF_Regsxreg_file_409_port, QN => 
                           n_2399);
   IF_Regsxreg_file_regx20xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468314, Q => IF_Regsxreg_file_377_port, QN => 
                           n_2400);
   IF_Regsxreg_file_regx21xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468309, Q => IF_Regsxreg_file_345_port, QN => 
                           n_2401);
   IF_Regsxreg_file_regx22xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468304, Q => IF_Regsxreg_file_313_port, QN => 
                           n_2402);
   IF_Regsxreg_file_regx23xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468299, Q => IF_Regsxreg_file_281_port, QN => 
                           n_2403);
   IF_Regsxreg_file_regx24xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468294, Q => IF_Regsxreg_file_249_port, QN => 
                           n_2404);
   IF_Regsxreg_file_regx25xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468289, Q => IF_Regsxreg_file_217_port, QN => 
                           n_2405);
   IF_Regsxreg_file_regx26xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468284, Q => IF_Regsxreg_file_185_port, QN => 
                           n_2406);
   IF_Regsxreg_file_regx27xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468279, Q => IF_Regsxreg_file_153_port, QN => 
                           n_2407);
   IF_Regsxreg_file_regx28xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468274, Q => IF_Regsxreg_file_121_port, QN => 
                           n_2408);
   IF_Regsxreg_file_regx29xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468269, Q => IF_Regsxreg_file_89_port, QN => 
                           n_2409);
   IF_Regsxreg_file_regx30xx25x : DFF_X1 port map( D => IF_RegsxN685, CK => 
                           net2468264, Q => IF_Regsxreg_file_57_port, QN => 
                           n_2410);
   IF_RegsxRegsToCtl_port_contents2_regx25x : DFF_X1 port map( D => 
                           IF_RegsxN652, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_25_port, QN => n_2411);
   IF_CPathxRegsToCtl_data_signal_contents2_regx25x : DFF_X1 port map( D => 
                           IF_CPathxN2149, CK => net2468199, Q => n_2412, QN =>
                           n6314);
   IF_CPathxCtlToMem_port_dataIn_regx25x : DFF_X1 port map( D => n6442, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(25), QN => 
                           n_2413);
   IF_CPathxCtlToALU_port_reg2_contents_regx25x : DFF_X1 port map( D => n6587, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_25_port, QN => n_2414);
   IF_RegsxRegsToCtl_port_contents1_regx25x : DFF_X1 port map( D => 
                           IF_RegsxN620, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_25_port, QN => n_2415);
   IF_CPathxRegsToCtl_data_signal_contents1_regx25x : DFF_X1 port map( D => 
                           n6399, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_25_port, QN
                           => n6349);
   IF_CPathxCtlToALU_port_reg1_contents_regx25x : DFF_X1 port map( D => n6586, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_25_port, QN => n_2416);
   IF_ALUxALUtoCtl_port_regx9x : DFF_X1 port map( D => IF_ALUxN947, CK => 
                           net2468144, Q => ALUtoCtl_port_9_port, QN => n6281);
   IF_CPathxALUtoCtl_data_signal_regx9x : DFF_X1 port map( D => IF_CPathxN1869,
                           CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_9_port, QN => n_2417);
   IF_CPathxCtlToMem_port_addrIn_regx9x : DFF_X1 port map( D => n6441, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(9), QN => 
                           n_2418);
   IF_CPathxCtlToRegs_port_dst_data_regx9x : DFF_X1 port map( D => n6550, CK =>
                           net2468214, Q => CtlToRegs_port_dst_data_9_port, QN 
                           => n_2419);
   IF_Regsxreg_file_regx31xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468259, Q => IF_Regsxreg_file_9_port, QN => 
                           n_2420);
   IF_Regsxreg_file_regx1xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468409, Q => IF_Regsxreg_file_969_port, QN => 
                           n_2421);
   IF_Regsxreg_file_regx2xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468404, Q => IF_Regsxreg_file_937_port, QN => 
                           n_2422);
   IF_Regsxreg_file_regx3xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468399, Q => IF_Regsxreg_file_905_port, QN => 
                           n_2423);
   IF_Regsxreg_file_regx4xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468394, Q => IF_Regsxreg_file_873_port, QN => 
                           n_2424);
   IF_Regsxreg_file_regx5xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468389, Q => IF_Regsxreg_file_841_port, QN => 
                           n_2425);
   IF_Regsxreg_file_regx6xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468384, Q => IF_Regsxreg_file_809_port, QN => 
                           n_2426);
   IF_Regsxreg_file_regx7xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468379, Q => IF_Regsxreg_file_777_port, QN => 
                           n_2427);
   IF_Regsxreg_file_regx8xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468374, Q => IF_Regsxreg_file_745_port, QN => 
                           n_2428);
   IF_Regsxreg_file_regx9xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468369, Q => IF_Regsxreg_file_713_port, QN => 
                           n_2429);
   IF_Regsxreg_file_regx10xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468364, Q => IF_Regsxreg_file_681_port, QN => 
                           n_2430);
   IF_Regsxreg_file_regx11xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468359, Q => IF_Regsxreg_file_649_port, QN => 
                           n_2431);
   IF_Regsxreg_file_regx12xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468354, Q => IF_Regsxreg_file_617_port, QN => 
                           n_2432);
   IF_Regsxreg_file_regx13xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468349, Q => IF_Regsxreg_file_585_port, QN => 
                           n_2433);
   IF_Regsxreg_file_regx14xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468344, Q => IF_Regsxreg_file_553_port, QN => 
                           n_2434);
   IF_Regsxreg_file_regx15xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468339, Q => IF_Regsxreg_file_521_port, QN => 
                           n_2435);
   IF_Regsxreg_file_regx16xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468334, Q => IF_Regsxreg_file_489_port, QN => 
                           n_2436);
   IF_Regsxreg_file_regx17xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468329, Q => IF_Regsxreg_file_457_port, QN => 
                           n_2437);
   IF_Regsxreg_file_regx18xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468324, Q => IF_Regsxreg_file_425_port, QN => 
                           n_2438);
   IF_Regsxreg_file_regx19xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468319, Q => IF_Regsxreg_file_393_port, QN => 
                           n_2439);
   IF_Regsxreg_file_regx20xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468314, Q => IF_Regsxreg_file_361_port, QN => 
                           n_2440);
   IF_Regsxreg_file_regx21xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468309, Q => IF_Regsxreg_file_329_port, QN => 
                           n_2441);
   IF_Regsxreg_file_regx22xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468304, Q => IF_Regsxreg_file_297_port, QN => 
                           n_2442);
   IF_Regsxreg_file_regx23xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468299, Q => IF_Regsxreg_file_265_port, QN => 
                           n_2443);
   IF_Regsxreg_file_regx24xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468294, Q => IF_Regsxreg_file_233_port, QN => 
                           n_2444);
   IF_Regsxreg_file_regx25xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468289, Q => IF_Regsxreg_file_201_port, QN => 
                           n_2445);
   IF_Regsxreg_file_regx26xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468284, Q => IF_Regsxreg_file_169_port, QN => 
                           n_2446);
   IF_Regsxreg_file_regx27xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468279, Q => IF_Regsxreg_file_137_port, QN => 
                           n_2447);
   IF_Regsxreg_file_regx28xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468274, Q => IF_Regsxreg_file_105_port, QN => 
                           n_2448);
   IF_Regsxreg_file_regx29xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468269, Q => IF_Regsxreg_file_73_port, QN => 
                           n_2449);
   IF_Regsxreg_file_regx30xx9x : DFF_X1 port map( D => IF_RegsxN669, CK => 
                           net2468264, Q => IF_Regsxreg_file_41_port, QN => 
                           n_2450);
   IF_RegsxRegsToCtl_port_contents2_regx9x : DFF_X1 port map( D => IF_RegsxN636
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents2_9_port, QN => n_2451);
   IF_CPathxRegsToCtl_data_signal_contents2_regx9x : DFF_X1 port map( D => 
                           IF_CPathxN2133, CK => net2468199, Q => n_2452, QN =>
                           n6315);
   IF_CPathxCtlToMem_port_dataIn_regx9x : DFF_X1 port map( D => n6440, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(9), QN => 
                           n_2453);
   IF_CPathxCtlToALU_port_reg2_contents_regx9x : DFF_X1 port map( D => n6585, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_9_port, QN => n_2454);
   IF_RegsxRegsToCtl_port_contents1_regx9x : DFF_X1 port map( D => IF_RegsxN604
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents1_9_port, QN => n_2455);
   IF_CPathxRegsToCtl_data_signal_contents1_regx9x : DFF_X1 port map( D => 
                           n6383, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_9_port, QN 
                           => n6359);
   IF_CPathxCtlToALU_port_reg1_contents_regx9x : DFF_X1 port map( D => n6584, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_9_port, QN => n_2456);
   IF_ALUxALUtoCtl_port_regx6x : DFF_X1 port map( D => IF_ALUxN944, CK => 
                           net2468144, Q => ALUtoCtl_port_6_port, QN => n_2457)
                           ;
   IF_CPathxALUtoCtl_data_signal_regx6x : DFF_X1 port map( D => IF_CPathxN1866,
                           CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_6_port, QN => n_2458);
   IF_CPathxCtlToMem_port_addrIn_regx6x : DFF_X1 port map( D => n6439, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(6), QN => 
                           n_2459);
   IF_CPathxCtlToRegs_port_dst_data_regx6x : DFF_X1 port map( D => n6549, CK =>
                           net2468214, Q => CtlToRegs_port_dst_data_6_port, QN 
                           => n_2460);
   IF_Regsxreg_file_regx31xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468259, Q => IF_Regsxreg_file_6_port, QN => 
                           n_2461);
   IF_Regsxreg_file_regx1xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468409, Q => IF_Regsxreg_file_966_port, QN => 
                           n_2462);
   IF_Regsxreg_file_regx2xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468404, Q => IF_Regsxreg_file_934_port, QN => 
                           n_2463);
   IF_Regsxreg_file_regx3xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468399, Q => IF_Regsxreg_file_902_port, QN => 
                           n_2464);
   IF_Regsxreg_file_regx4xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468394, Q => IF_Regsxreg_file_870_port, QN => 
                           n_2465);
   IF_Regsxreg_file_regx5xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468389, Q => IF_Regsxreg_file_838_port, QN => 
                           n_2466);
   IF_Regsxreg_file_regx6xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468384, Q => IF_Regsxreg_file_806_port, QN => 
                           n_2467);
   IF_Regsxreg_file_regx7xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468379, Q => IF_Regsxreg_file_774_port, QN => 
                           n_2468);
   IF_Regsxreg_file_regx8xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468374, Q => IF_Regsxreg_file_742_port, QN => 
                           n_2469);
   IF_Regsxreg_file_regx9xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468369, Q => IF_Regsxreg_file_710_port, QN => 
                           n_2470);
   IF_Regsxreg_file_regx10xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468364, Q => IF_Regsxreg_file_678_port, QN => 
                           n_2471);
   IF_Regsxreg_file_regx11xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468359, Q => IF_Regsxreg_file_646_port, QN => 
                           n_2472);
   IF_Regsxreg_file_regx12xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468354, Q => IF_Regsxreg_file_614_port, QN => 
                           n_2473);
   IF_Regsxreg_file_regx13xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468349, Q => IF_Regsxreg_file_582_port, QN => 
                           n_2474);
   IF_Regsxreg_file_regx14xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468344, Q => IF_Regsxreg_file_550_port, QN => 
                           n_2475);
   IF_Regsxreg_file_regx15xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468339, Q => IF_Regsxreg_file_518_port, QN => 
                           n_2476);
   IF_Regsxreg_file_regx16xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468334, Q => IF_Regsxreg_file_486_port, QN => 
                           n_2477);
   IF_Regsxreg_file_regx17xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468329, Q => IF_Regsxreg_file_454_port, QN => 
                           n_2478);
   IF_Regsxreg_file_regx18xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468324, Q => IF_Regsxreg_file_422_port, QN => 
                           n_2479);
   IF_Regsxreg_file_regx19xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468319, Q => IF_Regsxreg_file_390_port, QN => 
                           n_2480);
   IF_Regsxreg_file_regx20xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468314, Q => IF_Regsxreg_file_358_port, QN => 
                           n_2481);
   IF_Regsxreg_file_regx21xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468309, Q => IF_Regsxreg_file_326_port, QN => 
                           n_2482);
   IF_Regsxreg_file_regx22xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468304, Q => IF_Regsxreg_file_294_port, QN => 
                           n_2483);
   IF_Regsxreg_file_regx23xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468299, Q => IF_Regsxreg_file_262_port, QN => 
                           n_2484);
   IF_Regsxreg_file_regx24xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468294, Q => IF_Regsxreg_file_230_port, QN => 
                           n_2485);
   IF_Regsxreg_file_regx25xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468289, Q => IF_Regsxreg_file_198_port, QN => 
                           n_2486);
   IF_Regsxreg_file_regx26xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468284, Q => IF_Regsxreg_file_166_port, QN => 
                           n_2487);
   IF_Regsxreg_file_regx27xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468279, Q => IF_Regsxreg_file_134_port, QN => 
                           n_2488);
   IF_Regsxreg_file_regx28xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468274, Q => IF_Regsxreg_file_102_port, QN => 
                           n_2489);
   IF_Regsxreg_file_regx29xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468269, Q => IF_Regsxreg_file_70_port, QN => 
                           n_2490);
   IF_Regsxreg_file_regx30xx6x : DFF_X1 port map( D => IF_RegsxN666, CK => 
                           net2468264, Q => IF_Regsxreg_file_38_port, QN => 
                           n_2491);
   IF_RegsxRegsToCtl_port_contents2_regx6x : DFF_X1 port map( D => IF_RegsxN633
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents2_6_port, QN => n_2492);
   IF_CPathxRegsToCtl_data_signal_contents2_regx6x : DFF_X1 port map( D => 
                           IF_CPathxN2130, CK => net2468199, Q => n_2493, QN =>
                           n6316);
   IF_CPathxCtlToMem_port_dataIn_regx6x : DFF_X1 port map( D => n6438, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(6), QN => 
                           n_2494);
   IF_CPathxCtlToALU_port_reg2_contents_regx6x : DFF_X1 port map( D => n6583, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_6_port, QN => n_2495);
   IF_RegsxRegsToCtl_port_contents1_regx6x : DFF_X1 port map( D => IF_RegsxN601
                           , CK => net2468414, Q => 
                           RegsToCtl_port_contents1_6_port, QN => n_2496);
   IF_CPathxRegsToCtl_data_signal_contents1_regx6x : DFF_X1 port map( D => 
                           n6380, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_6_port, QN 
                           => n6361);
   IF_CPathxCtlToALU_port_reg1_contents_regx6x : DFF_X1 port map( D => n6582, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_6_port, QN => n_2497);
   IF_ALUxALUtoCtl_port_regx30x : DFF_X1 port map( D => IF_ALUxN968, CK => 
                           net2468144, Q => ALUtoCtl_port_30_port, QN => n_2498
                           );
   IF_CPathxALUtoCtl_data_signal_regx30x : DFF_X1 port map( D => IF_CPathxN1890
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_30_port, QN => n_2499)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx30x : DFF_X1 port map( D => n6437, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(30), QN => 
                           n_2500);
   IF_CPathxCtlToRegs_port_dst_data_regx30x : DFF_X1 port map( D => n6548, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_30_port,
                           QN => n_2501);
   IF_Regsxreg_file_regx31xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468259, Q => IF_Regsxreg_file_30_port, QN => 
                           n_2502);
   IF_Regsxreg_file_regx1xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468409, Q => IF_Regsxreg_file_990_port, QN => 
                           n_2503);
   IF_Regsxreg_file_regx2xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468404, Q => IF_Regsxreg_file_958_port, QN => 
                           n_2504);
   IF_Regsxreg_file_regx3xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468399, Q => IF_Regsxreg_file_926_port, QN => 
                           n_2505);
   IF_Regsxreg_file_regx4xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468394, Q => IF_Regsxreg_file_894_port, QN => 
                           n_2506);
   IF_Regsxreg_file_regx5xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468389, Q => IF_Regsxreg_file_862_port, QN => 
                           n_2507);
   IF_Regsxreg_file_regx6xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468384, Q => IF_Regsxreg_file_830_port, QN => 
                           n_2508);
   IF_Regsxreg_file_regx7xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468379, Q => IF_Regsxreg_file_798_port, QN => 
                           n_2509);
   IF_Regsxreg_file_regx8xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468374, Q => IF_Regsxreg_file_766_port, QN => 
                           n_2510);
   IF_Regsxreg_file_regx9xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468369, Q => IF_Regsxreg_file_734_port, QN => 
                           n_2511);
   IF_Regsxreg_file_regx10xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468364, Q => IF_Regsxreg_file_702_port, QN => 
                           n_2512);
   IF_Regsxreg_file_regx11xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468359, Q => IF_Regsxreg_file_670_port, QN => 
                           n_2513);
   IF_Regsxreg_file_regx12xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468354, Q => IF_Regsxreg_file_638_port, QN => 
                           n_2514);
   IF_Regsxreg_file_regx13xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468349, Q => IF_Regsxreg_file_606_port, QN => 
                           n_2515);
   IF_Regsxreg_file_regx14xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468344, Q => IF_Regsxreg_file_574_port, QN => 
                           n_2516);
   IF_Regsxreg_file_regx15xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468339, Q => IF_Regsxreg_file_542_port, QN => 
                           n_2517);
   IF_Regsxreg_file_regx16xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468334, Q => IF_Regsxreg_file_510_port, QN => 
                           n_2518);
   IF_Regsxreg_file_regx17xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468329, Q => IF_Regsxreg_file_478_port, QN => 
                           n_2519);
   IF_Regsxreg_file_regx18xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468324, Q => IF_Regsxreg_file_446_port, QN => 
                           n_2520);
   IF_Regsxreg_file_regx19xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468319, Q => IF_Regsxreg_file_414_port, QN => 
                           n_2521);
   IF_Regsxreg_file_regx20xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468314, Q => IF_Regsxreg_file_382_port, QN => 
                           n_2522);
   IF_Regsxreg_file_regx21xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468309, Q => IF_Regsxreg_file_350_port, QN => 
                           n_2523);
   IF_Regsxreg_file_regx22xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468304, Q => IF_Regsxreg_file_318_port, QN => 
                           n_2524);
   IF_Regsxreg_file_regx23xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468299, Q => IF_Regsxreg_file_286_port, QN => 
                           n_2525);
   IF_Regsxreg_file_regx24xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468294, Q => IF_Regsxreg_file_254_port, QN => 
                           n_2526);
   IF_Regsxreg_file_regx25xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468289, Q => IF_Regsxreg_file_222_port, QN => 
                           n_2527);
   IF_Regsxreg_file_regx26xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468284, Q => IF_Regsxreg_file_190_port, QN => 
                           n_2528);
   IF_Regsxreg_file_regx27xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468279, Q => IF_Regsxreg_file_158_port, QN => 
                           n_2529);
   IF_Regsxreg_file_regx28xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468274, Q => IF_Regsxreg_file_126_port, QN => 
                           n_2530);
   IF_Regsxreg_file_regx29xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468269, Q => IF_Regsxreg_file_94_port, QN => 
                           n_2531);
   IF_Regsxreg_file_regx30xx30x : DFF_X1 port map( D => IF_RegsxN690, CK => 
                           net2468264, Q => IF_Regsxreg_file_62_port, QN => 
                           n_2532);
   IF_RegsxRegsToCtl_port_contents2_regx30x : DFF_X1 port map( D => 
                           IF_RegsxN657, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_30_port, QN => n_2533);
   IF_CPathxRegsToCtl_data_signal_contents2_regx30x : DFF_X1 port map( D => 
                           IF_CPathxN2154, CK => net2468199, Q => n_2534, QN =>
                           n6317);
   IF_CPathxCtlToMem_port_dataIn_regx30x : DFF_X1 port map( D => n6436, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(30), QN => 
                           n_2535);
   IF_CPathxCtlToALU_port_reg2_contents_regx30x : DFF_X1 port map( D => n6581, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_30_port, QN => n_2536);
   IF_RegsxRegsToCtl_port_contents1_regx30x : DFF_X1 port map( D => 
                           IF_RegsxN625, CK => net2468414, Q => 
                           RegsToCtl_port_contents1_30_port, QN => n_2537);
   IF_CPathxRegsToCtl_data_signal_contents1_regx30x : DFF_X1 port map( D => 
                           n6404, CK => net2468199, Q => 
                           IF_CPathxRegsToCtl_data_signal_contents1_30_port, QN
                           => n6372);
   IF_CPathxCtlToALU_port_reg1_contents_regx30x : DFF_X1 port map( D => n6580, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg1_contents_30_port, QN => n_2538);
   IF_CPathxpc_next_signal_regx31x : DFF_X1 port map( D => IF_CPathxN2273, CK 
                           => net2468179, Q => IF_CPathxpc_next_signal_31_port,
                           QN => n_2539);
   IF_CPathxpc_reg_signal_regx31x : DFF_X1 port map( D => n6506, CK => 
                           net2468174, Q => IF_CPathxpc_reg_signal_31_port, QN 
                           => n_2540);
   IF_CPathxCtlToALU_port_pc_reg_regx31x : DFF_X1 port map( D => IF_CPathxN1967
                           , CK => net2468224, Q => 
                           CtlToALU_port_pc_reg_31_port, QN => n_2541);
   IF_CPathxALUtoCtl_data_signal_regx31x : DFF_X1 port map( D => IF_CPathxN1891
                           , CK => net2468179, Q => 
                           IF_CPathxALUtoCtl_data_signal_31_port, QN => n_2542)
                           ;
   IF_CPathxCtlToMem_port_addrIn_regx31x : DFF_X1 port map( D => n6435, CK => 
                           net2468164, Q => CtlToMem_port_addrIn(31), QN => 
                           n_2543);
   IF_CPathxCtlToRegs_port_dst_data_regx31x : DFF_X1 port map( D => n6547, CK 
                           => net2468214, Q => CtlToRegs_port_dst_data_31_port,
                           QN => n_2544);
   IF_Regsxreg_file_regx31xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468259, Q => IF_Regsxreg_file_31_port, QN => 
                           n_2545);
   IF_Regsxreg_file_regx1xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468409, Q => IF_Regsxreg_file_991_port, QN => 
                           n_2546);
   IF_Regsxreg_file_regx2xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468404, Q => IF_Regsxreg_file_959_port, QN => 
                           n_2547);
   IF_Regsxreg_file_regx3xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468399, Q => IF_Regsxreg_file_927_port, QN => 
                           n_2548);
   IF_Regsxreg_file_regx4xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468394, Q => IF_Regsxreg_file_895_port, QN => 
                           n_2549);
   IF_Regsxreg_file_regx5xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468389, Q => IF_Regsxreg_file_863_port, QN => 
                           n_2550);
   IF_Regsxreg_file_regx6xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468384, Q => IF_Regsxreg_file_831_port, QN => 
                           n_2551);
   IF_Regsxreg_file_regx7xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468379, Q => IF_Regsxreg_file_799_port, QN => 
                           n_2552);
   IF_Regsxreg_file_regx8xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468374, Q => IF_Regsxreg_file_767_port, QN => 
                           n_2553);
   IF_Regsxreg_file_regx9xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468369, Q => IF_Regsxreg_file_735_port, QN => 
                           n_2554);
   IF_Regsxreg_file_regx10xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468364, Q => IF_Regsxreg_file_703_port, QN => 
                           n_2555);
   IF_Regsxreg_file_regx11xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468359, Q => IF_Regsxreg_file_671_port, QN => 
                           n_2556);
   IF_Regsxreg_file_regx12xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468354, Q => IF_Regsxreg_file_639_port, QN => 
                           n_2557);
   IF_Regsxreg_file_regx13xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468349, Q => IF_Regsxreg_file_607_port, QN => 
                           n_2558);
   IF_Regsxreg_file_regx14xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468344, Q => IF_Regsxreg_file_575_port, QN => 
                           n_2559);
   IF_Regsxreg_file_regx15xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468339, Q => IF_Regsxreg_file_543_port, QN => 
                           n_2560);
   IF_Regsxreg_file_regx16xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468334, Q => IF_Regsxreg_file_511_port, QN => 
                           n_2561);
   IF_Regsxreg_file_regx17xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468329, Q => IF_Regsxreg_file_479_port, QN => 
                           n_2562);
   IF_Regsxreg_file_regx18xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468324, Q => IF_Regsxreg_file_447_port, QN => 
                           n_2563);
   IF_Regsxreg_file_regx19xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468319, Q => IF_Regsxreg_file_415_port, QN => 
                           n_2564);
   IF_Regsxreg_file_regx20xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468314, Q => IF_Regsxreg_file_383_port, QN => 
                           n_2565);
   IF_Regsxreg_file_regx21xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468309, Q => IF_Regsxreg_file_351_port, QN => 
                           n_2566);
   IF_Regsxreg_file_regx22xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468304, Q => IF_Regsxreg_file_319_port, QN => 
                           n_2567);
   IF_Regsxreg_file_regx23xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468299, Q => IF_Regsxreg_file_287_port, QN => 
                           n_2568);
   IF_Regsxreg_file_regx24xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468294, Q => IF_Regsxreg_file_255_port, QN => 
                           n_2569);
   IF_Regsxreg_file_regx25xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468289, Q => IF_Regsxreg_file_223_port, QN => 
                           n_2570);
   IF_Regsxreg_file_regx26xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468284, Q => IF_Regsxreg_file_191_port, QN => 
                           n_2571);
   IF_Regsxreg_file_regx27xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468279, Q => IF_Regsxreg_file_159_port, QN => 
                           n_2572);
   IF_Regsxreg_file_regx28xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468274, Q => IF_Regsxreg_file_127_port, QN => 
                           n_2573);
   IF_Regsxreg_file_regx29xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468269, Q => IF_Regsxreg_file_95_port, QN => 
                           n_2574);
   IF_Regsxreg_file_regx30xx31x : DFF_X1 port map( D => IF_RegsxN691, CK => 
                           net2468264, Q => IF_Regsxreg_file_63_port, QN => 
                           n_2575);
   IF_RegsxRegsToCtl_port_contents2_regx31x : DFF_X1 port map( D => 
                           IF_RegsxN658, CK => net2468414, Q => 
                           RegsToCtl_port_contents2_31_port, QN => n_2576);
   IF_CPathxRegsToCtl_data_signal_contents2_regx31x : DFF_X1 port map( D => 
                           IF_CPathxN2155, CK => net2468199, Q => n_2577, QN =>
                           n6318);
   IF_CPathxCtlToMem_port_dataIn_regx31x : DFF_X1 port map( D => n6434, CK => 
                           net2468164, Q => CtlToMem_port_dataIn(31), QN => 
                           n_2578);
   IF_CPathxCtlToALU_port_reg2_contents_regx31x : DFF_X1 port map( D => n6579, 
                           CK => net2468224, Q => 
                           CtlToALU_port_reg2_contents_31_port, QN => n_2579);
   DP_OP_1698J95_122_4028xU33 : FA_X1 port map( A => IF_ALUxN112, B => n6378, 
                           CI => DP_OP_1698J95_122_4028xn68, CO => 
                           DP_OP_1698J95_122_4028xn32, S => C596xDATA2_0);
   DP_OP_1698J95_122_4028xU32 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn67
                           , B => IF_ALUxN113, CI => DP_OP_1698J95_122_4028xn32
                           , CO => DP_OP_1698J95_122_4028xn31, S => 
                           C596xDATA2_1);
   DP_OP_1698J95_122_4028xU31 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn66
                           , B => IF_ALUxN114, CI => DP_OP_1698J95_122_4028xn31
                           , CO => DP_OP_1698J95_122_4028xn30, S => 
                           C596xDATA2_2);
   DP_OP_1698J95_122_4028xU30 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn65
                           , B => IF_ALUxN115, CI => DP_OP_1698J95_122_4028xn30
                           , CO => DP_OP_1698J95_122_4028xn29, S => 
                           C596xDATA2_3);
   DP_OP_1698J95_122_4028xU29 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn64
                           , B => IF_ALUxN116, CI => DP_OP_1698J95_122_4028xn29
                           , CO => DP_OP_1698J95_122_4028xn28, S => 
                           C596xDATA2_4);
   DP_OP_1698J95_122_4028xU28 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn63
                           , B => IF_ALUxN117, CI => DP_OP_1698J95_122_4028xn28
                           , CO => DP_OP_1698J95_122_4028xn27, S => 
                           C596xDATA2_5);
   DP_OP_1698J95_122_4028xU27 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn62
                           , B => IF_ALUxN118, CI => DP_OP_1698J95_122_4028xn27
                           , CO => DP_OP_1698J95_122_4028xn26, S => 
                           C596xDATA2_6);
   DP_OP_1698J95_122_4028xU26 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn61
                           , B => IF_ALUxN119, CI => DP_OP_1698J95_122_4028xn26
                           , CO => DP_OP_1698J95_122_4028xn25, S => 
                           C596xDATA2_7);
   DP_OP_1698J95_122_4028xU25 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn60
                           , B => IF_ALUxN120, CI => DP_OP_1698J95_122_4028xn25
                           , CO => DP_OP_1698J95_122_4028xn24, S => 
                           C596xDATA2_8);
   DP_OP_1698J95_122_4028xU24 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn59
                           , B => IF_ALUxN121, CI => DP_OP_1698J95_122_4028xn24
                           , CO => DP_OP_1698J95_122_4028xn23, S => 
                           C596xDATA2_9);
   DP_OP_1698J95_122_4028xU23 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn58
                           , B => IF_ALUxN122, CI => DP_OP_1698J95_122_4028xn23
                           , CO => DP_OP_1698J95_122_4028xn22, S => 
                           C596xDATA2_10);
   DP_OP_1698J95_122_4028xU22 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn57
                           , B => IF_ALUxN123, CI => DP_OP_1698J95_122_4028xn22
                           , CO => DP_OP_1698J95_122_4028xn21, S => 
                           C596xDATA2_11);
   DP_OP_1698J95_122_4028xU21 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn56
                           , B => IF_ALUxN124, CI => DP_OP_1698J95_122_4028xn21
                           , CO => DP_OP_1698J95_122_4028xn20, S => 
                           C596xDATA2_12);
   DP_OP_1698J95_122_4028xU20 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn55
                           , B => IF_ALUxN125, CI => DP_OP_1698J95_122_4028xn20
                           , CO => DP_OP_1698J95_122_4028xn19, S => 
                           C596xDATA2_13);
   DP_OP_1698J95_122_4028xU19 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn54
                           , B => IF_ALUxN126, CI => DP_OP_1698J95_122_4028xn19
                           , CO => DP_OP_1698J95_122_4028xn18, S => 
                           C596xDATA2_14);
   DP_OP_1698J95_122_4028xU18 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn53
                           , B => IF_ALUxN127, CI => DP_OP_1698J95_122_4028xn18
                           , CO => DP_OP_1698J95_122_4028xn17, S => 
                           C596xDATA2_15);
   DP_OP_1698J95_122_4028xU17 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn52
                           , B => IF_ALUxN128, CI => DP_OP_1698J95_122_4028xn17
                           , CO => DP_OP_1698J95_122_4028xn16, S => 
                           C596xDATA2_16);
   DP_OP_1698J95_122_4028xU16 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn51
                           , B => IF_ALUxN129, CI => DP_OP_1698J95_122_4028xn16
                           , CO => DP_OP_1698J95_122_4028xn15, S => 
                           C596xDATA2_17);
   DP_OP_1698J95_122_4028xU15 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn50
                           , B => IF_ALUxN130, CI => DP_OP_1698J95_122_4028xn15
                           , CO => DP_OP_1698J95_122_4028xn14, S => 
                           C596xDATA2_18);
   DP_OP_1698J95_122_4028xU14 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn49
                           , B => IF_ALUxN131, CI => DP_OP_1698J95_122_4028xn14
                           , CO => DP_OP_1698J95_122_4028xn13, S => 
                           C596xDATA2_19);
   DP_OP_1698J95_122_4028xU13 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn48
                           , B => IF_ALUxN132, CI => DP_OP_1698J95_122_4028xn13
                           , CO => DP_OP_1698J95_122_4028xn12, S => 
                           C596xDATA2_20);
   DP_OP_1698J95_122_4028xU12 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn47
                           , B => IF_ALUxN133, CI => DP_OP_1698J95_122_4028xn12
                           , CO => DP_OP_1698J95_122_4028xn11, S => 
                           C596xDATA2_21);
   DP_OP_1698J95_122_4028xU11 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn46
                           , B => IF_ALUxN134, CI => DP_OP_1698J95_122_4028xn11
                           , CO => DP_OP_1698J95_122_4028xn10, S => 
                           C596xDATA2_22);
   DP_OP_1698J95_122_4028xU10 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn45
                           , B => IF_ALUxN135, CI => DP_OP_1698J95_122_4028xn10
                           , CO => DP_OP_1698J95_122_4028xn9, S => 
                           C596xDATA2_23);
   DP_OP_1698J95_122_4028xU9 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn44,
                           B => IF_ALUxN136, CI => DP_OP_1698J95_122_4028xn9, 
                           CO => DP_OP_1698J95_122_4028xn8, S => C596xDATA2_24)
                           ;
   DP_OP_1698J95_122_4028xU8 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn43,
                           B => IF_ALUxN137, CI => DP_OP_1698J95_122_4028xn8, 
                           CO => DP_OP_1698J95_122_4028xn7, S => C596xDATA2_25)
                           ;
   DP_OP_1698J95_122_4028xU7 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn42,
                           B => IF_ALUxN138, CI => DP_OP_1698J95_122_4028xn7, 
                           CO => DP_OP_1698J95_122_4028xn6, S => C596xDATA2_26)
                           ;
   DP_OP_1698J95_122_4028xU6 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn41,
                           B => IF_ALUxN139, CI => DP_OP_1698J95_122_4028xn6, 
                           CO => DP_OP_1698J95_122_4028xn5, S => C596xDATA2_27)
                           ;
   DP_OP_1698J95_122_4028xU5 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn40,
                           B => IF_ALUxN140, CI => DP_OP_1698J95_122_4028xn5, 
                           CO => DP_OP_1698J95_122_4028xn4, S => C596xDATA2_28)
                           ;
   DP_OP_1698J95_122_4028xU4 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn39,
                           B => IF_ALUxN141, CI => DP_OP_1698J95_122_4028xn4, 
                           CO => DP_OP_1698J95_122_4028xn3, S => C596xDATA2_29)
                           ;
   DP_OP_1698J95_122_4028xU3 : FA_X1 port map( A => DP_OP_1698J95_122_4028xn38,
                           B => IF_ALUxN142, CI => DP_OP_1698J95_122_4028xn3, 
                           CO => DP_OP_1698J95_122_4028xn2, S => C596xDATA2_30)
                           ;
   DP_OP_1703J95_125_7309xU33 : HA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn101, B => 
                           IF_CPathxDecToCtl_data_signal_imm_0_port, CO => 
                           DP_OP_1703J95_125_7309xn32, S => IF_CPathxN866);
   DP_OP_1703J95_125_7309xU32 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn102, B => 
                           IF_CPathxDecToCtl_data_signal_imm_1_port, CI => 
                           DP_OP_1703J95_125_7309xn32, CO => 
                           DP_OP_1703J95_125_7309xn31, S => IF_CPathxN867);
   DP_OP_1703J95_125_7309xU31 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn103, B => 
                           IF_CPathxDecToCtl_data_signal_imm_2_port, CI => 
                           DP_OP_1703J95_125_7309xn31, CO => 
                           DP_OP_1703J95_125_7309xn30, S => IF_CPathxN868);
   DP_OP_1703J95_125_7309xU30 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn104, B => 
                           IF_CPathxDecToCtl_data_signal_imm_3_port, CI => 
                           DP_OP_1703J95_125_7309xn30, CO => 
                           DP_OP_1703J95_125_7309xn29, S => IF_CPathxN869);
   DP_OP_1703J95_125_7309xU29 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn105, B => 
                           IF_CPathxDecToCtl_data_signal_imm_4_port, CI => 
                           DP_OP_1703J95_125_7309xn29, CO => 
                           DP_OP_1703J95_125_7309xn28, S => IF_CPathxN870);
   DP_OP_1703J95_125_7309xU28 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn106, B => 
                           IF_CPathxDecToCtl_data_signal_imm_5_port, CI => 
                           DP_OP_1703J95_125_7309xn28, CO => 
                           DP_OP_1703J95_125_7309xn27, S => IF_CPathxN871);
   DP_OP_1703J95_125_7309xU27 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn107, B => 
                           IF_CPathxDecToCtl_data_signal_imm_6_port, CI => 
                           DP_OP_1703J95_125_7309xn27, CO => 
                           DP_OP_1703J95_125_7309xn26, S => IF_CPathxN872);
   DP_OP_1703J95_125_7309xU26 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn108, B => 
                           IF_CPathxDecToCtl_data_signal_imm_7_port, CI => 
                           DP_OP_1703J95_125_7309xn26, CO => 
                           DP_OP_1703J95_125_7309xn25, S => IF_CPathxN873);
   DP_OP_1703J95_125_7309xU25 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn109, B => 
                           IF_CPathxDecToCtl_data_signal_imm_8_port, CI => 
                           DP_OP_1703J95_125_7309xn25, CO => 
                           DP_OP_1703J95_125_7309xn24, S => IF_CPathxN874);
   DP_OP_1703J95_125_7309xU24 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn110, B => 
                           IF_CPathxDecToCtl_data_signal_imm_9_port, CI => 
                           DP_OP_1703J95_125_7309xn24, CO => 
                           DP_OP_1703J95_125_7309xn23, S => IF_CPathxN875);
   DP_OP_1703J95_125_7309xU23 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn111, B => 
                           IF_CPathxDecToCtl_data_signal_imm_10_port, CI => 
                           DP_OP_1703J95_125_7309xn23, CO => 
                           DP_OP_1703J95_125_7309xn22, S => IF_CPathxN876);
   DP_OP_1703J95_125_7309xU22 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn112, B => 
                           IF_CPathxDecToCtl_data_signal_imm_11_port, CI => 
                           DP_OP_1703J95_125_7309xn22, CO => 
                           DP_OP_1703J95_125_7309xn21, S => IF_CPathxN877);
   DP_OP_1703J95_125_7309xU21 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn113, B => 
                           IF_CPathxDecToCtl_data_signal_imm_12_port, CI => 
                           DP_OP_1703J95_125_7309xn21, CO => 
                           DP_OP_1703J95_125_7309xn20, S => IF_CPathxN878);
   DP_OP_1703J95_125_7309xU20 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn114, B => 
                           IF_CPathxDecToCtl_data_signal_imm_13_port, CI => 
                           DP_OP_1703J95_125_7309xn20, CO => 
                           DP_OP_1703J95_125_7309xn19, S => IF_CPathxN879);
   DP_OP_1703J95_125_7309xU19 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn115, B => 
                           IF_CPathxDecToCtl_data_signal_imm_14_port, CI => 
                           DP_OP_1703J95_125_7309xn19, CO => 
                           DP_OP_1703J95_125_7309xn18, S => IF_CPathxN880);
   DP_OP_1703J95_125_7309xU18 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn116, B => 
                           IF_CPathxDecToCtl_data_signal_imm_15_port, CI => 
                           DP_OP_1703J95_125_7309xn18, CO => 
                           DP_OP_1703J95_125_7309xn17, S => IF_CPathxN881);
   DP_OP_1703J95_125_7309xU17 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn117, B => 
                           IF_CPathxDecToCtl_data_signal_imm_16_port, CI => 
                           DP_OP_1703J95_125_7309xn17, CO => 
                           DP_OP_1703J95_125_7309xn16, S => IF_CPathxN882);
   DP_OP_1703J95_125_7309xU16 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn118, B => 
                           IF_CPathxDecToCtl_data_signal_imm_17_port, CI => 
                           DP_OP_1703J95_125_7309xn16, CO => 
                           DP_OP_1703J95_125_7309xn15, S => IF_CPathxN883);
   DP_OP_1703J95_125_7309xU15 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn119, B => 
                           IF_CPathxDecToCtl_data_signal_imm_18_port, CI => 
                           DP_OP_1703J95_125_7309xn15, CO => 
                           DP_OP_1703J95_125_7309xn14, S => IF_CPathxN884);
   DP_OP_1703J95_125_7309xU14 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn120, B => 
                           IF_CPathxDecToCtl_data_signal_imm_19_port, CI => 
                           DP_OP_1703J95_125_7309xn14, CO => 
                           DP_OP_1703J95_125_7309xn13, S => IF_CPathxN885);
   DP_OP_1703J95_125_7309xU13 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn121, B => 
                           IF_CPathxDecToCtl_data_signal_imm_20_port, CI => 
                           DP_OP_1703J95_125_7309xn13, CO => 
                           DP_OP_1703J95_125_7309xn12, S => IF_CPathxN886);
   DP_OP_1703J95_125_7309xU12 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn122, B => 
                           IF_CPathxDecToCtl_data_signal_imm_21_port, CI => 
                           DP_OP_1703J95_125_7309xn12, CO => 
                           DP_OP_1703J95_125_7309xn11, S => IF_CPathxN887);
   DP_OP_1703J95_125_7309xU11 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn123, B => 
                           IF_CPathxDecToCtl_data_signal_imm_22_port, CI => 
                           DP_OP_1703J95_125_7309xn11, CO => 
                           DP_OP_1703J95_125_7309xn10, S => IF_CPathxN888);
   DP_OP_1703J95_125_7309xU10 : FA_X1 port map( A => 
                           DP_OP_1703J95_125_7309xn124, B => 
                           IF_CPathxDecToCtl_data_signal_imm_23_port, CI => 
                           DP_OP_1703J95_125_7309xn10, CO => 
                           DP_OP_1703J95_125_7309xn9, S => IF_CPathxN889);
   DP_OP_1703J95_125_7309xU9 : FA_X1 port map( A => DP_OP_1703J95_125_7309xn125
                           , B => IF_CPathxDecToCtl_data_signal_imm_24_port, CI
                           => DP_OP_1703J95_125_7309xn9, CO => 
                           DP_OP_1703J95_125_7309xn8, S => IF_CPathxN890);
   DP_OP_1703J95_125_7309xU8 : FA_X1 port map( A => DP_OP_1703J95_125_7309xn126
                           , B => IF_CPathxDecToCtl_data_signal_imm_25_port, CI
                           => DP_OP_1703J95_125_7309xn8, CO => 
                           DP_OP_1703J95_125_7309xn7, S => IF_CPathxN891);
   DP_OP_1703J95_125_7309xU7 : FA_X1 port map( A => DP_OP_1703J95_125_7309xn127
                           , B => IF_CPathxDecToCtl_data_signal_imm_26_port, CI
                           => DP_OP_1703J95_125_7309xn7, CO => 
                           DP_OP_1703J95_125_7309xn6, S => IF_CPathxN892);
   DP_OP_1703J95_125_7309xU6 : FA_X1 port map( A => DP_OP_1703J95_125_7309xn128
                           , B => IF_CPathxDecToCtl_data_signal_imm_27_port, CI
                           => DP_OP_1703J95_125_7309xn6, CO => 
                           DP_OP_1703J95_125_7309xn5, S => IF_CPathxN893);
   DP_OP_1703J95_125_7309xU5 : FA_X1 port map( A => DP_OP_1703J95_125_7309xn129
                           , B => IF_CPathxDecToCtl_data_signal_imm_28_port, CI
                           => DP_OP_1703J95_125_7309xn5, CO => 
                           DP_OP_1703J95_125_7309xn4, S => IF_CPathxN894);
   DP_OP_1703J95_125_7309xU4 : FA_X1 port map( A => DP_OP_1703J95_125_7309xn130
                           , B => IF_CPathxDecToCtl_data_signal_imm_29_port, CI
                           => DP_OP_1703J95_125_7309xn4, CO => 
                           DP_OP_1703J95_125_7309xn3, S => IF_CPathxN895);
   DP_OP_1703J95_125_7309xU3 : FA_X1 port map( A => DP_OP_1703J95_125_7309xn131
                           , B => IF_CPathxDecToCtl_data_signal_imm_30_port, CI
                           => DP_OP_1703J95_125_7309xn3, CO => 
                           DP_OP_1703J95_125_7309xn2, S => IF_CPathxN896);
   IF_DecoderxDecToCtl_port_encType_regx1x : DFF_X1 port map( D => 
                           IF_DecoderxN550, CK => net2468249, Q => 
                           DecToCtl_port_encType_1_port, QN => n6225);
   IF_DecoderxDecToCtl_port_instrType_regx2x : DFF_X1 port map( D => 
                           IF_DecoderxN587, CK => net2468249, Q => 
                           DecToCtl_port_instrType_2_port, QN => n6195);
   IF_DecoderxDecToCtl_port_instrType_regx4x : DFF_X1 port map( D => 
                           IF_DecoderxN589, CK => net2468249, Q => 
                           DecToCtl_port_instrType_4_port, QN => n6191);
   IF_CPathxCtlToALU_port_alu_fun_regx0x : DFF_X1 port map( D => IF_CPathxN1628
                           , CK => net2468149, Q => 
                           CtlToALU_port_alu_fun_0_port, QN => n6201);
   U3810 : NOR2_X4 port map( A1 => IF_CPathxwb_sel_signal_0_port, A2 => n4280, 
                           ZN => n4392);
   U3811 : OAI211_X2 port map( C1 => n3042, C2 => n3041, A => n3040, B => n3039
                           , ZN => n3113);
   U3812 : INV_X1 port map( A => rst, ZN => n4671);
   U3813 : CLKBUF_X1 port map( A => n4671, Z => n6180);
   U3814 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_22_port, A2 => n6180
                           , ZN => IF_RegsxN682);
   U3815 : CLKBUF_X1 port map( A => n4671, Z => n4547);
   U3816 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_20_port, A2 => n4547
                           , ZN => IF_RegsxN680);
   U3817 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_15_port, A2 => n6180
                           , ZN => IF_RegsxN675);
   U3818 : CLKBUF_X1 port map( A => n4671, Z => n4571);
   U3819 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_13_port, A2 => n4571
                           , ZN => IF_RegsxN673);
   U3820 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_11_port, A2 => n4547
                           , ZN => IF_RegsxN671);
   U3821 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_8_port, A2 => n6180,
                           ZN => IF_RegsxN668);
   U3822 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_23_port, A2 => n6180
                           , ZN => IF_RegsxN683);
   U3823 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_28_port, A2 => n6180
                           , ZN => IF_RegsxN688);
   U3824 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_16_port, A2 => n6180
                           , ZN => IF_RegsxN676);
   U3825 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_27_port, A2 => n4547
                           , ZN => IF_RegsxN687);
   U3826 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_12_port, A2 => n4547
                           , ZN => IF_RegsxN672);
   U3827 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_26_port, A2 => n4547
                           , ZN => IF_RegsxN686);
   U3828 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_10_port, A2 => n6180
                           , ZN => IF_RegsxN670);
   U3829 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_29_port, A2 => n4547
                           , ZN => IF_RegsxN689);
   U3830 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_0_port, A2 => n6180,
                           ZN => IF_RegsxN660);
   U3831 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_7_port, A2 => n6180,
                           ZN => IF_RegsxN667);
   U3832 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_5_port, A2 => n6180,
                           ZN => IF_RegsxN665);
   U3833 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_1_port, A2 => n6180,
                           ZN => IF_RegsxN661);
   U3834 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_3_port, A2 => n6180,
                           ZN => IF_RegsxN663);
   U3835 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_30_port, A2 => n4547
                           , ZN => IF_RegsxN690);
   U3836 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_31_port, A2 => n4571
                           , ZN => IF_RegsxN691);
   U3837 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_6_port, A2 => n6180,
                           ZN => IF_RegsxN666);
   U3838 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_9_port, A2 => n4547,
                           ZN => IF_RegsxN669);
   U3839 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_25_port, A2 => n6180
                           , ZN => IF_RegsxN685);
   U3840 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_18_port, A2 => n4547
                           , ZN => IF_RegsxN678);
   U3841 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_21_port, A2 => n4547
                           , ZN => IF_RegsxN681);
   U3842 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_19_port, A2 => n6180
                           , ZN => IF_RegsxN679);
   U3843 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_24_port, A2 => n4547
                           , ZN => IF_RegsxN684);
   U3844 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_17_port, A2 => n4547
                           , ZN => IF_RegsxN677);
   U3845 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_2_port, A2 => n6180,
                           ZN => IF_RegsxN662);
   U3846 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_14_port, A2 => n4547
                           , ZN => IF_RegsxN674);
   U3847 : AND2_X1 port map( A1 => CtlToRegs_port_dst_data_4_port, A2 => n6180,
                           ZN => IF_RegsxN664);
   U3848 : NOR2_X1 port map( A1 => n6193, A2 => CtlToALU_port_alu_fun_2_port, 
                           ZN => n3263);
   U3849 : INV_X1 port map( A => n3263, ZN => n2954);
   U3850 : NOR3_X1 port map( A1 => n2954, A2 => CtlToALU_port_alu_fun_1_port, 
                           A3 => n6201, ZN => n3276);
   U3851 : CLKBUF_X2 port map( A => n3276, Z => n6378);
   U3852 : AND2_X1 port map( A1 => n6203, A2 => CtlToALU_port_op1_sel_0_port, 
                           ZN => n3207);
   U3853 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_24_port, 
                           ZN => n2957);
   U3854 : AND2_X1 port map( A1 => n6242, A2 => CtlToALU_port_op1_sel_1_port, 
                           ZN => n3242);
   U3855 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_24_port, ZN => n2956);
   U3856 : NOR2_X1 port map( A1 => CtlToALU_port_op1_sel_1_port, A2 => 
                           CtlToALU_port_op1_sel_0_port, ZN => n3208);
   U3857 : CLKBUF_X1 port map( A => n3208, Z => n3258);
   U3858 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_24_port, ZN 
                           => n2955);
   U3859 : NAND3_X1 port map( A1 => n2957, A2 => n2956, A3 => n2955, ZN => 
                           IF_ALUxN136);
   U3860 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_30_port, 
                           ZN => n2960);
   U3861 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_30_port, ZN => n2959);
   U3862 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_30_port, ZN 
                           => n2958);
   U3863 : NAND3_X1 port map( A1 => n2960, A2 => n2959, A3 => n2958, ZN => 
                           IF_ALUxN142);
   U3864 : AND2_X1 port map( A1 => n6241, A2 => CtlToALU_port_op2_sel_1_port, 
                           ZN => n3932);
   U3865 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_30_port, ZN => n2963);
   U3866 : AND2_X1 port map( A1 => n6202, A2 => CtlToALU_port_op2_sel_0_port, 
                           ZN => n3931);
   U3867 : CLKBUF_X1 port map( A => n3931, Z => n3023);
   U3868 : NAND2_X1 port map( A1 => n3023, A2 => CtlToALU_port_pc_reg_30_port, 
                           ZN => n2962);
   U3869 : NOR2_X1 port map( A1 => CtlToALU_port_op2_sel_1_port, A2 => 
                           CtlToALU_port_op2_sel_0_port, ZN => n3018);
   U3870 : CLKBUF_X1 port map( A => n3018, Z => n3930);
   U3871 : NAND2_X1 port map( A1 => n3930, A2 => CtlToALU_port_imm_30_port, ZN 
                           => n2961);
   U3872 : NAND3_X1 port map( A1 => n2963, A2 => n2962, A3 => n2961, ZN => 
                           n4040);
   U3873 : XOR2_X1 port map( A => n6378, B => n4040, Z => 
                           DP_OP_1698J95_122_4028xn38);
   U3874 : AOI222_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_29_port, B1 => n3931, B2
                           => CtlToALU_port_pc_reg_29_port, C1 => n3930, C2 => 
                           CtlToALU_port_imm_29_port, ZN => n3840);
   U3875 : INV_X1 port map( A => n3840, ZN => n3829);
   U3876 : XOR2_X1 port map( A => n6378, B => n3829, Z => 
                           DP_OP_1698J95_122_4028xn39);
   U3877 : AOI222_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_28_port, B1 => n3931, B2
                           => CtlToALU_port_pc_reg_28_port, C1 => n3930, C2 => 
                           CtlToALU_port_imm_28_port, ZN => n3846);
   U3878 : INV_X1 port map( A => n3846, ZN => n4032);
   U3879 : XOR2_X1 port map( A => n6378, B => n4032, Z => 
                           DP_OP_1698J95_122_4028xn40);
   U3880 : CLKBUF_X1 port map( A => n3932, Z => n3022);
   U3881 : NAND2_X1 port map( A1 => n3022, A2 => 
                           CtlToALU_port_reg2_contents_27_port, ZN => n2966);
   U3882 : NAND2_X1 port map( A1 => n3931, A2 => CtlToALU_port_pc_reg_27_port, 
                           ZN => n2965);
   U3883 : NAND2_X1 port map( A1 => n3930, A2 => CtlToALU_port_imm_27_port, ZN 
                           => n2964);
   U3884 : NAND3_X1 port map( A1 => n2966, A2 => n2965, A3 => n2964, ZN => 
                           n3762);
   U3885 : XOR2_X1 port map( A => n6378, B => n3762, Z => 
                           DP_OP_1698J95_122_4028xn41);
   U3886 : NAND2_X1 port map( A1 => n3022, A2 => 
                           CtlToALU_port_reg2_contents_26_port, ZN => n2969);
   U3887 : NAND2_X1 port map( A1 => n3931, A2 => CtlToALU_port_pc_reg_26_port, 
                           ZN => n2968);
   U3888 : NAND2_X1 port map( A1 => n3930, A2 => CtlToALU_port_imm_26_port, ZN 
                           => n2967);
   U3889 : NAND3_X1 port map( A1 => n2969, A2 => n2968, A3 => n2967, ZN => 
                           n3788);
   U3890 : XOR2_X1 port map( A => n6378, B => n3788, Z => 
                           DP_OP_1698J95_122_4028xn42);
   U3891 : AOI222_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_25_port, B1 => n3931, B2
                           => CtlToALU_port_pc_reg_25_port, C1 => n3930, C2 => 
                           CtlToALU_port_imm_25_port, ZN => n3331);
   U3892 : INV_X1 port map( A => n3331, ZN => n3319);
   U3893 : XOR2_X1 port map( A => n6378, B => n3319, Z => 
                           DP_OP_1698J95_122_4028xn43);
   U3894 : AOI222_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_24_port, B1 => n3931, B2
                           => CtlToALU_port_pc_reg_24_port, C1 => n3930, C2 => 
                           CtlToALU_port_imm_24_port, ZN => n4020);
   U3895 : INV_X1 port map( A => n4020, ZN => n3881);
   U3896 : XOR2_X1 port map( A => n6378, B => n3881, Z => 
                           DP_OP_1698J95_122_4028xn44);
   U3897 : AOI222_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_23_port, B1 => n3931, B2
                           => CtlToALU_port_pc_reg_23_port, C1 => n3930, C2 => 
                           CtlToALU_port_imm_23_port, ZN => n3680);
   U3898 : INV_X1 port map( A => n3680, ZN => n3669);
   U3899 : XOR2_X1 port map( A => n3276, B => n3669, Z => 
                           DP_OP_1698J95_122_4028xn45);
   U3900 : NAND2_X1 port map( A1 => n3022, A2 => 
                           CtlToALU_port_reg2_contents_22_port, ZN => n2972);
   U3901 : NAND2_X1 port map( A1 => n3931, A2 => CtlToALU_port_pc_reg_22_port, 
                           ZN => n2971);
   U3902 : NAND2_X1 port map( A1 => n3930, A2 => CtlToALU_port_imm_22_port, ZN 
                           => n2970);
   U3903 : NAND3_X1 port map( A1 => n2972, A2 => n2971, A3 => n2970, ZN => 
                           n3688);
   U3904 : XOR2_X1 port map( A => n3276, B => n3688, Z => 
                           DP_OP_1698J95_122_4028xn46);
   U3905 : NAND2_X1 port map( A1 => n3022, A2 => 
                           CtlToALU_port_reg2_contents_21_port, ZN => n2975);
   U3906 : NAND2_X1 port map( A1 => n3931, A2 => CtlToALU_port_pc_reg_21_port, 
                           ZN => n2974);
   U3907 : NAND2_X1 port map( A1 => n3930, A2 => CtlToALU_port_imm_21_port, ZN 
                           => n2973);
   U3908 : NAND3_X1 port map( A1 => n2975, A2 => n2974, A3 => n2973, ZN => 
                           n3532);
   U3909 : XOR2_X1 port map( A => n3276, B => n3532, Z => 
                           DP_OP_1698J95_122_4028xn47);
   U3910 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_20_port, ZN => n2978);
   U3911 : NAND2_X1 port map( A1 => n3023, A2 => CtlToALU_port_pc_reg_20_port, 
                           ZN => n2977);
   U3912 : NAND2_X1 port map( A1 => n3930, A2 => CtlToALU_port_imm_20_port, ZN 
                           => n2976);
   U3913 : NAND3_X1 port map( A1 => n2978, A2 => n2977, A3 => n2976, ZN => 
                           n3709);
   U3914 : XOR2_X1 port map( A => n3276, B => n3709, Z => 
                           DP_OP_1698J95_122_4028xn48);
   U3915 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_19_port, ZN => n2981);
   U3916 : NAND2_X1 port map( A1 => n3023, A2 => CtlToALU_port_pc_reg_19_port, 
                           ZN => n2980);
   U3917 : NAND2_X1 port map( A1 => n3930, A2 => CtlToALU_port_imm_19_port, ZN 
                           => n2979);
   U3918 : NAND3_X1 port map( A1 => n2981, A2 => n2980, A3 => n2979, ZN => 
                           n4007);
   U3919 : XOR2_X1 port map( A => n6378, B => n4007, Z => 
                           DP_OP_1698J95_122_4028xn49);
   U3920 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_18_port, ZN => n2984);
   U3921 : NAND2_X1 port map( A1 => n3023, A2 => CtlToALU_port_pc_reg_18_port, 
                           ZN => n2983);
   U3922 : NAND2_X1 port map( A1 => n3930, A2 => CtlToALU_port_imm_18_port, ZN 
                           => n2982);
   U3923 : NAND3_X1 port map( A1 => n2984, A2 => n2983, A3 => n2982, ZN => 
                           n3996);
   U3924 : XOR2_X1 port map( A => n6378, B => n3996, Z => 
                           DP_OP_1698J95_122_4028xn50);
   U3925 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_17_port, ZN => n2987);
   U3926 : NAND2_X1 port map( A1 => n3023, A2 => CtlToALU_port_pc_reg_17_port, 
                           ZN => n2986);
   U3927 : NAND2_X1 port map( A1 => n3930, A2 => CtlToALU_port_imm_17_port, ZN 
                           => n2985);
   U3928 : NAND3_X1 port map( A1 => n2987, A2 => n2986, A3 => n2985, ZN => 
                           n4001);
   U3929 : XOR2_X1 port map( A => n6378, B => n4001, Z => 
                           DP_OP_1698J95_122_4028xn51);
   U3930 : AOI222_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_16_port, B1 => n3931, B2
                           => CtlToALU_port_pc_reg_16_port, C1 => n3930, C2 => 
                           CtlToALU_port_imm_16_port, ZN => n3919);
   U3931 : INV_X1 port map( A => n3919, ZN => n4003);
   U3932 : XOR2_X1 port map( A => n6378, B => n4003, Z => 
                           DP_OP_1698J95_122_4028xn52);
   U3933 : NAND2_X1 port map( A1 => n3022, A2 => 
                           CtlToALU_port_reg2_contents_15_port, ZN => n2990);
   U3934 : NAND2_X1 port map( A1 => n3931, A2 => CtlToALU_port_pc_reg_15_port, 
                           ZN => n2989);
   U3935 : NAND2_X1 port map( A1 => n3930, A2 => CtlToALU_port_imm_15_port, ZN 
                           => n2988);
   U3936 : NAND3_X1 port map( A1 => n2990, A2 => n2989, A3 => n2988, ZN => 
                           n3944);
   U3937 : XOR2_X1 port map( A => n6378, B => n3944, Z => 
                           DP_OP_1698J95_122_4028xn53);
   U3938 : NAND2_X1 port map( A1 => n3022, A2 => 
                           CtlToALU_port_reg2_contents_14_port, ZN => n2993);
   U3939 : NAND2_X1 port map( A1 => n3931, A2 => CtlToALU_port_pc_reg_14_port, 
                           ZN => n2992);
   U3940 : NAND2_X1 port map( A1 => n3930, A2 => CtlToALU_port_imm_14_port, ZN 
                           => n2991);
   U3941 : NAND3_X1 port map( A1 => n2993, A2 => n2992, A3 => n2991, ZN => 
                           n3942);
   U3942 : XOR2_X1 port map( A => n6378, B => n3942, Z => 
                           DP_OP_1698J95_122_4028xn54);
   U3943 : AOI222_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_13_port, B1 => n3931, B2
                           => CtlToALU_port_pc_reg_13_port, C1 => n3018, C2 => 
                           CtlToALU_port_imm_13_port, ZN => n3618);
   U3944 : INV_X1 port map( A => n3618, ZN => n3610);
   U3945 : XOR2_X1 port map( A => n6378, B => n3610, Z => 
                           DP_OP_1698J95_122_4028xn55);
   U3946 : AOI222_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_12_port, B1 => n3931, B2
                           => CtlToALU_port_pc_reg_12_port, C1 => n3018, C2 => 
                           CtlToALU_port_imm_12_port, ZN => n3752);
   U3947 : INV_X1 port map( A => n3752, ZN => n3739);
   U3948 : XOR2_X1 port map( A => n6378, B => n3739, Z => 
                           DP_OP_1698J95_122_4028xn56);
   U3949 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_11_port, ZN => n2996);
   U3950 : NAND2_X1 port map( A1 => n3023, A2 => CtlToALU_port_pc_reg_11_port, 
                           ZN => n2995);
   U3951 : NAND2_X1 port map( A1 => n3018, A2 => CtlToALU_port_imm_11_port, ZN 
                           => n2994);
   U3952 : NAND3_X1 port map( A1 => n2996, A2 => n2995, A3 => n2994, ZN => 
                           n3631);
   U3953 : XOR2_X1 port map( A => n6378, B => n3631, Z => 
                           DP_OP_1698J95_122_4028xn57);
   U3954 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_10_port, ZN => n2999);
   U3955 : NAND2_X1 port map( A1 => n3023, A2 => CtlToALU_port_pc_reg_10_port, 
                           ZN => n2998);
   U3956 : NAND2_X1 port map( A1 => n3018, A2 => CtlToALU_port_imm_10_port, ZN 
                           => n2997);
   U3957 : NAND3_X1 port map( A1 => n2999, A2 => n2998, A3 => n2997, ZN => 
                           n3982);
   U3958 : XOR2_X1 port map( A => n6378, B => n3982, Z => 
                           DP_OP_1698J95_122_4028xn58);
   U3959 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_9_port, ZN => n3002);
   U3960 : NAND2_X1 port map( A1 => n3931, A2 => CtlToALU_port_pc_reg_9_port, 
                           ZN => n3001);
   U3961 : NAND2_X1 port map( A1 => n3018, A2 => CtlToALU_port_imm_9_port, ZN 
                           => n3000);
   U3962 : NAND3_X1 port map( A1 => n3002, A2 => n3001, A3 => n3000, ZN => 
                           n3949);
   U3963 : XOR2_X1 port map( A => n6378, B => n3949, Z => 
                           DP_OP_1698J95_122_4028xn59);
   U3964 : NAND2_X1 port map( A1 => n3022, A2 => 
                           CtlToALU_port_reg2_contents_8_port, ZN => n3005);
   U3965 : NAND2_X1 port map( A1 => n3931, A2 => CtlToALU_port_pc_reg_8_port, 
                           ZN => n3004);
   U3966 : NAND2_X1 port map( A1 => n3018, A2 => CtlToALU_port_imm_8_port, ZN 
                           => n3003);
   U3967 : NAND3_X1 port map( A1 => n3005, A2 => n3004, A3 => n3003, ZN => 
                           n3951);
   U3968 : XOR2_X1 port map( A => n6378, B => n3951, Z => 
                           DP_OP_1698J95_122_4028xn60);
   U3969 : AOI222_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_7_port, B1 => n3931, B2 
                           => CtlToALU_port_pc_reg_7_port, C1 => n3930, C2 => 
                           CtlToALU_port_imm_7_port, ZN => n3361);
   U3970 : INV_X1 port map( A => n3361, ZN => n3975);
   U3971 : XOR2_X1 port map( A => n6378, B => n3975, Z => 
                           DP_OP_1698J95_122_4028xn61);
   U3972 : AOI222_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_6_port, B1 => n3931, B2 
                           => CtlToALU_port_pc_reg_6_port, C1 => n3018, C2 => 
                           CtlToALU_port_imm_6_port, ZN => n3298);
   U3973 : INV_X1 port map( A => n3298, ZN => n3965);
   U3974 : XOR2_X1 port map( A => n6378, B => n3965, Z => 
                           DP_OP_1698J95_122_4028xn62);
   U3975 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_5_port, ZN => n3008);
   U3976 : NAND2_X1 port map( A1 => n3023, A2 => CtlToALU_port_pc_reg_5_port, 
                           ZN => n3007);
   U3977 : NAND2_X1 port map( A1 => n3018, A2 => CtlToALU_port_imm_5_port, ZN 
                           => n3006);
   U3978 : NAND3_X1 port map( A1 => n3008, A2 => n3007, A3 => n3006, ZN => 
                           n3967);
   U3979 : XOR2_X1 port map( A => n6378, B => n3967, Z => 
                           DP_OP_1698J95_122_4028xn63);
   U3980 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_4_port, ZN => n3011);
   U3981 : NAND2_X1 port map( A1 => n3023, A2 => CtlToALU_port_pc_reg_4_port, 
                           ZN => n3010);
   U3982 : NAND2_X1 port map( A1 => n3018, A2 => CtlToALU_port_imm_4_port, ZN 
                           => n3009);
   U3983 : NAND3_X1 port map( A1 => n3011, A2 => n3010, A3 => n3009, ZN => 
                           n3271);
   U3984 : XOR2_X1 port map( A => n6378, B => n3271, Z => 
                           DP_OP_1698J95_122_4028xn64);
   U3985 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_3_port, ZN => n3014);
   U3986 : NAND2_X1 port map( A1 => n3023, A2 => CtlToALU_port_pc_reg_3_port, 
                           ZN => n3013);
   U3987 : NAND2_X1 port map( A1 => n3018, A2 => CtlToALU_port_imm_3_port, ZN 
                           => n3012);
   U3988 : NAND3_X1 port map( A1 => n3014, A2 => n3013, A3 => n3012, ZN => 
                           n3782);
   U3989 : INV_X1 port map( A => n3782, ZN => n3866);
   U3990 : INV_X1 port map( A => n3866, ZN => n4056);
   U3991 : XOR2_X1 port map( A => n6378, B => n4056, Z => 
                           DP_OP_1698J95_122_4028xn65);
   U3992 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_2_port, ZN => n3017);
   U3993 : NAND2_X1 port map( A1 => n3023, A2 => CtlToALU_port_pc_reg_2_port, 
                           ZN => n3016);
   U3994 : NAND2_X1 port map( A1 => n3018, A2 => CtlToALU_port_imm_2_port, ZN 
                           => n3015);
   U3995 : NAND3_X1 port map( A1 => n3017, A2 => n3016, A3 => n3015, ZN => 
                           n3875);
   U3996 : XOR2_X1 port map( A => n6378, B => n3875, Z => 
                           DP_OP_1698J95_122_4028xn66);
   U3997 : NAND2_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_1_port, ZN => n3021);
   U3998 : NAND2_X1 port map( A1 => n3023, A2 => CtlToALU_port_pc_reg_1_port, 
                           ZN => n3020);
   U3999 : NAND2_X1 port map( A1 => n3018, A2 => CtlToALU_port_imm_1_port, ZN 
                           => n3019);
   U4000 : NAND3_X1 port map( A1 => n3021, A2 => n3020, A3 => n3019, ZN => 
                           n4118);
   U4001 : XOR2_X1 port map( A => n6378, B => n4118, Z => 
                           DP_OP_1698J95_122_4028xn67);
   U4002 : AOI222_X1 port map( A1 => CtlToALU_port_pc_reg_0_port, A2 => n3023, 
                           B1 => n3022, B2 => 
                           CtlToALU_port_reg2_contents_0_port, C1 => n3930, C2 
                           => CtlToALU_port_imm_0_port, ZN => n3024);
   U4003 : INV_X1 port map( A => n3024, ZN => n3487);
   U4004 : INV_X1 port map( A => n3487, ZN => n4045);
   U4005 : INV_X2 port map( A => n4045, ZN => n4116);
   U4006 : XOR2_X1 port map( A => n6378, B => n4116, Z => 
                           DP_OP_1698J95_122_4028xn68);
   U4007 : CLKBUF_X1 port map( A => n4671, Z => n4546);
   U4008 : AND2_X1 port map( A1 => n4546, A2 => DecToCtl_port_imm_0_port, ZN =>
                           IF_CPathxN2158);
   U4009 : AND2_X1 port map( A1 => n4546, A2 => DecToCtl_port_imm_1_port, ZN =>
                           IF_CPathxN2159);
   U4010 : AND2_X1 port map( A1 => n4546, A2 => DecToCtl_port_imm_2_port, ZN =>
                           IF_CPathxN2160);
   U4011 : NOR2_X1 port map( A1 => rst, A2 => n6224, ZN => IF_CPathxN2161);
   U4012 : AND2_X1 port map( A1 => n4546, A2 => DecToCtl_port_imm_4_port, ZN =>
                           IF_CPathxN2162);
   U4013 : NOR2_X1 port map( A1 => rst, A2 => n6373, ZN => IF_CPathxN2090);
   U4014 : NOR2_X1 port map( A1 => rst, A2 => n6374, ZN => IF_CPathxN2096);
   U4015 : NOR2_X1 port map( A1 => rst, A2 => n6375, ZN => IF_CPathxN2094);
   U4016 : NOR2_X1 port map( A1 => rst, A2 => n6376, ZN => IF_CPathxN2095);
   U4017 : NOR2_X1 port map( A1 => rst, A2 => n6377, ZN => IF_CPathxN2092);
   U4018 : AND2_X1 port map( A1 => 
                           IF_CPathxDecToCtl_data_signal_instrType_0_port, A2 
                           => IF_CPathxDecToCtl_data_signal_instrType_1_port, 
                           ZN => n3043);
   U4019 : OR4_X1 port map( A1 => ALUtoCtl_port_29_port, A2 => 
                           ALUtoCtl_port_28_port, A3 => ALUtoCtl_port_27_port, 
                           A4 => ALUtoCtl_port_26_port, ZN => n3025);
   U4020 : NOR4_X1 port map( A1 => ALUtoCtl_port_1_port, A2 => 
                           ALUtoCtl_port_31_port, A3 => ALUtoCtl_port_30_port, 
                           A4 => n3025, ZN => n3033);
   U4021 : NOR4_X1 port map( A1 => ALUtoCtl_port_21_port, A2 => 
                           ALUtoCtl_port_20_port, A3 => ALUtoCtl_port_19_port, 
                           A4 => ALUtoCtl_port_18_port, ZN => n3032);
   U4022 : NOR4_X1 port map( A1 => ALUtoCtl_port_25_port, A2 => 
                           ALUtoCtl_port_24_port, A3 => ALUtoCtl_port_23_port, 
                           A4 => ALUtoCtl_port_22_port, ZN => n3031);
   U4023 : NOR4_X1 port map( A1 => ALUtoCtl_port_13_port, A2 => 
                           ALUtoCtl_port_12_port, A3 => ALUtoCtl_port_11_port, 
                           A4 => ALUtoCtl_port_10_port, ZN => n3029);
   U4024 : NOR4_X1 port map( A1 => ALUtoCtl_port_17_port, A2 => 
                           ALUtoCtl_port_16_port, A3 => ALUtoCtl_port_15_port, 
                           A4 => ALUtoCtl_port_14_port, ZN => n3028);
   U4025 : NOR4_X1 port map( A1 => ALUtoCtl_port_5_port, A2 => 
                           ALUtoCtl_port_4_port, A3 => ALUtoCtl_port_3_port, A4
                           => ALUtoCtl_port_2_port, ZN => n3027);
   U4026 : NOR4_X1 port map( A1 => ALUtoCtl_port_9_port, A2 => 
                           ALUtoCtl_port_8_port, A3 => ALUtoCtl_port_7_port, A4
                           => ALUtoCtl_port_6_port, ZN => n3026);
   U4027 : AND4_X1 port map( A1 => n3029, A2 => n3028, A3 => n3027, A4 => n3026
                           , ZN => n3030);
   U4028 : NAND4_X1 port map( A1 => n3033, A2 => n3032, A3 => n3031, A4 => 
                           n3030, ZN => n3037);
   U4029 : INV_X1 port map( A => n3037, ZN => n3035);
   U4030 : OAI21_X1 port map( B1 => 
                           IF_CPathxDecToCtl_data_signal_instrType_0_port, B2 
                           => n3035, A => IF_CPathxbr_en_signal, ZN => n3034);
   U4031 : AOI21_X1 port map( B1 => n3035, B2 => n6238, A => n3034, ZN => n3042
                           );
   U4032 : NAND2_X1 port map( A1 => n6240, A2 => 
                           IF_CPathxDecToCtl_data_signal_instrType_2_port, ZN 
                           => n3041);
   U4033 : NOR3_X1 port map( A1 => n6239, A2 => 
                           IF_CPathxDecToCtl_data_signal_instrType_4_port, A3 
                           => IF_CPathxDecToCtl_data_signal_instrType_5_port, 
                           ZN => n3040);
   U4034 : OAI21_X1 port map( B1 => n3043, B2 => n6238, A => 
                           IF_CPathxbr_en_signal, ZN => n3036);
   U4035 : AOI211_X1 port map( C1 => n3043, C2 => n6238, A => n3037, B => n3036
                           , ZN => n3038);
   U4036 : OR2_X1 port map( A1 => n3038, A2 => 
                           IF_CPathxDecToCtl_data_signal_instrType_2_port, ZN 
                           => n3039);
   U4037 : AOI21_X1 port map( B1 => 
                           IF_CPathxDecToCtl_data_signal_instrType_2_port, B2 
                           => n3043, A => n3113, ZN => n3093);
   U4038 : CLKBUF_X1 port map( A => n3093, Z => n3112);
   U4039 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_31_port, B 
                           => IF_CPathxpc_reg_signal_31_port, S => n3112, Z => 
                           n3044);
   U4040 : XOR2_X1 port map( A => n3044, B => 
                           IF_CPathxDecToCtl_data_signal_imm_31_port, Z => 
                           n3045);
   U4041 : XOR2_X1 port map( A => DP_OP_1703J95_125_7309xn2, B => n3045, Z => 
                           n3048);
   U4042 : INV_X1 port map( A => n3113, ZN => n3115);
   U4043 : CLKBUF_X1 port map( A => n3115, Z => n3111);
   U4044 : NOR2_X1 port map( A1 => n6204, A2 => n6245, ZN => n3108);
   U4045 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_4_port, A2 => n3108,
                           ZN => n3105);
   U4046 : NOR2_X1 port map( A1 => n6243, A2 => n3105, ZN => n3103);
   U4047 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_6_port, A2 => n3103,
                           ZN => n3101);
   U4048 : NOR2_X1 port map( A1 => n6244, A2 => n3101, ZN => n3098);
   U4049 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_8_port, A2 => n3098,
                           ZN => n3096);
   U4050 : NOR2_X1 port map( A1 => n6247, A2 => n3096, ZN => n3094);
   U4051 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_10_port, A2 => n3094
                           , ZN => n3091);
   U4052 : NOR2_X1 port map( A1 => n6248, A2 => n3091, ZN => n3088);
   U4053 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_12_port, A2 => n3088
                           , ZN => n3086);
   U4054 : NOR2_X1 port map( A1 => n6249, A2 => n3086, ZN => n3084);
   U4055 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_14_port, A2 => n3084
                           , ZN => n3082);
   U4056 : NOR2_X1 port map( A1 => n6250, A2 => n3082, ZN => n3080);
   U4057 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_16_port, A2 => n3080
                           , ZN => n3078);
   U4058 : NOR2_X1 port map( A1 => n6251, A2 => n3078, ZN => n3076);
   U4059 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_18_port, A2 => n3076
                           , ZN => n3074);
   U4060 : NOR2_X1 port map( A1 => n6252, A2 => n3074, ZN => n3072);
   U4061 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_20_port, A2 => n3072
                           , ZN => n3070);
   U4062 : NOR2_X1 port map( A1 => n6253, A2 => n3070, ZN => n3068);
   U4063 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_22_port, A2 => n3068
                           , ZN => n3066);
   U4064 : NOR2_X1 port map( A1 => n6254, A2 => n3066, ZN => n3064);
   U4065 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_24_port, A2 => n3064
                           , ZN => n3062);
   U4066 : NOR2_X1 port map( A1 => n6255, A2 => n3062, ZN => n3060);
   U4067 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_26_port, A2 => n3060
                           , ZN => n3058);
   U4068 : NOR2_X1 port map( A1 => n6262, A2 => n3058, ZN => n3056);
   U4069 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_28_port, A2 => n3056
                           , ZN => n3054);
   U4070 : NOR2_X1 port map( A1 => n6263, A2 => n3054, ZN => n3052);
   U4071 : NAND2_X1 port map( A1 => IF_CPathxpc_reg_signal_30_port, A2 => n3052
                           , ZN => n3046);
   U4072 : XNOR2_X1 port map( A => IF_CPathxpc_reg_signal_31_port, B => n3046, 
                           ZN => n4393);
   U4073 : AND2_X1 port map( A1 => n3113, A2 => n4393, ZN => n3047);
   U4074 : AOI21_X1 port map( B1 => n3048, B2 => n3111, A => n3047, ZN => n3250
                           );
   U4075 : NOR2_X1 port map( A1 => n6196, A2 => rst, ZN => n4279);
   U4076 : INV_X1 port map( A => n4279, ZN => n3100);
   U4077 : NAND2_X1 port map( A1 => n4571, A2 => n6196, ZN => n4281);
   U4078 : INV_X1 port map( A => n4281, ZN => n3090);
   U4079 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_31_port, ZN => n3248);
   U4080 : OAI21_X1 port map( B1 => n3250, B2 => n3100, A => n3248, ZN => n6506
                           );
   U4081 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_31_port, ZN => n6405);
   U4082 : INV_X1 port map( A => n3052, ZN => n3049);
   U4083 : XOR2_X1 port map( A => IF_CPathxpc_reg_signal_30_port, B => n3049, Z
                           => n4389);
   U4084 : NAND2_X1 port map( A1 => n3113, A2 => n4389, ZN => n3050);
   U4085 : OAI21_X1 port map( B1 => IF_CPathxN896, B2 => n3113, A => n3050, ZN 
                           => n3254);
   U4086 : NOR2_X1 port map( A1 => rst, A2 => n3254, ZN => n6423);
   U4087 : INV_X1 port map( A => n6423, ZN => n3051);
   U4088 : CLKBUF_X1 port map( A => n3090, Z => n4181);
   U4089 : NAND2_X1 port map( A1 => n4181, A2 => 
                           IF_CPathxpc_next_signal_30_port, ZN => n3252);
   U4090 : OAI21_X1 port map( B1 => n6196, B2 => n3051, A => n3252, ZN => n6507
                           );
   U4091 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_30_port, ZN => n6404);
   U4092 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_30_port, B 
                           => IF_CPathxpc_reg_signal_30_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn131);
   U4093 : AOI21_X1 port map( B1 => n6263, B2 => n3054, A => n3052, ZN => n4296
                           );
   U4094 : AND2_X1 port map( A1 => n3113, A2 => n4296, ZN => n3053);
   U4095 : AOI21_X1 port map( B1 => IF_CPathxN895, B2 => n3111, A => n3053, ZN 
                           => n4085);
   U4096 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_29_port, ZN => n3821);
   U4097 : OAI21_X1 port map( B1 => n4085, B2 => n3100, A => n3821, ZN => n6508
                           );
   U4098 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_29_port, ZN => n6403);
   U4099 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_29_port, B 
                           => IF_CPathxpc_reg_signal_29_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn130);
   U4100 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_28_port, B2 => n3056
                           , A => n3054, ZN => n4292);
   U4101 : NOR2_X1 port map( A1 => n3115, A2 => n4292, ZN => n3055);
   U4102 : AOI21_X1 port map( B1 => IF_CPathxN894, B2 => n3111, A => n3055, ZN 
                           => n4086);
   U4103 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_28_port, ZN => n3844);
   U4104 : OAI21_X1 port map( B1 => n4086, B2 => n3100, A => n3844, ZN => n6509
                           );
   U4105 : CLKBUF_X1 port map( A => n4671, Z => n4545);
   U4106 : AND2_X1 port map( A1 => n4545, A2 => 
                           RegsToCtl_port_contents1_28_port, ZN => n6402);
   U4107 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_28_port, B 
                           => IF_CPathxpc_reg_signal_28_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn129);
   U4108 : AOI21_X1 port map( B1 => n6262, B2 => n3058, A => n3056, ZN => n4306
                           );
   U4109 : AND2_X1 port map( A1 => n3113, A2 => n4306, ZN => n3057);
   U4110 : AOI21_X1 port map( B1 => IF_CPathxN893, B2 => n3111, A => n3057, ZN 
                           => n4087);
   U4111 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_27_port, ZN => n3756);
   U4112 : OAI21_X1 port map( B1 => n4087, B2 => n3100, A => n3756, ZN => n6510
                           );
   U4113 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_27_port, ZN => n6401);
   U4114 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_27_port, B 
                           => IF_CPathxpc_reg_signal_27_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn128);
   U4115 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_26_port, B2 => n3060
                           , A => n3058, ZN => n4305);
   U4116 : NOR2_X1 port map( A1 => n3115, A2 => n4305, ZN => n3059);
   U4117 : AOI21_X1 port map( B1 => IF_CPathxN892, B2 => n3111, A => n3059, ZN 
                           => n4088);
   U4118 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_26_port, ZN => n3779);
   U4119 : OAI21_X1 port map( B1 => n4088, B2 => n3100, A => n3779, ZN => n6511
                           );
   U4120 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_26_port, ZN => n6400);
   U4121 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_26_port, B 
                           => IF_CPathxpc_reg_signal_26_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn127);
   U4122 : AOI21_X1 port map( B1 => n6255, B2 => n3062, A => n3060, ZN => n4373
                           );
   U4123 : AND2_X1 port map( A1 => n3113, A2 => n4373, ZN => n3061);
   U4124 : AOI21_X1 port map( B1 => IF_CPathxN891, B2 => n3115, A => n3061, ZN 
                           => n4089);
   U4125 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_25_port, ZN => n3316);
   U4126 : OAI21_X1 port map( B1 => n4089, B2 => n3100, A => n3316, ZN => n6512
                           );
   U4127 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_25_port, ZN => n6399);
   U4128 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_25_port, B 
                           => IF_CPathxpc_reg_signal_25_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn126);
   U4129 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_24_port, B2 => n3064
                           , A => n3062, ZN => n4291);
   U4130 : NOR2_X1 port map( A1 => n3115, A2 => n4291, ZN => n3063);
   U4131 : AOI21_X1 port map( B1 => IF_CPathxN890, B2 => n3111, A => n3063, ZN 
                           => n4090);
   U4132 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_24_port, ZN => n3873);
   U4133 : OAI21_X1 port map( B1 => n4090, B2 => n3100, A => n3873, ZN => n6513
                           );
   U4134 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_24_port, ZN => n6398);
   U4135 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_24_port, B 
                           => IF_CPathxpc_reg_signal_24_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn125);
   U4136 : AOI21_X1 port map( B1 => n6254, B2 => n3066, A => n3064, ZN => n4320
                           );
   U4137 : AND2_X1 port map( A1 => n3113, A2 => n4320, ZN => n3065);
   U4138 : AOI21_X1 port map( B1 => IF_CPathxN889, B2 => n3111, A => n3065, ZN 
                           => n4091);
   U4139 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_23_port, ZN => n3662);
   U4140 : OAI21_X1 port map( B1 => n4091, B2 => n3100, A => n3662, ZN => n6514
                           );
   U4141 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_23_port, ZN => n6397);
   U4142 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_23_port, B 
                           => IF_CPathxpc_reg_signal_23_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn124);
   U4143 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_22_port, B2 => n3068
                           , A => n3066, ZN => n4316);
   U4144 : NOR2_X1 port map( A1 => n3115, A2 => n4316, ZN => n3067);
   U4145 : AOI21_X1 port map( B1 => IF_CPathxN888, B2 => n3115, A => n3067, ZN 
                           => n4092);
   U4146 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_22_port, ZN => n3684);
   U4147 : OAI21_X1 port map( B1 => n4092, B2 => n3100, A => n3684, ZN => n6515
                           );
   U4148 : AND2_X1 port map( A1 => n4545, A2 => 
                           RegsToCtl_port_contents1_22_port, ZN => n6396);
   U4149 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_22_port, B 
                           => IF_CPathxpc_reg_signal_22_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn123);
   U4150 : AOI21_X1 port map( B1 => n6253, B2 => n3070, A => n3068, ZN => n4342
                           );
   U4151 : AND2_X1 port map( A1 => n3113, A2 => n4342, ZN => n3069);
   U4152 : AOI21_X1 port map( B1 => IF_CPathxN887, B2 => n3111, A => n3069, ZN 
                           => n4093);
   U4153 : CLKBUF_X1 port map( A => n3100, Z => n4282);
   U4154 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_21_port, ZN => n3526);
   U4155 : OAI21_X1 port map( B1 => n4093, B2 => n4282, A => n3526, ZN => n6516
                           );
   U4156 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_21_port, ZN => n6395);
   U4157 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_21_port, B 
                           => IF_CPathxpc_reg_signal_21_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn122);
   U4158 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_20_port, B2 => n3072
                           , A => n3070, ZN => n4312);
   U4159 : NOR2_X1 port map( A1 => n3115, A2 => n4312, ZN => n3071);
   U4160 : AOI21_X1 port map( B1 => IF_CPathxN886, B2 => n3115, A => n3071, ZN 
                           => n4094);
   U4161 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_20_port, ZN => n3705);
   U4162 : OAI21_X1 port map( B1 => n4094, B2 => n4282, A => n3705, ZN => n6517
                           );
   U4163 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_20_port, ZN => n6394);
   U4164 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_20_port, B 
                           => IF_CPathxpc_reg_signal_20_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn121);
   U4165 : AOI21_X1 port map( B1 => n6252, B2 => n3074, A => n3072, ZN => n4338
                           );
   U4166 : AND2_X1 port map( A1 => n3113, A2 => n4338, ZN => n3073);
   U4167 : AOI21_X1 port map( B1 => IF_CPathxN885, B2 => n3115, A => n3073, ZN 
                           => n4095);
   U4168 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_19_port, ZN => n3545);
   U4169 : OAI21_X1 port map( B1 => n4095, B2 => n4282, A => n3545, ZN => n6518
                           );
   U4170 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_19_port, ZN => n6393);
   U4171 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_19_port, B 
                           => IF_CPathxpc_reg_signal_19_port, S => n3093, Z => 
                           DP_OP_1703J95_125_7309xn120);
   U4172 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_18_port, B2 => n3076
                           , A => n3074, ZN => n4346);
   U4173 : NOR2_X1 port map( A1 => n3115, A2 => n4346, ZN => n3075);
   U4174 : AOI21_X1 port map( B1 => IF_CPathxN884, B2 => n3115, A => n3075, ZN 
                           => n4096);
   U4175 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_18_port, ZN => n3507);
   U4176 : OAI21_X1 port map( B1 => n4096, B2 => n3100, A => n3507, ZN => n6519
                           );
   U4177 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_18_port, ZN => n6392);
   U4178 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_18_port, B 
                           => IF_CPathxpc_reg_signal_18_port, S => n3093, Z => 
                           DP_OP_1703J95_125_7309xn119);
   U4179 : AOI21_X1 port map( B1 => n6251, B2 => n3078, A => n3076, ZN => n4335
                           );
   U4180 : AND2_X1 port map( A1 => n3113, A2 => n4335, ZN => n3077);
   U4181 : AOI21_X1 port map( B1 => IF_CPathxN883, B2 => n3115, A => n3077, ZN 
                           => n4097);
   U4182 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_17_port, ZN => n3566);
   U4183 : OAI21_X1 port map( B1 => n4097, B2 => n3100, A => n3566, ZN => n6520
                           );
   U4184 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_17_port, ZN => n6391);
   U4185 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_17_port, B 
                           => IF_CPathxpc_reg_signal_17_port, S => n3093, Z => 
                           DP_OP_1703J95_125_7309xn118);
   U4186 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_16_port, B2 => n3080
                           , A => n3078, ZN => n4285);
   U4187 : NOR2_X1 port map( A1 => n3111, A2 => n4285, ZN => n3079);
   U4188 : AOI21_X1 port map( B1 => IF_CPathxN882, B2 => n3115, A => n3079, ZN 
                           => n4098);
   U4189 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_16_port, ZN => n3901);
   U4190 : OAI21_X1 port map( B1 => n4098, B2 => n3100, A => n3901, ZN => n6521
                           );
   U4191 : AND2_X1 port map( A1 => n4545, A2 => 
                           RegsToCtl_port_contents1_16_port, ZN => n6390);
   U4192 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_16_port, B 
                           => IF_CPathxpc_reg_signal_16_port, S => n3093, Z => 
                           DP_OP_1703J95_125_7309xn117);
   U4193 : AOI21_X1 port map( B1 => n6250, B2 => n3082, A => n3080, ZN => n4332
                           );
   U4194 : AND2_X1 port map( A1 => n3113, A2 => n4332, ZN => n3081);
   U4195 : AOI21_X1 port map( B1 => IF_CPathxN881, B2 => n3115, A => n3081, ZN 
                           => n4099);
   U4196 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_15_port, ZN => n3584);
   U4197 : OAI21_X1 port map( B1 => n4099, B2 => n3100, A => n3584, ZN => n6522
                           );
   U4198 : AND2_X1 port map( A1 => n4546, A2 => 
                           RegsToCtl_port_contents1_15_port, ZN => n6389);
   U4199 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_15_port, B 
                           => IF_CPathxpc_reg_signal_15_port, S => n3093, Z => 
                           DP_OP_1703J95_125_7309xn116);
   U4200 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_14_port, B2 => n3084
                           , A => n3082, ZN => n4353);
   U4201 : NOR2_X1 port map( A1 => n3115, A2 => n4353, ZN => n3083);
   U4202 : AOI21_X1 port map( B1 => IF_CPathxN880, B2 => n3115, A => n3083, ZN 
                           => n4100);
   U4203 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_14_port, ZN => n3455);
   U4204 : OAI21_X1 port map( B1 => n4100, B2 => n3100, A => n3455, ZN => n6523
                           );
   U4205 : AND2_X1 port map( A1 => n4545, A2 => 
                           RegsToCtl_port_contents1_14_port, ZN => n6388);
   U4206 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_14_port, B 
                           => IF_CPathxpc_reg_signal_14_port, S => n3093, Z => 
                           DP_OP_1703J95_125_7309xn115);
   U4207 : AOI21_X1 port map( B1 => n6249, B2 => n3086, A => n3084, ZN => n4329
                           );
   U4208 : AND2_X1 port map( A1 => n3113, A2 => n4329, ZN => n3085);
   U4209 : AOI21_X1 port map( B1 => IF_CPathxN879, B2 => n3115, A => n3085, ZN 
                           => n4101);
   U4210 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_13_port, ZN => n3602);
   U4211 : OAI21_X1 port map( B1 => n4101, B2 => n3100, A => n3602, ZN => n6524
                           );
   U4212 : AND2_X1 port map( A1 => n4545, A2 => 
                           RegsToCtl_port_contents1_13_port, ZN => n6387);
   U4213 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_13_port, B 
                           => IF_CPathxpc_reg_signal_13_port, S => n3093, Z => 
                           DP_OP_1703J95_125_7309xn114);
   U4214 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_12_port, B2 => n3088
                           , A => n3086, ZN => n4311);
   U4215 : NOR2_X1 port map( A1 => n3115, A2 => n4311, ZN => n3087);
   U4216 : AOI21_X1 port map( B1 => IF_CPathxN878, B2 => n3115, A => n3087, ZN 
                           => n4102);
   U4217 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_12_port, ZN => n3733);
   U4218 : OAI21_X1 port map( B1 => n4102, B2 => n3100, A => n3733, ZN => n6525
                           );
   U4219 : AND2_X1 port map( A1 => n4545, A2 => 
                           RegsToCtl_port_contents1_12_port, ZN => n6386);
   U4220 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_12_port, B 
                           => IF_CPathxpc_reg_signal_12_port, S => n3093, Z => 
                           DP_OP_1703J95_125_7309xn113);
   U4221 : AOI21_X1 port map( B1 => n6248, B2 => n3091, A => n3088, ZN => n4326
                           );
   U4222 : AND2_X1 port map( A1 => n3113, A2 => n4326, ZN => n3089);
   U4223 : AOI21_X1 port map( B1 => IF_CPathxN877, B2 => n3111, A => n3089, ZN 
                           => n4103);
   U4224 : NAND2_X1 port map( A1 => n3090, A2 => 
                           IF_CPathxpc_next_signal_11_port, ZN => n3622);
   U4225 : OAI21_X1 port map( B1 => n4103, B2 => n3100, A => n3622, ZN => n6526
                           );
   U4226 : AND2_X1 port map( A1 => n4545, A2 => 
                           RegsToCtl_port_contents1_11_port, ZN => n6385);
   U4227 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_11_port, B 
                           => IF_CPathxpc_reg_signal_11_port, S => n3093, Z => 
                           DP_OP_1703J95_125_7309xn112);
   U4228 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_10_port, B2 => n3094
                           , A => n3091, ZN => n4299);
   U4229 : NOR2_X1 port map( A1 => n3115, A2 => n4299, ZN => n3092);
   U4230 : AOI21_X1 port map( B1 => IF_CPathxN876, B2 => n3111, A => n3092, ZN 
                           => n4104);
   U4231 : NAND2_X1 port map( A1 => n4181, A2 => 
                           IF_CPathxpc_next_signal_10_port, ZN => n3802);
   U4232 : OAI21_X1 port map( B1 => n4104, B2 => n3100, A => n3802, ZN => n6527
                           );
   U4233 : AND2_X1 port map( A1 => n4545, A2 => 
                           RegsToCtl_port_contents1_10_port, ZN => n6384);
   U4234 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_10_port, B 
                           => IF_CPathxpc_reg_signal_10_port, S => n3093, Z => 
                           DP_OP_1703J95_125_7309xn111);
   U4235 : AOI21_X1 port map( B1 => n6247, B2 => n3096, A => n3094, ZN => n4376
                           );
   U4236 : AND2_X1 port map( A1 => n3113, A2 => n4376, ZN => n3095);
   U4237 : AOI21_X1 port map( B1 => IF_CPathxN875, B2 => n3111, A => n3095, ZN 
                           => n4105);
   U4238 : NAND2_X1 port map( A1 => n4181, A2 => IF_CPathxpc_next_signal_9_port
                           , ZN => n3302);
   U4239 : OAI21_X1 port map( B1 => n4105, B2 => n3100, A => n3302, ZN => n6528
                           );
   U4240 : AND2_X1 port map( A1 => n4545, A2 => RegsToCtl_port_contents1_9_port
                           , ZN => n6383);
   U4241 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_9_port, B 
                           => IF_CPathxpc_reg_signal_9_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn110);
   U4242 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_8_port, B2 => n3098,
                           A => n3096, ZN => n4325);
   U4243 : NOR2_X1 port map( A1 => n3115, A2 => n4325, ZN => n3097);
   U4244 : AOI21_X1 port map( B1 => IF_CPathxN874, B2 => n3111, A => n3097, ZN 
                           => n4106);
   U4245 : NAND2_X1 port map( A1 => n4181, A2 => IF_CPathxpc_next_signal_8_port
                           , ZN => n3643);
   U4246 : OAI21_X1 port map( B1 => n4106, B2 => n3100, A => n3643, ZN => n6529
                           );
   U4247 : AND2_X1 port map( A1 => n4545, A2 => RegsToCtl_port_contents1_8_port
                           , ZN => n6382);
   U4248 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_8_port, B 
                           => IF_CPathxpc_reg_signal_8_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn109);
   U4249 : AOI21_X1 port map( B1 => n6244, B2 => n3101, A => n3098, ZN => n4368
                           );
   U4250 : AND2_X1 port map( A1 => n3113, A2 => n4368, ZN => n3099);
   U4251 : AOI21_X1 port map( B1 => IF_CPathxN873, B2 => n3111, A => n3099, ZN 
                           => n4107);
   U4252 : NAND2_X1 port map( A1 => n4181, A2 => IF_CPathxpc_next_signal_7_port
                           , ZN => n3335);
   U4253 : OAI21_X1 port map( B1 => n4107, B2 => n3100, A => n3335, ZN => n6530
                           );
   U4254 : AND2_X1 port map( A1 => n4545, A2 => RegsToCtl_port_contents1_7_port
                           , ZN => n6381);
   U4255 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_7_port, B 
                           => IF_CPathxpc_reg_signal_7_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn108);
   U4256 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_6_port, B2 => n3103,
                           A => n3101, ZN => n4379);
   U4257 : NOR2_X1 port map( A1 => n3115, A2 => n4379, ZN => n3102);
   U4258 : AOI21_X1 port map( B1 => IF_CPathxN872, B2 => n3111, A => n3102, ZN 
                           => n4108);
   U4259 : NAND2_X1 port map( A1 => n4181, A2 => IF_CPathxpc_next_signal_6_port
                           , ZN => n3283);
   U4260 : OAI21_X1 port map( B1 => n4108, B2 => n4282, A => n3283, ZN => n6531
                           );
   U4261 : AND2_X1 port map( A1 => n4545, A2 => RegsToCtl_port_contents1_6_port
                           , ZN => n6380);
   U4262 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_6_port, B 
                           => IF_CPathxpc_reg_signal_6_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn107);
   U4263 : AOI21_X1 port map( B1 => n6243, B2 => n3105, A => n3103, ZN => n4365
                           );
   U4264 : AND2_X1 port map( A1 => n3113, A2 => n4365, ZN => n3104);
   U4265 : AOI21_X1 port map( B1 => IF_CPathxN871, B2 => n3111, A => n3104, ZN 
                           => n4109);
   U4266 : NAND2_X1 port map( A1 => n4181, A2 => IF_CPathxpc_next_signal_5_port
                           , ZN => n3365);
   U4267 : OAI21_X1 port map( B1 => n4109, B2 => n4282, A => n3365, ZN => n6532
                           );
   U4268 : AND2_X1 port map( A1 => n4545, A2 => RegsToCtl_port_contents1_5_port
                           , ZN => n6379);
   U4269 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_5_port, B 
                           => IF_CPathxpc_reg_signal_5_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn106);
   U4270 : OAI21_X1 port map( B1 => IF_CPathxpc_reg_signal_4_port, B2 => n3108,
                           A => n3105, ZN => n4352);
   U4271 : NOR2_X1 port map( A1 => n3111, A2 => n4352, ZN => n3106);
   U4272 : AOI21_X1 port map( B1 => IF_CPathxN870, B2 => n3111, A => n3106, ZN 
                           => n4110);
   U4273 : NAND2_X1 port map( A1 => n4181, A2 => IF_CPathxpc_next_signal_4_port
                           , ZN => n3473);
   U4274 : OAI21_X1 port map( B1 => n4110, B2 => n4282, A => n3473, ZN => n6533
                           );
   U4275 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_4_port, B 
                           => IF_CPathxpc_reg_signal_4_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn105);
   U4276 : NOR2_X1 port map( A1 => n3115, A2 => IF_CPathxpc_reg_signal_2_port, 
                           ZN => n3107);
   U4277 : AOI21_X1 port map( B1 => IF_CPathxN868, B2 => n3111, A => n3107, ZN 
                           => n4112);
   U4278 : NAND2_X1 port map( A1 => n4181, A2 => IF_CPathxpc_next_signal_2_port
                           , ZN => n3432);
   U4279 : OAI21_X1 port map( B1 => n4112, B2 => n4282, A => n3432, ZN => n6535
                           );
   U4280 : AOI21_X1 port map( B1 => n6245, B2 => n6204, A => n3108, ZN => n4359
                           );
   U4281 : AND2_X1 port map( A1 => n3113, A2 => n4359, ZN => n3109);
   U4282 : AOI21_X1 port map( B1 => IF_CPathxN869, B2 => n3111, A => n3109, ZN 
                           => n4111);
   U4283 : NAND2_X1 port map( A1 => n4181, A2 => IF_CPathxpc_next_signal_3_port
                           , ZN => n3411);
   U4284 : OAI21_X1 port map( B1 => n4111, B2 => n4282, A => n3411, ZN => n6534
                           );
   U4285 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_3_port, B 
                           => IF_CPathxpc_reg_signal_3_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn104);
   U4286 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_2_port, B 
                           => IF_CPathxpc_reg_signal_2_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn103);
   U4287 : AND2_X1 port map( A1 => n3113, A2 => IF_CPathxpc_reg_signal_1_port, 
                           ZN => n3110);
   U4288 : AOI21_X1 port map( B1 => IF_CPathxN867, B2 => n3111, A => n3110, ZN 
                           => n4113);
   U4289 : NAND2_X1 port map( A1 => n4181, A2 => IF_CPathxpc_next_signal_1_port
                           , ZN => n3389);
   U4290 : OAI21_X1 port map( B1 => n4113, B2 => n4282, A => n3389, ZN => n6536
                           );
   U4291 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_1_port, B 
                           => IF_CPathxpc_reg_signal_1_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn102);
   U4292 : MUX2_X1 port map( A => 
                           IF_CPathxRegsToCtl_data_signal_contents1_0_port, B 
                           => IF_CPathxpc_reg_signal_0_port, S => n3112, Z => 
                           DP_OP_1703J95_125_7309xn101);
   U4293 : AND2_X1 port map( A1 => n4545, A2 => DecToCtl_port_imm_31_port, ZN 
                           => n6422);
   U4294 : AND2_X1 port map( A1 => n4545, A2 => DecToCtl_port_imm_30_port, ZN 
                           => n6421);
   U4295 : AND2_X1 port map( A1 => n4545, A2 => DecToCtl_port_imm_29_port, ZN 
                           => n6420);
   U4296 : NOR2_X1 port map( A1 => rst, A2 => n6223, ZN => IF_CPathxN2186);
   U4297 : AND2_X1 port map( A1 => n4545, A2 => DecToCtl_port_imm_27_port, ZN 
                           => n6419);
   U4298 : AND2_X1 port map( A1 => n4545, A2 => DecToCtl_port_imm_26_port, ZN 
                           => n6418);
   U4299 : NOR2_X1 port map( A1 => rst, A2 => n6214, ZN => IF_CPathxN2183);
   U4300 : NOR2_X1 port map( A1 => rst, A2 => n6216, ZN => IF_CPathxN2182);
   U4301 : NOR2_X1 port map( A1 => rst, A2 => n6215, ZN => IF_CPathxN2181);
   U4302 : AND2_X1 port map( A1 => n4545, A2 => DecToCtl_port_imm_22_port, ZN 
                           => n6417);
   U4303 : AND2_X1 port map( A1 => n6180, A2 => DecToCtl_port_imm_21_port, ZN 
                           => n6416);
   U4304 : CLKBUF_X1 port map( A => n4671, Z => n4667);
   U4305 : AND2_X1 port map( A1 => n4667, A2 => DecToCtl_port_imm_20_port, ZN 
                           => n6415);
   U4306 : AND2_X1 port map( A1 => n4671, A2 => DecToCtl_port_imm_19_port, ZN 
                           => n6414);
   U4307 : NOR2_X1 port map( A1 => rst, A2 => n6222, ZN => IF_CPathxN2176);
   U4308 : AND2_X1 port map( A1 => n4671, A2 => DecToCtl_port_imm_17_port, ZN 
                           => n6413);
   U4309 : NOR2_X1 port map( A1 => rst, A2 => n6221, ZN => IF_CPathxN2174);
   U4310 : AND2_X1 port map( A1 => n4545, A2 => DecToCtl_port_imm_15_port, ZN 
                           => n6412);
   U4311 : AND2_X1 port map( A1 => n4547, A2 => DecToCtl_port_imm_14_port, ZN 
                           => n6411);
   U4312 : AND2_X1 port map( A1 => n6180, A2 => DecToCtl_port_imm_13_port, ZN 
                           => n6410);
   U4313 : AND2_X1 port map( A1 => n4546, A2 => DecToCtl_port_imm_12_port, ZN 
                           => n6409);
   U4314 : AND2_X1 port map( A1 => n4667, A2 => DecToCtl_port_imm_11_port, ZN 
                           => n6408);
   U4315 : NOR2_X1 port map( A1 => rst, A2 => n6220, ZN => IF_CPathxN2168);
   U4316 : NOR2_X1 port map( A1 => rst, A2 => n6217, ZN => IF_CPathxN2167);
   U4317 : AND2_X1 port map( A1 => n4545, A2 => DecToCtl_port_imm_8_port, ZN =>
                           n6407);
   U4318 : NOR2_X1 port map( A1 => rst, A2 => n6219, ZN => IF_CPathxN2165);
   U4319 : AND2_X1 port map( A1 => n4571, A2 => DecToCtl_port_imm_6_port, ZN =>
                           n6406);
   U4320 : NOR2_X1 port map( A1 => rst, A2 => n6218, ZN => IF_CPathxN2163);
   U4321 : AND2_X1 port map( A1 => n3113, A2 => IF_CPathxpc_reg_signal_0_port, 
                           ZN => n3114);
   U4322 : AOI21_X1 port map( B1 => IF_CPathxN866, B2 => n3115, A => n3114, ZN 
                           => n4114);
   U4323 : NAND2_X1 port map( A1 => n4181, A2 => IF_CPathxpc_next_signal_0_port
                           , ZN => n3923);
   U4324 : OAI21_X1 port map( B1 => n4114, B2 => n4282, A => n3923, ZN => n6537
                           );
   U4325 : INV_X2 port map( A => n6227, ZN => n4275);
   U4326 : NAND2_X1 port map( A1 => IF_CPathxsection_0_port, A2 => n4275, ZN =>
                           n4188);
   U4327 : NAND2_X1 port map( A1 => n6196, A2 => n6228, ZN => n6182);
   U4328 : NOR2_X1 port map( A1 => n4188, A2 => n6182, ZN => n4541);
   U4329 : NAND2_X1 port map( A1 => n6197, A2 => DecToCtl_port_encType_2_port, 
                           ZN => n4225);
   U4330 : INV_X1 port map( A => n4225, ZN => n4533);
   U4331 : NAND2_X1 port map( A1 => DecToCtl_port_encType_1_port, A2 => n4533, 
                           ZN => n4454);
   U4332 : NAND3_X1 port map( A1 => DecToCtl_port_instrType_2_port, A2 => n6226
                           , A3 => n6189, ZN => n4460);
   U4333 : NOR2_X1 port map( A1 => DecToCtl_port_instrType_4_port, A2 => n4460,
                           ZN => n4527);
   U4334 : NAND2_X1 port map( A1 => DecToCtl_port_instrType_0_port, A2 => 
                           DecToCtl_port_instrType_1_port, ZN => n4266);
   U4335 : INV_X1 port map( A => n4266, ZN => n4409);
   U4336 : NAND2_X1 port map( A1 => n4527, A2 => n4409, ZN => n4437);
   U4337 : NOR2_X1 port map( A1 => n4454, A2 => n4437, ZN => n4434);
   U4338 : NAND2_X1 port map( A1 => n4541, A2 => n4434, ZN => n4430);
   U4339 : NOR2_X1 port map( A1 => DecToCtl_port_instrType_5_port, A2 => n6189,
                           ZN => n4244);
   U4340 : NOR2_X1 port map( A1 => n2953, A2 => DecToCtl_port_instrType_0_port,
                           ZN => n4532);
   U4341 : INV_X1 port map( A => n4532, ZN => n4184);
   U4342 : NAND3_X1 port map( A1 => DecToCtl_port_encType_0_port, A2 => 
                           DecToCtl_port_encType_1_port, A3 => n6230, ZN => 
                           n4517);
   U4343 : NOR2_X1 port map( A1 => n4184, A2 => n4517, ZN => n4408);
   U4344 : NOR2_X1 port map( A1 => DecToCtl_port_instrType_4_port, A2 => n6195,
                           ZN => n4242);
   U4345 : NAND3_X1 port map( A1 => n4244, A2 => n4408, A3 => n4242, ZN => 
                           n4443);
   U4346 : NAND2_X1 port map( A1 => n6232, A2 => n2953, ZN => n4241);
   U4347 : INV_X1 port map( A => n4241, ZN => n4528);
   U4348 : NAND2_X1 port map( A1 => DecToCtl_port_instrType_4_port, A2 => n4528
                           , ZN => n4182);
   U4349 : NOR3_X1 port map( A1 => DecToCtl_port_instrType_3_port, A2 => n6195,
                           A3 => n4182, ZN => n4262);
   U4350 : NAND2_X1 port map( A1 => n4262, A2 => n6226, ZN => n4438);
   U4351 : NOR2_X1 port map( A1 => n4454, A2 => n4438, ZN => n4435);
   U4352 : INV_X1 port map( A => n4435, ZN => n4432);
   U4353 : INV_X1 port map( A => n4541, ZN => n4521);
   U4354 : AOI21_X1 port map( B1 => n4443, B2 => n4432, A => n4521, ZN => n4429
                           );
   U4355 : AOI21_X1 port map( B1 => 
                           IF_CPathxCtlToALU_data_signal_alu_fun_1_port, B2 => 
                           n4430, A => n4429, ZN => n3116);
   U4356 : INV_X1 port map( A => n3116, ZN => IF_CPathxN1629);
   U4357 : AOI21_X1 port map( B1 => 
                           IF_CPathxCtlToALU_data_signal_op2_sel_0_port, B2 => 
                           n4430, A => n4429, ZN => n3117);
   U4358 : INV_X1 port map( A => n3117, ZN => IF_CPathxN1667);
   U4359 : AND2_X1 port map( A1 => n4547, A2 => IF_CPathxpc_reg_signal_0_port, 
                           ZN => IF_CPathxN1936);
   U4360 : CLKBUF_X1 port map( A => n3207, Z => n3257);
   U4361 : CLKBUF_X1 port map( A => n3242, Z => n3256);
   U4362 : AOI222_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_0_port, 
                           B1 => n3256, B2 => 
                           CtlToALU_port_reg1_contents_0_port, C1 => n3258, C2 
                           => CtlToALU_port_imm_0_port, ZN => n3118);
   U4363 : INV_X1 port map( A => n3118, ZN => IF_ALUxN112);
   U4364 : INV_X1 port map( A => n6227, ZN => n4277);
   U4365 : NAND2_X1 port map( A1 => n4571, A2 => n6227, ZN => n4268);
   U4366 : INV_X1 port map( A => n4268, ZN => n4210);
   U4367 : AOI22_X1 port map( A1 => n6422, A2 => n4277, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_31_port, ZN => 
                           n3119);
   U4368 : INV_X1 port map( A => n3119, ZN => n6643);
   U4369 : INV_X1 port map( A => n6405, ZN => n3120);
   U4370 : NAND2_X1 port map( A1 => n4275, A2 => n4671, ZN => n3235);
   U4371 : CLKBUF_X2 port map( A => n3235, Z => n4276);
   U4372 : OAI22_X1 port map( A1 => n3120, A2 => n6207, B1 => n4276, B2 => 
                           n6346, ZN => n6642);
   U4373 : AND2_X1 port map( A1 => n4671, A2 => IF_CPathxpc_reg_signal_31_port,
                           ZN => IF_CPathxN1967);
   U4374 : AOI22_X1 port map( A1 => n6419, A2 => n4277, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_27_port, ZN => 
                           n3121);
   U4375 : INV_X1 port map( A => n3121, ZN => n6647);
   U4376 : NOR2_X1 port map( A1 => rst, A2 => n6262, ZN => IF_CPathxN1963);
   U4377 : INV_X1 port map( A => n6401, ZN => n3122);
   U4378 : OAI22_X1 port map( A1 => n3122, A2 => n6207, B1 => n4276, B2 => 
                           n6347, ZN => n6626);
   U4379 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_27_port, 
                           ZN => n3125);
   U4380 : NAND2_X1 port map( A1 => n3256, A2 => 
                           CtlToALU_port_reg1_contents_27_port, ZN => n3124);
   U4381 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_27_port, ZN 
                           => n3123);
   U4382 : NAND3_X1 port map( A1 => n3125, A2 => n3124, A3 => n3123, ZN => 
                           IF_ALUxN139);
   U4383 : AOI22_X1 port map( A1 => n6418, A2 => n4277, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_26_port, ZN => 
                           n3126);
   U4384 : INV_X1 port map( A => n3126, ZN => n6648);
   U4385 : AND2_X1 port map( A1 => n4545, A2 => IF_CPathxpc_reg_signal_26_port,
                           ZN => IF_CPathxN1962);
   U4386 : INV_X1 port map( A => n6400, ZN => n3127);
   U4387 : OAI22_X1 port map( A1 => n3127, A2 => n6207, B1 => n4276, B2 => 
                           n6348, ZN => n6628);
   U4388 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_26_port, 
                           ZN => n3130);
   U4389 : NAND2_X1 port map( A1 => n3256, A2 => 
                           CtlToALU_port_reg1_contents_26_port, ZN => n3129);
   U4390 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_26_port, ZN 
                           => n3128);
   U4391 : NAND3_X1 port map( A1 => n3130, A2 => n3129, A3 => n3128, ZN => 
                           IF_ALUxN138);
   U4392 : OAI22_X1 port map( A1 => n4268, A2 => n6330, B1 => n4276, B2 => 
                           n6214, ZN => n6649);
   U4393 : NOR2_X1 port map( A1 => rst, A2 => n6255, ZN => IF_CPathxN1961);
   U4394 : INV_X1 port map( A => n6399, ZN => n3131);
   U4395 : OAI22_X1 port map( A1 => n3131, A2 => n4275, B1 => n4276, B2 => 
                           n6349, ZN => n6586);
   U4396 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_25_port, 
                           ZN => n3134);
   U4397 : NAND2_X1 port map( A1 => n3256, A2 => 
                           CtlToALU_port_reg1_contents_25_port, ZN => n3133);
   U4398 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_25_port, ZN 
                           => n3132);
   U4399 : NAND3_X1 port map( A1 => n3134, A2 => n3133, A3 => n3132, ZN => 
                           IF_ALUxN137);
   U4400 : OAI22_X1 port map( A1 => n4268, A2 => n6331, B1 => n4276, B2 => 
                           n6215, ZN => n6651);
   U4401 : NOR2_X1 port map( A1 => rst, A2 => n6254, ZN => IF_CPathxN1959);
   U4402 : INV_X1 port map( A => n6397, ZN => n3135);
   U4403 : OAI22_X1 port map( A1 => n3135, A2 => n4277, B1 => n4276, B2 => 
                           n6350, ZN => n6618);
   U4404 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_23_port, 
                           ZN => n3138);
   U4405 : NAND2_X1 port map( A1 => n3256, A2 => 
                           CtlToALU_port_reg1_contents_23_port, ZN => n3137);
   U4406 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_23_port, ZN 
                           => n3136);
   U4407 : NAND3_X1 port map( A1 => n3138, A2 => n3137, A3 => n3136, ZN => 
                           IF_ALUxN135);
   U4408 : AOI22_X1 port map( A1 => n6417, A2 => n4277, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_22_port, ZN => 
                           n3139);
   U4409 : INV_X1 port map( A => n3139, ZN => n6652);
   U4410 : AND2_X1 port map( A1 => n4547, A2 => IF_CPathxpc_reg_signal_22_port,
                           ZN => IF_CPathxN1958);
   U4411 : INV_X1 port map( A => n6396, ZN => n3140);
   U4412 : OAI22_X1 port map( A1 => n3140, A2 => n6207, B1 => n4276, B2 => 
                           n6351, ZN => n6620);
   U4413 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_22_port, 
                           ZN => n3143);
   U4414 : NAND2_X1 port map( A1 => n3256, A2 => 
                           CtlToALU_port_reg1_contents_22_port, ZN => n3142);
   U4415 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_22_port, ZN 
                           => n3141);
   U4416 : NAND3_X1 port map( A1 => n3143, A2 => n3142, A3 => n3141, ZN => 
                           IF_ALUxN134);
   U4417 : AOI22_X1 port map( A1 => n6416, A2 => n4277, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_21_port, ZN => 
                           n3144);
   U4418 : INV_X1 port map( A => n3144, ZN => n6653);
   U4419 : NOR2_X1 port map( A1 => rst, A2 => n6253, ZN => IF_CPathxN1957);
   U4420 : INV_X1 port map( A => n6395, ZN => n3145);
   U4421 : OAI22_X1 port map( A1 => n3145, A2 => n6207, B1 => n4276, B2 => 
                           n6352, ZN => n6604);
   U4422 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_21_port, 
                           ZN => n3148);
   U4423 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_21_port, ZN => n3147);
   U4424 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_21_port, ZN 
                           => n3146);
   U4425 : NAND3_X1 port map( A1 => n3148, A2 => n3147, A3 => n3146, ZN => 
                           IF_ALUxN133);
   U4426 : OAI22_X1 port map( A1 => n4268, A2 => n6332, B1 => n4276, B2 => 
                           n6216, ZN => n6650);
   U4427 : AND2_X1 port map( A1 => n6180, A2 => IF_CPathxpc_reg_signal_24_port,
                           ZN => IF_CPathxN1960);
   U4428 : INV_X1 port map( A => n6398, ZN => n3149);
   U4429 : OAI22_X1 port map( A1 => n3149, A2 => n6207, B1 => n4276, B2 => 
                           n6353, ZN => n6636);
   U4430 : AOI22_X1 port map( A1 => n6412, A2 => n4277, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_15_port, ZN => 
                           n3150);
   U4431 : INV_X1 port map( A => n3150, ZN => n6659);
   U4432 : NOR2_X1 port map( A1 => rst, A2 => n6250, ZN => IF_CPathxN1951);
   U4433 : INV_X1 port map( A => n6389, ZN => n3151);
   U4434 : OAI22_X1 port map( A1 => n3151, A2 => n4275, B1 => n4276, B2 => 
                           n6354, ZN => n6610);
   U4435 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_15_port, 
                           ZN => n3154);
   U4436 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_15_port, ZN => n3153);
   U4437 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_15_port, ZN 
                           => n3152);
   U4438 : NAND3_X1 port map( A1 => n3154, A2 => n3153, A3 => n3152, ZN => 
                           IF_ALUxN127);
   U4439 : AOI22_X1 port map( A1 => n6411, A2 => n6207, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_14_port, ZN => 
                           n3155);
   U4440 : INV_X1 port map( A => n3155, ZN => n6660);
   U4441 : AND2_X1 port map( A1 => n4546, A2 => IF_CPathxpc_reg_signal_14_port,
                           ZN => IF_CPathxN1950);
   U4442 : INV_X1 port map( A => n6388, ZN => n3156);
   U4443 : OAI22_X1 port map( A1 => n3156, A2 => n4275, B1 => n3235, B2 => 
                           n6355, ZN => n6598);
   U4444 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_14_port, 
                           ZN => n3159);
   U4445 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_14_port, ZN => n3158);
   U4446 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_14_port, ZN 
                           => n3157);
   U4447 : NAND3_X1 port map( A1 => n3159, A2 => n3158, A3 => n3157, ZN => 
                           IF_ALUxN126);
   U4448 : AOI22_X1 port map( A1 => n6410, A2 => n6207, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_13_port, ZN => 
                           n3160);
   U4449 : INV_X1 port map( A => n3160, ZN => n6661);
   U4450 : NOR2_X1 port map( A1 => rst, A2 => n6249, ZN => IF_CPathxN1949);
   U4451 : INV_X1 port map( A => n6387, ZN => n3161);
   U4452 : OAI22_X1 port map( A1 => n3161, A2 => n6207, B1 => n4276, B2 => 
                           n6356, ZN => n6612);
   U4453 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_13_port, 
                           ZN => n3164);
   U4454 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_13_port, ZN => n3163);
   U4455 : NAND2_X1 port map( A1 => n3208, A2 => CtlToALU_port_imm_13_port, ZN 
                           => n3162);
   U4456 : NAND3_X1 port map( A1 => n3164, A2 => n3163, A3 => n3162, ZN => 
                           IF_ALUxN125);
   U4457 : AOI22_X1 port map( A1 => n6409, A2 => n6207, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_12_port, ZN => 
                           n3165);
   U4458 : INV_X1 port map( A => n3165, ZN => n6662);
   U4459 : AND2_X1 port map( A1 => n4667, A2 => IF_CPathxpc_reg_signal_12_port,
                           ZN => IF_CPathxN1948);
   U4460 : INV_X1 port map( A => n6386, ZN => n3166);
   U4461 : OAI22_X1 port map( A1 => n3166, A2 => n6207, B1 => n4276, B2 => 
                           n6357, ZN => n6624);
   U4462 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_12_port, 
                           ZN => n3169);
   U4463 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_12_port, ZN => n3168);
   U4464 : NAND2_X1 port map( A1 => n3208, A2 => CtlToALU_port_imm_12_port, ZN 
                           => n3167);
   U4465 : NAND3_X1 port map( A1 => n3169, A2 => n3168, A3 => n3167, ZN => 
                           IF_ALUxN124);
   U4466 : AOI22_X1 port map( A1 => n6407, A2 => n6207, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_8_port, ZN => 
                           n3170);
   U4467 : INV_X1 port map( A => n3170, ZN => n6666);
   U4468 : CLKBUF_X1 port map( A => n4671, Z => n6178);
   U4469 : AND2_X1 port map( A1 => n6178, A2 => IF_CPathxpc_reg_signal_8_port, 
                           ZN => IF_CPathxN1944);
   U4470 : INV_X1 port map( A => n6382, ZN => n3171);
   U4471 : OAI22_X1 port map( A1 => n3171, A2 => n6207, B1 => n4276, B2 => 
                           n6358, ZN => n6616);
   U4472 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_8_port, 
                           ZN => n3174);
   U4473 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_8_port, ZN => n3173);
   U4474 : NAND2_X1 port map( A1 => n3208, A2 => CtlToALU_port_imm_8_port, ZN 
                           => n3172);
   U4475 : NAND3_X1 port map( A1 => n3174, A2 => n3173, A3 => n3172, ZN => 
                           IF_ALUxN120);
   U4476 : OAI22_X1 port map( A1 => n4268, A2 => n6333, B1 => n4276, B2 => 
                           n6217, ZN => n6665);
   U4477 : NOR2_X1 port map( A1 => rst, A2 => n6247, ZN => IF_CPathxN1945);
   U4478 : INV_X1 port map( A => n6383, ZN => n3175);
   U4479 : OAI22_X1 port map( A1 => n3175, A2 => n6207, B1 => n4276, B2 => 
                           n6359, ZN => n6584);
   U4480 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_9_port, 
                           ZN => n3178);
   U4481 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_9_port, ZN => n3177);
   U4482 : NAND2_X1 port map( A1 => n3208, A2 => CtlToALU_port_imm_9_port, ZN 
                           => n3176);
   U4483 : NAND3_X1 port map( A1 => n3178, A2 => n3177, A3 => n3176, ZN => 
                           IF_ALUxN121);
   U4484 : NOR2_X1 port map( A1 => rst, A2 => n6204, ZN => IF_CPathxN1939);
   U4485 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_3_port, 
                           ZN => n3181);
   U4486 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_3_port, ZN => n3180);
   U4487 : NAND2_X1 port map( A1 => n3208, A2 => CtlToALU_port_imm_3_port, ZN 
                           => n3179);
   U4488 : NAND3_X1 port map( A1 => n3181, A2 => n3180, A3 => n3179, ZN => 
                           IF_ALUxN115);
   U4489 : AND2_X1 port map( A1 => n4571, A2 => IF_CPathxpc_reg_signal_4_port, 
                           ZN => IF_CPathxN1940);
   U4490 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_4_port, 
                           ZN => n3184);
   U4491 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_4_port, ZN => n3183);
   U4492 : NAND2_X1 port map( A1 => n3208, A2 => CtlToALU_port_imm_4_port, ZN 
                           => n3182);
   U4493 : NAND3_X1 port map( A1 => n3184, A2 => n3183, A3 => n3182, ZN => 
                           IF_ALUxN116);
   U4494 : NOR2_X1 port map( A1 => rst, A2 => n6323, ZN => IF_CPathxN1937);
   U4495 : AOI222_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_1_port, 
                           B1 => n3256, B2 => 
                           CtlToALU_port_reg1_contents_1_port, C1 => n3258, C2 
                           => CtlToALU_port_imm_1_port, ZN => n3407);
   U4496 : INV_X1 port map( A => n3407, ZN => IF_ALUxN113);
   U4497 : NOR2_X1 port map( A1 => rst, A2 => n6245, ZN => IF_CPathxN1938);
   U4498 : NAND2_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_2_port, 
                           ZN => n3187);
   U4499 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_2_port, ZN => n3186);
   U4500 : NAND2_X1 port map( A1 => n3208, A2 => CtlToALU_port_imm_2_port, ZN 
                           => n3185);
   U4501 : NAND3_X1 port map( A1 => n3187, A2 => n3186, A3 => n3185, ZN => 
                           IF_ALUxN114);
   U4502 : OAI22_X1 port map( A1 => n4268, A2 => n6334, B1 => n4276, B2 => 
                           n6218, ZN => n6669);
   U4503 : NOR2_X1 port map( A1 => rst, A2 => n6243, ZN => IF_CPathxN1941);
   U4504 : INV_X1 port map( A => n6379, ZN => n3188);
   U4505 : OAI22_X1 port map( A1 => n3188, A2 => n6207, B1 => n4276, B2 => 
                           n6360, ZN => n6590);
   U4506 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_5_port, 
                           ZN => n3191);
   U4507 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_5_port, ZN => n3190);
   U4508 : NAND2_X1 port map( A1 => n3208, A2 => CtlToALU_port_imm_5_port, ZN 
                           => n3189);
   U4509 : NAND3_X1 port map( A1 => n3191, A2 => n3190, A3 => n3189, ZN => 
                           IF_ALUxN117);
   U4510 : AOI22_X1 port map( A1 => n6406, A2 => n6207, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_6_port, ZN => 
                           n3192);
   U4511 : INV_X1 port map( A => n3192, ZN => n6668);
   U4512 : AND2_X1 port map( A1 => n4546, A2 => IF_CPathxpc_reg_signal_6_port, 
                           ZN => IF_CPathxN1942);
   U4513 : INV_X1 port map( A => n6380, ZN => n3193);
   U4514 : OAI22_X1 port map( A1 => n3193, A2 => n6207, B1 => n3235, B2 => 
                           n6361, ZN => n6582);
   U4515 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_6_port, 
                           ZN => n3196);
   U4516 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_6_port, ZN => n3195);
   U4517 : NAND2_X1 port map( A1 => n3208, A2 => CtlToALU_port_imm_6_port, ZN 
                           => n3194);
   U4518 : NAND3_X1 port map( A1 => n3196, A2 => n3195, A3 => n3194, ZN => 
                           IF_ALUxN118);
   U4519 : OAI22_X1 port map( A1 => n4268, A2 => n6335, B1 => n4276, B2 => 
                           n6219, ZN => n6667);
   U4520 : NOR2_X1 port map( A1 => rst, A2 => n6244, ZN => IF_CPathxN1943);
   U4521 : INV_X1 port map( A => n6381, ZN => n3197);
   U4522 : OAI22_X1 port map( A1 => n3197, A2 => n4277, B1 => n4276, B2 => 
                           n6362, ZN => n6588);
   U4523 : NAND2_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_7_port, 
                           ZN => n3200);
   U4524 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_7_port, ZN => n3199);
   U4525 : NAND2_X1 port map( A1 => n3208, A2 => CtlToALU_port_imm_7_port, ZN 
                           => n3198);
   U4526 : NAND3_X1 port map( A1 => n3200, A2 => n3199, A3 => n3198, ZN => 
                           IF_ALUxN119);
   U4527 : AOI22_X1 port map( A1 => n6408, A2 => n6207, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_11_port, ZN => 
                           n3201);
   U4528 : INV_X1 port map( A => n3201, ZN => n6663);
   U4529 : NOR2_X1 port map( A1 => rst, A2 => n6248, ZN => IF_CPathxN1947);
   U4530 : INV_X1 port map( A => n6385, ZN => n3202);
   U4531 : OAI22_X1 port map( A1 => n3202, A2 => n6207, B1 => n4276, B2 => 
                           n6363, ZN => n6614);
   U4532 : NAND2_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_11_port, 
                           ZN => n3205);
   U4533 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_11_port, ZN => n3204);
   U4534 : NAND2_X1 port map( A1 => n3208, A2 => CtlToALU_port_imm_11_port, ZN 
                           => n3203);
   U4535 : NAND3_X1 port map( A1 => n3205, A2 => n3204, A3 => n3203, ZN => 
                           IF_ALUxN123);
   U4536 : OAI22_X1 port map( A1 => n4268, A2 => n6336, B1 => n4276, B2 => 
                           n6220, ZN => n6664);
   U4537 : AND2_X1 port map( A1 => n6178, A2 => IF_CPathxpc_reg_signal_10_port,
                           ZN => IF_CPathxN1946);
   U4538 : INV_X1 port map( A => n6384, ZN => n3206);
   U4539 : OAI22_X1 port map( A1 => n3206, A2 => n6207, B1 => n3235, B2 => 
                           n6364, ZN => n6630);
   U4540 : NAND2_X1 port map( A1 => n3207, A2 => CtlToALU_port_pc_reg_10_port, 
                           ZN => n3211);
   U4541 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_10_port, ZN => n3210);
   U4542 : NAND2_X1 port map( A1 => n3208, A2 => CtlToALU_port_imm_10_port, ZN 
                           => n3209);
   U4543 : NAND3_X1 port map( A1 => n3211, A2 => n3210, A3 => n3209, ZN => 
                           IF_ALUxN122);
   U4544 : OAI22_X1 port map( A1 => n4268, A2 => n6337, B1 => n3235, B2 => 
                           n6221, ZN => n6658);
   U4545 : AND2_X1 port map( A1 => n4571, A2 => IF_CPathxpc_reg_signal_16_port,
                           ZN => IF_CPathxN1952);
   U4546 : INV_X1 port map( A => n6390, ZN => n3212);
   U4547 : OAI22_X1 port map( A1 => n3212, A2 => n6207, B1 => n3235, B2 => 
                           n6365, ZN => n6638);
   U4548 : NAND2_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_16_port, 
                           ZN => n3215);
   U4549 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_16_port, ZN => n3214);
   U4550 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_16_port, ZN 
                           => n3213);
   U4551 : NAND3_X1 port map( A1 => n3215, A2 => n3214, A3 => n3213, ZN => 
                           IF_ALUxN128);
   U4552 : AOI22_X1 port map( A1 => n6413, A2 => n6207, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_17_port, ZN => 
                           n3216);
   U4553 : INV_X1 port map( A => n3216, ZN => n6657);
   U4554 : NOR2_X1 port map( A1 => rst, A2 => n6251, ZN => IF_CPathxN1953);
   U4555 : INV_X1 port map( A => n6391, ZN => n3217);
   U4556 : OAI22_X1 port map( A1 => n3217, A2 => n6207, B1 => n4276, B2 => 
                           n6366, ZN => n6608);
   U4557 : NAND2_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_17_port, 
                           ZN => n3220);
   U4558 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_17_port, ZN => n3219);
   U4559 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_17_port, ZN 
                           => n3218);
   U4560 : NAND3_X1 port map( A1 => n3220, A2 => n3219, A3 => n3218, ZN => 
                           IF_ALUxN129);
   U4561 : AOI22_X1 port map( A1 => n6414, A2 => n6207, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_19_port, ZN => 
                           n3221);
   U4562 : INV_X1 port map( A => n3221, ZN => n6655);
   U4563 : NOR2_X1 port map( A1 => rst, A2 => n6252, ZN => IF_CPathxN1955);
   U4564 : INV_X1 port map( A => n6393, ZN => n3222);
   U4565 : OAI22_X1 port map( A1 => n3222, A2 => n4277, B1 => n3235, B2 => 
                           n6367, ZN => n6606);
   U4566 : NAND2_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_19_port, 
                           ZN => n3225);
   U4567 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_19_port, ZN => n3224);
   U4568 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_19_port, ZN 
                           => n3223);
   U4569 : NAND3_X1 port map( A1 => n3225, A2 => n3224, A3 => n3223, ZN => 
                           IF_ALUxN131);
   U4570 : OAI22_X1 port map( A1 => n4268, A2 => n6338, B1 => n4276, B2 => 
                           n6222, ZN => n6656);
   U4571 : AND2_X1 port map( A1 => n4671, A2 => IF_CPathxpc_reg_signal_18_port,
                           ZN => IF_CPathxN1954);
   U4572 : INV_X1 port map( A => n6392, ZN => n3226);
   U4573 : CLKBUF_X1 port map( A => n3235, Z => n4270);
   U4574 : OAI22_X1 port map( A1 => n3226, A2 => n4277, B1 => n4270, B2 => 
                           n6368, ZN => n6602);
   U4575 : NAND2_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_18_port, 
                           ZN => n3229);
   U4576 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_18_port, ZN => n3228);
   U4577 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_18_port, ZN 
                           => n3227);
   U4578 : NAND3_X1 port map( A1 => n3229, A2 => n3228, A3 => n3227, ZN => 
                           IF_ALUxN130);
   U4579 : AOI22_X1 port map( A1 => n6415, A2 => n4277, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_20_port, ZN => 
                           n3230);
   U4580 : INV_X1 port map( A => n3230, ZN => n6654);
   U4581 : AND2_X1 port map( A1 => n6178, A2 => IF_CPathxpc_reg_signal_20_port,
                           ZN => IF_CPathxN1956);
   U4582 : INV_X1 port map( A => n6394, ZN => n3231);
   U4583 : OAI22_X1 port map( A1 => n3231, A2 => n4277, B1 => n4270, B2 => 
                           n6369, ZN => n6622);
   U4584 : NAND2_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_20_port, 
                           ZN => n3234);
   U4585 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_20_port, ZN => n3233);
   U4586 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_20_port, ZN 
                           => n3232);
   U4587 : NAND3_X1 port map( A1 => n3234, A2 => n3233, A3 => n3232, ZN => 
                           IF_ALUxN132);
   U4588 : OAI22_X1 port map( A1 => n4268, A2 => n6339, B1 => n3235, B2 => 
                           n6223, ZN => n6646);
   U4589 : AND2_X1 port map( A1 => n4667, A2 => IF_CPathxpc_reg_signal_28_port,
                           ZN => IF_CPathxN1964);
   U4590 : INV_X1 port map( A => n6402, ZN => n3236);
   U4591 : OAI22_X1 port map( A1 => n3236, A2 => n4277, B1 => n4276, B2 => 
                           n6370, ZN => n6634);
   U4592 : NAND2_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_28_port, 
                           ZN => n3239);
   U4593 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_28_port, ZN => n3238);
   U4594 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_28_port, ZN 
                           => n3237);
   U4595 : NAND3_X1 port map( A1 => n3239, A2 => n3238, A3 => n3237, ZN => 
                           IF_ALUxN140);
   U4596 : AOI22_X1 port map( A1 => n6420, A2 => n6207, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_29_port, ZN => 
                           n3240);
   U4597 : INV_X1 port map( A => n3240, ZN => n6645);
   U4598 : NOR2_X1 port map( A1 => rst, A2 => n6263, ZN => IF_CPathxN1965);
   U4599 : INV_X1 port map( A => n6403, ZN => n3241);
   U4600 : OAI22_X1 port map( A1 => n3241, A2 => n4277, B1 => n4276, B2 => 
                           n6371, ZN => n6632);
   U4601 : NAND2_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_29_port, 
                           ZN => n3245);
   U4602 : NAND2_X1 port map( A1 => n3242, A2 => 
                           CtlToALU_port_reg1_contents_29_port, ZN => n3244);
   U4603 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_29_port, ZN 
                           => n3243);
   U4604 : NAND3_X1 port map( A1 => n3245, A2 => n3244, A3 => n3243, ZN => 
                           IF_ALUxN141);
   U4605 : AOI22_X1 port map( A1 => n6421, A2 => n6207, B1 => n4210, B2 => 
                           IF_CPathxDecToCtl_data_signal_imm_30_port, ZN => 
                           n3246);
   U4606 : INV_X1 port map( A => n3246, ZN => n6644);
   U4607 : AND2_X1 port map( A1 => n4545, A2 => IF_CPathxpc_reg_signal_30_port,
                           ZN => IF_CPathxN1966);
   U4608 : INV_X1 port map( A => n6404, ZN => n3247);
   U4609 : OAI22_X1 port map( A1 => n3247, A2 => n4277, B1 => n4270, B2 => 
                           n6372, ZN => n6580);
   U4610 : NAND2_X1 port map( A1 => n4279, A2 => n6199, ZN => n3735);
   U4611 : NAND2_X1 port map( A1 => n4279, A2 => IF_CPathxmem_en_signal, ZN => 
                           n3251);
   U4612 : INV_X1 port map( A => n3251, ZN => n4413);
   U4613 : NAND2_X1 port map( A1 => ALUtoCtl_port_31_port, A2 => n4413, ZN => 
                           n3249);
   U4614 : OAI211_X1 port map( C1 => n3735, C2 => n3250, A => n3249, B => n3248
                           , ZN => n6435);
   U4615 : NOR2_X1 port map( A1 => rst, A2 => n3250, ZN => IF_CPathxN2273);
   U4616 : INV_X1 port map( A => n3251, ZN => n4415);
   U4617 : NAND2_X1 port map( A1 => ALUtoCtl_port_30_port, A2 => n4415, ZN => 
                           n3253);
   U4618 : OAI211_X1 port map( C1 => n3735, C2 => n3254, A => n3253, B => n3252
                           , ZN => n6437);
   U4619 : INV_X1 port map( A => n3271, ZN => n3953);
   U4620 : NAND2_X1 port map( A1 => n6193, A2 => CtlToALU_port_alu_fun_2_port, 
                           ZN => n4043);
   U4621 : NOR3_X1 port map( A1 => CtlToALU_port_alu_fun_0_port, A2 => 
                           CtlToALU_port_alu_fun_1_port, A3 => n4043, ZN => 
                           n3272);
   U4622 : NAND2_X1 port map( A1 => n3953, A2 => n3272, ZN => n3862);
   U4623 : INV_X1 port map( A => n3782, ZN => n3954);
   U4624 : NOR2_X1 port map( A1 => n3862, A2 => n3954, ZN => n3912);
   U4625 : CLKBUF_X1 port map( A => n3875, Z => n3726);
   U4626 : INV_X1 port map( A => n3726, ZN => n3878);
   U4627 : INV_X1 port map( A => n4118, ZN => n4120);
   U4628 : INV_X1 port map( A => n3487, ZN => n3758);
   U4629 : INV_X1 port map( A => IF_ALUxN134, ZN => n3701);
   U4630 : INV_X1 port map( A => IF_ALUxN133, ZN => n3540);
   U4631 : AOI22_X1 port map( A1 => n3758, A2 => n3701, B1 => n3540, B2 => 
                           n4116, ZN => n3857);
   U4632 : INV_X1 port map( A => IF_ALUxN132, ZN => n3707);
   U4633 : INV_X1 port map( A => IF_ALUxN131, ZN => n4008);
   U4634 : AOI22_X1 port map( A1 => n3758, A2 => n3707, B1 => n4008, B2 => 
                           n4116, ZN => n3720);
   U4635 : INV_X1 port map( A => n4118, ZN => n3725);
   U4636 : INV_X1 port map( A => n3725, ZN => n3856);
   U4637 : AOI22_X1 port map( A1 => n4120, A2 => n3857, B1 => n3720, B2 => 
                           n3856, ZN => n3790);
   U4638 : INV_X1 port map( A => n3487, ZN => n3320);
   U4639 : INV_X1 port map( A => IF_ALUxN130, ZN => n3997);
   U4640 : INV_X1 port map( A => IF_ALUxN129, ZN => n4002);
   U4641 : AOI22_X1 port map( A1 => n3320, A2 => n3997, B1 => n4002, B2 => 
                           n4116, ZN => n3719);
   U4642 : INV_X1 port map( A => IF_ALUxN128, ZN => n4004);
   U4643 : INV_X1 port map( A => IF_ALUxN127, ZN => n3943);
   U4644 : AOI22_X1 port map( A1 => n3320, A2 => n4004, B1 => n3943, B2 => 
                           n4116, ZN => n3722);
   U4645 : AOI22_X1 port map( A1 => n3725, A2 => n3719, B1 => n3722, B2 => 
                           n3856, ZN => n3513);
   U4646 : AOI22_X1 port map( A1 => n3878, A2 => n3790, B1 => n3513, B2 => 
                           n3875, ZN => n3687);
   U4647 : INV_X1 port map( A => n3726, ZN => n3490);
   U4648 : NOR2_X1 port map( A1 => CtlToALU_port_alu_fun_0_port, A2 => 
                           CtlToALU_port_alu_fun_1_port, ZN => n3255);
   U4649 : NAND2_X1 port map( A1 => n3255, A2 => n3263, ZN => n3285);
   U4650 : NOR2_X1 port map( A1 => n3271, A2 => n3285, ZN => n3696);
   U4651 : INV_X1 port map( A => n3696, ZN => n3713);
   U4652 : NOR2_X1 port map( A1 => n4056, A2 => n3713, ZN => n3880);
   U4653 : NAND2_X1 port map( A1 => n3490, A2 => n3880, ZN => n3828);
   U4654 : NAND2_X1 port map( A1 => n3256, A2 => 
                           CtlToALU_port_reg1_contents_31_port, ZN => n3261);
   U4655 : NAND2_X1 port map( A1 => n3257, A2 => CtlToALU_port_pc_reg_31_port, 
                           ZN => n3260);
   U4656 : NAND2_X1 port map( A1 => n3258, A2 => CtlToALU_port_imm_31_port, ZN 
                           => n3259);
   U4657 : NAND3_X1 port map( A1 => n3261, A2 => n3260, A3 => n3259, ZN => 
                           n4144);
   U4658 : INV_X1 port map( A => IF_ALUxN142, ZN => n4041);
   U4659 : AOI21_X1 port map( B1 => n3024, B2 => n4041, A => n4118, ZN => n3265
                           );
   U4660 : OAI21_X1 port map( B1 => n4045, B2 => n4144, A => n3265, ZN => n3286
                           );
   U4661 : NOR2_X1 port map( A1 => n6201, A2 => n6246, ZN => n3262);
   U4662 : NAND2_X1 port map( A1 => n3263, A2 => n3262, ZN => n4131);
   U4663 : INV_X1 port map( A => n4131, ZN => n4073);
   U4664 : INV_X1 port map( A => n4040, ZN => n3279);
   U4665 : NAND2_X1 port map( A1 => n3279, A2 => IF_ALUxN142, ZN => n4038);
   U4666 : OAI21_X1 port map( B1 => n3279, B2 => IF_ALUxN142, A => n4038, ZN =>
                           n3268);
   U4667 : INV_X1 port map( A => n4043, ZN => n3928);
   U4668 : NAND3_X1 port map( A1 => CtlToALU_port_alu_fun_0_port, A2 => 
                           CtlToALU_port_alu_fun_1_port, A3 => n3928, ZN => 
                           n4122);
   U4669 : NOR2_X1 port map( A1 => n3953, A2 => n4122, ZN => n4063);
   U4670 : NAND2_X1 port map( A1 => n4144, A2 => n4063, ZN => n3882);
   U4671 : INV_X1 port map( A => n3882, ZN => n3908);
   U4672 : INV_X1 port map( A => IF_ALUxN138, ZN => n3798);
   U4673 : INV_X1 port map( A => IF_ALUxN137, ZN => n3330);
   U4674 : AOI22_X1 port map( A1 => n3758, A2 => n3798, B1 => n3330, B2 => 
                           n4116, ZN => n3859);
   U4675 : INV_X1 port map( A => IF_ALUxN136, ZN => n3897);
   U4676 : INV_X1 port map( A => IF_ALUxN135, ZN => n3679);
   U4677 : AOI22_X1 port map( A1 => n3758, A2 => n3897, B1 => n3679, B2 => 
                           n4116, ZN => n3858);
   U4678 : AOI22_X1 port map( A1 => n4120, A2 => n3859, B1 => n3858, B2 => 
                           n3856, ZN => n3789);
   U4679 : NOR2_X1 port map( A1 => n4056, A2 => n3490, ZN => n3864);
   U4680 : INV_X1 port map( A => n3864, ZN => n4053);
   U4681 : NOR2_X1 port map( A1 => n3862, A2 => n4053, ZN => n4141);
   U4682 : INV_X1 port map( A => n4141, ZN => n3886);
   U4683 : INV_X1 port map( A => IF_ALUxN141, ZN => n3839);
   U4684 : NAND2_X1 port map( A1 => n3839, A2 => n4116, ZN => n3264);
   U4685 : INV_X1 port map( A => IF_ALUxN140, ZN => n4033);
   U4686 : INV_X1 port map( A => IF_ALUxN139, ZN => n3775);
   U4687 : AOI22_X1 port map( A1 => n3758, A2 => n4033, B1 => n3775, B2 => 
                           n4116, ZN => n3861);
   U4688 : AOI22_X1 port map( A1 => n3265, A2 => n3264, B1 => n3861, B2 => 
                           n3856, ZN => n3266);
   U4689 : INV_X1 port map( A => n3862, ZN => n3636);
   U4690 : NAND2_X1 port map( A1 => n3954, A2 => n3636, ZN => n3671);
   U4691 : NOR2_X1 port map( A1 => n3726, A2 => n3671, ZN => n3761);
   U4692 : INV_X1 port map( A => n3761, ZN => n4117);
   U4693 : OAI22_X1 port map( A1 => n3789, A2 => n3886, B1 => n3266, B2 => 
                           n4117, ZN => n3267);
   U4694 : AOI211_X1 port map( C1 => n4073, C2 => n3268, A => n3908, B => n3267
                           , ZN => n3270);
   U4695 : NOR2_X2 port map( A1 => CtlToALU_port_alu_fun_2_port, A2 => 
                           CtlToALU_port_alu_fun_3_port, ZN => n4060);
   U4696 : OAI221_X1 port map( B1 => IF_ALUxN142, B2 => 
                           CtlToALU_port_alu_fun_0_port, C1 => IF_ALUxN142, C2 
                           => n4040, A => n4060, ZN => n3269);
   U4697 : OAI211_X1 port map( C1 => n3828, C2 => n3286, A => n3270, B => n3269
                           , ZN => n3274);
   U4698 : INV_X1 port map( A => n3725, ZN => n3494);
   U4699 : NAND2_X1 port map( A1 => n3494, A2 => n4144, ZN => n3375);
   U4700 : NAND2_X1 port map( A1 => n3875, A2 => n4144, ZN => n3491);
   U4701 : OAI211_X1 port map( C1 => n3286, C2 => n3875, A => n3375, B => n3491
                           , ZN => n3292);
   U4702 : INV_X1 port map( A => n4144, ZN => n4147);
   U4703 : NOR2_X1 port map( A1 => n3866, A2 => n4147, ZN => n3743);
   U4704 : AOI21_X1 port map( B1 => n3954, B2 => n3292, A => n3743, ZN => n3464
                           );
   U4705 : NOR2_X1 port map( A1 => n4122, A2 => n3271, ZN => n3891);
   U4706 : INV_X1 port map( A => n3891, ZN => n3851);
   U4707 : INV_X1 port map( A => n4118, ZN => n3860);
   U4708 : INV_X1 port map( A => IF_ALUxN126, ZN => n3941);
   U4709 : INV_X1 port map( A => IF_ALUxN125, ZN => n3617);
   U4710 : AOI22_X1 port map( A1 => n3320, A2 => n3941, B1 => n3617, B2 => 
                           n4116, ZN => n3721);
   U4711 : INV_X1 port map( A => IF_ALUxN124, ZN => n3751);
   U4712 : INV_X1 port map( A => IF_ALUxN123, ZN => n3638);
   U4713 : AOI22_X1 port map( A1 => n3320, A2 => n3751, B1 => n3638, B2 => 
                           n4116, ZN => n3724);
   U4714 : AOI22_X1 port map( A1 => n3860, A2 => n3721, B1 => n3724, B2 => 
                           n3856, ZN => n3512);
   U4715 : INV_X1 port map( A => IF_ALUxN122, ZN => n3983);
   U4716 : INV_X1 port map( A => IF_ALUxN121, ZN => n3950);
   U4717 : AOI22_X1 port map( A1 => n3024, A2 => n3983, B1 => n3950, B2 => 
                           n4116, ZN => n3723);
   U4718 : INV_X1 port map( A => IF_ALUxN120, ZN => n3952);
   U4719 : INV_X1 port map( A => IF_ALUxN119, ZN => n3976);
   U4720 : AOI22_X1 port map( A1 => n3320, A2 => n3952, B1 => n3976, B2 => 
                           n4116, ZN => n3651);
   U4721 : AOI22_X1 port map( A1 => n3725, A2 => n3723, B1 => n3651, B2 => 
                           n3856, ZN => n3510);
   U4722 : AOI22_X1 port map( A1 => n3878, A2 => n3512, B1 => n3510, B2 => 
                           n3726, ZN => n3686);
   U4723 : INV_X1 port map( A => IF_ALUxN118, ZN => n3966);
   U4724 : INV_X1 port map( A => IF_ALUxN117, ZN => n3968);
   U4725 : AOI22_X1 port map( A1 => n3758, A2 => n3966, B1 => n3968, B2 => 
                           n3487, ZN => n3650);
   U4726 : INV_X1 port map( A => IF_ALUxN116, ZN => n3503);
   U4727 : INV_X1 port map( A => IF_ALUxN115, ZN => n3428);
   U4728 : AOI22_X1 port map( A1 => n3758, A2 => n3503, B1 => n3428, B2 => 
                           n3487, ZN => n3485);
   U4729 : AOI22_X1 port map( A1 => n3860, A2 => n3650, B1 => n3485, B2 => 
                           n3856, ZN => n3509);
   U4730 : INV_X1 port map( A => IF_ALUxN114, ZN => n3440);
   U4731 : OAI22_X1 port map( A1 => n4116, A2 => n3440, B1 => n3407, B2 => 
                           n3024, ZN => n3484);
   U4732 : AND2_X1 port map( A1 => IF_ALUxN112, A2 => n4045, ZN => n3927);
   U4733 : OAI22_X1 port map( A1 => n4118, A2 => n3484, B1 => n3927, B2 => 
                           n3860, ZN => n3441);
   U4734 : AOI22_X1 port map( A1 => n3878, A2 => n3509, B1 => n3441, B2 => 
                           n3875, ZN => n3690);
   U4735 : AOI22_X1 port map( A1 => n3866, A2 => n3686, B1 => n3690, B2 => 
                           n3782, ZN => n3463);
   U4736 : NAND2_X1 port map( A1 => n3272, A2 => n3271, ZN => n3894);
   U4737 : OAI22_X1 port map( A1 => n3464, A2 => n3851, B1 => n3463, B2 => 
                           n3894, ZN => n3273);
   U4738 : AOI211_X1 port map( C1 => n3912, C2 => n3687, A => n3274, B => n3273
                           , ZN => n3282);
   U4739 : NOR2_X1 port map( A1 => CtlToALU_port_alu_fun_1_port, A2 => n6201, 
                           ZN => n3929);
   U4740 : INV_X1 port map( A => n3929, ZN => n3275);
   U4741 : NAND3_X1 port map( A1 => n4060, A2 => n6246, A3 => n6201, ZN => 
                           n3278);
   U4742 : OAI211_X1 port map( C1 => CtlToALU_port_alu_fun_2_port, C2 => n3275,
                           A => n4667, B => n3278, ZN => n4154);
   U4743 : CLKBUF_X1 port map( A => n4154, Z => n4078);
   U4744 : INV_X1 port map( A => n3276, ZN => n3277);
   U4745 : AOI21_X1 port map( B1 => n3278, B2 => n3277, A => rst, ZN => n3640);
   U4746 : CLKBUF_X1 port map( A => n3640, Z => n4152);
   U4747 : NAND4_X1 port map( A1 => n3929, A2 => n4571, A3 => n6193, A4 => 
                           n6268, ZN => n3816);
   U4748 : NOR3_X1 port map( A1 => n3279, A2 => n4041, A3 => n3816, ZN => n3280
                           );
   U4749 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_30, A => n3280, ZN 
                           => n3281);
   U4750 : OAI21_X1 port map( B1 => n3282, B2 => n4078, A => n3281, ZN => 
                           IF_ALUxN968);
   U4751 : NAND2_X1 port map( A1 => ALUtoCtl_port_6_port, A2 => n4415, ZN => 
                           n3284);
   U4752 : OAI211_X1 port map( C1 => n3735, C2 => n4108, A => n3284, B => n3283
                           , ZN => n6439);
   U4753 : NOR2_X1 port map( A1 => n3953, A2 => n3285, ZN => n4062);
   U4754 : INV_X1 port map( A => n3286, ZN => n3436);
   U4755 : NAND2_X1 port map( A1 => n3490, A2 => n3436, ZN => n3460);
   U4756 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN134, B1 => IF_ALUxN135
                           , B2 => n3487, ZN => n3492);
   U4757 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN136, B1 => IF_ALUxN137
                           , B2 => n3487, ZN => n3496);
   U4758 : AOI22_X1 port map( A1 => n3860, A2 => n3492, B1 => n3496, B2 => 
                           n3494, ZN => n3434);
   U4759 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN138, B1 => IF_ALUxN139
                           , B2 => n3487, ZN => n3495);
   U4760 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN140, B1 => IF_ALUxN141
                           , B2 => n4116, ZN => n3489);
   U4761 : AOI22_X1 port map( A1 => n3860, A2 => n3495, B1 => n3489, B2 => 
                           n3856, ZN => n3287);
   U4762 : MUX2_X1 port map( A => n3434, B => n3287, S => n3875, Z => n3288);
   U4763 : INV_X1 port map( A => n3288, ZN => n3457);
   U4764 : NOR2_X1 port map( A1 => n4056, A2 => n3457, ZN => n3291);
   U4765 : INV_X1 port map( A => n3291, ZN => n3289);
   U4766 : OAI21_X1 port map( B1 => n3954, B2 => n3460, A => n3289, ZN => n3695
                           );
   U4767 : AOI22_X1 port map( A1 => n3024, A2 => IF_ALUxN126, B1 => IF_ALUxN127
                           , B2 => n3487, ZN => n3475);
   U4768 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN128, B1 => IF_ALUxN129
                           , B2 => n3487, ZN => n3478);
   U4769 : AOI22_X1 port map( A1 => n3725, A2 => n3475, B1 => n3478, B2 => 
                           n3494, ZN => n3443);
   U4770 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN130, B1 => IF_ALUxN131
                           , B2 => n3487, ZN => n3477);
   U4771 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN132, B1 => IF_ALUxN133
                           , B2 => n3487, ZN => n3493);
   U4772 : AOI22_X1 port map( A1 => n3725, A2 => n3477, B1 => n3493, B2 => 
                           n3494, ZN => n3435);
   U4773 : AOI22_X1 port map( A1 => n3490, A2 => n3443, B1 => n3435, B2 => 
                           n3726, ZN => n3458);
   U4774 : NOR2_X2 port map( A1 => n3696, A2 => n3891, ZN => n4055);
   U4775 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN122, B1 => IF_ALUxN123
                           , B2 => n3487, ZN => n3479);
   U4776 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN124, B1 => IF_ALUxN125
                           , B2 => n3487, ZN => n3476);
   U4777 : AOI22_X1 port map( A1 => n3725, A2 => n3479, B1 => n3476, B2 => 
                           n3494, ZN => n3444);
   U4778 : NAND2_X1 port map( A1 => n3954, A2 => n3878, ZN => n4051);
   U4779 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN118, B1 => IF_ALUxN119
                           , B2 => n3487, ZN => n3481);
   U4780 : AOI22_X1 port map( A1 => n3024, A2 => IF_ALUxN120, B1 => IF_ALUxN121
                           , B2 => n3487, ZN => n3480);
   U4781 : AOI22_X1 port map( A1 => n3725, A2 => n3481, B1 => n3480, B2 => 
                           n3856, ZN => n3446);
   U4782 : OAI22_X1 port map( A1 => n4053, A2 => n3444, B1 => n4051, B2 => 
                           n3446, ZN => n3290);
   U4783 : AOI211_X1 port map( C1 => n3458, C2 => n4056, A => n4055, B => n3290
                           , ZN => n3297);
   U4784 : AOI21_X1 port map( B1 => n3782, B2 => n3292, A => n3291, ZN => n3699
                           );
   U4785 : INV_X1 port map( A => n4063, ZN => n3747);
   U4786 : NAND2_X1 port map( A1 => CtlToALU_port_alu_fun_0_port, A2 => n4060, 
                           ZN => n4079);
   U4787 : INV_X1 port map( A => n4079, ZN => n4127);
   U4788 : INV_X1 port map( A => n3671, ZN => n3914);
   U4789 : AOI22_X1 port map( A1 => n4127, A2 => n3965, B1 => n3914, B2 => 
                           n3690, ZN => n3295);
   U4790 : NAND2_X1 port map( A1 => n3966, A2 => n3965, ZN => n3969);
   U4791 : OAI21_X1 port map( B1 => n3966, B2 => n3965, A => n3969, ZN => n3293
                           );
   U4792 : AOI22_X1 port map( A1 => n4060, A2 => IF_ALUxN118, B1 => n4073, B2 
                           => n3293, ZN => n3294);
   U4793 : OAI211_X1 port map( C1 => n3699, C2 => n3747, A => n3295, B => n3294
                           , ZN => n3296);
   U4794 : AOI211_X1 port map( C1 => n4062, C2 => n3695, A => n3297, B => n3296
                           , ZN => n3301);
   U4795 : CLKBUF_X1 port map( A => n3816, Z => n4148);
   U4796 : NOR3_X1 port map( A1 => n3298, A2 => n4148, A3 => n3966, ZN => n3299
                           );
   U4797 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_6, A => n3299, ZN 
                           => n3300);
   U4798 : OAI21_X1 port map( B1 => n3301, B2 => n4078, A => n3300, ZN => 
                           IF_ALUxN944);
   U4799 : NAND2_X1 port map( A1 => ALUtoCtl_port_9_port, A2 => n4415, ZN => 
                           n3303);
   U4800 : OAI211_X1 port map( C1 => n3735, C2 => n4105, A => n3303, B => n3302
                           , ZN => n6441);
   U4801 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN121, B1 => IF_ALUxN120
                           , B2 => n4116, ZN => n3556);
   U4802 : OAI22_X1 port map( A1 => n4116, A2 => IF_ALUxN119, B1 => IF_ALUxN118
                           , B2 => n4045, ZN => n3352);
   U4803 : AOI22_X1 port map( A1 => n3725, A2 => n3556, B1 => n3352, B2 => 
                           n3856, ZN => n3528);
   U4804 : AOI22_X1 port map( A1 => n4045, A2 => IF_ALUxN117, B1 => IF_ALUxN116
                           , B2 => n4116, ZN => n3351);
   U4805 : AOI22_X1 port map( A1 => n3320, A2 => n3428, B1 => n3440, B2 => 
                           n3487, ZN => n3354);
   U4806 : INV_X1 port map( A => n3354, ZN => n3304);
   U4807 : AOI22_X1 port map( A1 => n3860, A2 => n3351, B1 => n3304, B2 => 
                           n3494, ZN => n3372);
   U4808 : AOI22_X1 port map( A1 => n3878, A2 => n3528, B1 => n3372, B2 => 
                           n3726, ZN => n3576);
   U4809 : NAND2_X1 port map( A1 => n3782, A2 => n3878, ZN => n3625);
   U4810 : NAND2_X1 port map( A1 => IF_ALUxN112, A2 => n4116, ZN => n3926);
   U4811 : OAI21_X1 port map( B1 => n3407, B2 => n4116, A => n3926, ZN => n3353
                           );
   U4812 : NAND2_X1 port map( A1 => n3860, A2 => n3353, ZN => n3397);
   U4813 : OAI22_X1 port map( A1 => n3576, A2 => n3782, B1 => n3625, B2 => 
                           n3397, ZN => n3325);
   U4814 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN121, B1 => IF_ALUxN122
                           , B2 => n4116, ZN => n3345);
   U4815 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN123, B1 => IF_ALUxN124
                           , B2 => n4116, ZN => n3347);
   U4816 : AOI22_X1 port map( A1 => n4120, A2 => n3345, B1 => n3347, B2 => 
                           n3494, ZN => n3370);
   U4817 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN125, B1 => IF_ALUxN126
                           , B2 => n4116, ZN => n3346);
   U4818 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN127, B1 => IF_ALUxN128
                           , B2 => n4116, ZN => n3342);
   U4819 : AOI22_X1 port map( A1 => n4120, A2 => n3346, B1 => n3342, B2 => 
                           n3494, ZN => n3368);
   U4820 : AOI22_X1 port map( A1 => n3490, A2 => n3370, B1 => n3368, B2 => 
                           n3726, ZN => n3395);
   U4821 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN129, B1 => IF_ALUxN130
                           , B2 => n4116, ZN => n3341);
   U4822 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN131, B1 => IF_ALUxN132
                           , B2 => n4116, ZN => n3344);
   U4823 : AOI22_X1 port map( A1 => n3725, A2 => n3341, B1 => n3344, B2 => 
                           n3494, ZN => n3367);
   U4824 : AOI22_X1 port map( A1 => n4045, A2 => IF_ALUxN133, B1 => IF_ALUxN134
                           , B2 => n4116, ZN => n3343);
   U4825 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN135, B1 => IF_ALUxN136
                           , B2 => n4116, ZN => n3340);
   U4826 : AOI22_X1 port map( A1 => n3860, A2 => n3343, B1 => n3340, B2 => 
                           n3494, ZN => n3378);
   U4827 : AOI22_X1 port map( A1 => n3490, A2 => n3367, B1 => n3378, B2 => 
                           n3875, ZN => n3399);
   U4828 : AOI221_X1 port map( B1 => n3866, B2 => n3395, C1 => n3782, C2 => 
                           n3399, A => n4055, ZN => n3311);
   U4829 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN141, B1 => IF_ALUxN142
                           , B2 => n4116, ZN => n3337);
   U4830 : NOR2_X1 port map( A1 => n3337, A2 => n4118, ZN => n3374);
   U4831 : INV_X1 port map( A => n3375, ZN => n3438);
   U4832 : NOR3_X1 port map( A1 => n3374, A2 => n3878, A3 => n3438, ZN => n3305
                           );
   U4833 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN137, B1 => IF_ALUxN138
                           , B2 => n4116, ZN => n3339);
   U4834 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN139, B1 => IF_ALUxN140
                           , B2 => n4116, ZN => n3338);
   U4835 : AOI22_X1 port map( A1 => n3860, A2 => n3339, B1 => n3338, B2 => 
                           n3494, ZN => n3377);
   U4836 : NOR2_X1 port map( A1 => n3377, A2 => n3875, ZN => n3306);
   U4837 : NOR2_X1 port map( A1 => n3305, A2 => n3306, ZN => n3400);
   U4838 : AOI21_X1 port map( B1 => n3954, B2 => n3400, A => n3743, ZN => n3328
                           );
   U4839 : NAND2_X1 port map( A1 => n3954, A2 => n4062, ZN => n3461);
   U4840 : INV_X1 port map( A => n3461, ZN => n3806);
   U4841 : NOR2_X1 port map( A1 => n4147, A2 => n4116, ZN => n4115);
   U4842 : AOI21_X1 port map( B1 => n4115, B2 => n4118, A => n3374, ZN => n3379
                           );
   U4843 : AOI21_X1 port map( B1 => n3379, B2 => n3875, A => n3306, ZN => n3402
                           );
   U4844 : AOI22_X1 port map( A1 => n4127, A2 => n3949, B1 => n3806, B2 => 
                           n3402, ZN => n3309);
   U4845 : INV_X1 port map( A => n3949, ZN => n3312);
   U4846 : NAND2_X1 port map( A1 => n3312, A2 => IF_ALUxN121, ZN => n3981);
   U4847 : OAI21_X1 port map( B1 => n3312, B2 => IF_ALUxN121, A => n3981, ZN =>
                           n3307);
   U4848 : AOI22_X1 port map( A1 => n4060, A2 => IF_ALUxN121, B1 => n4073, B2 
                           => n3307, ZN => n3308);
   U4849 : OAI211_X1 port map( C1 => n3328, C2 => n3747, A => n3309, B => n3308
                           , ZN => n3310);
   U4850 : AOI211_X1 port map( C1 => n3636, C2 => n3325, A => n3311, B => n3310
                           , ZN => n3315);
   U4851 : NOR3_X1 port map( A1 => n3950, A2 => n3312, A3 => n3816, ZN => n3313
                           );
   U4852 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_9, A => n3313, ZN 
                           => n3314);
   U4853 : OAI21_X1 port map( B1 => n3315, B2 => n4154, A => n3314, ZN => 
                           IF_ALUxN947);
   U4854 : NAND2_X1 port map( A1 => ALUtoCtl_port_25_port, A2 => n4415, ZN => 
                           n3317);
   U4855 : OAI211_X1 port map( C1 => n3735, C2 => n4089, A => n3317, B => n3316
                           , ZN => n6443);
   U4856 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN129, B1 => IF_ALUxN128
                           , B2 => n4116, ZN => n3548);
   U4857 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN127, B1 => IF_ALUxN126
                           , B2 => n4116, ZN => n3551);
   U4858 : AOI22_X1 port map( A1 => n3725, A2 => n3548, B1 => n3551, B2 => 
                           n3494, ZN => n3530);
   U4859 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN125, B1 => IF_ALUxN124
                           , B2 => n4116, ZN => n3550);
   U4860 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN123, B1 => IF_ALUxN122
                           , B2 => n4116, ZN => n3557);
   U4861 : AOI22_X1 port map( A1 => n3725, A2 => n3550, B1 => n3557, B2 => 
                           n3856, ZN => n3529);
   U4862 : AOI22_X1 port map( A1 => n3878, A2 => n3530, B1 => n3529, B2 => 
                           n3726, ZN => n3574);
   U4863 : INV_X1 port map( A => n3574, ZN => n3318);
   U4864 : AOI22_X1 port map( A1 => n3402, A2 => n3880, B1 => n3912, B2 => 
                           n3318, ZN => n3327);
   U4865 : INV_X1 port map( A => n3894, ZN => n4135);
   U4866 : OR2_X1 port map( A1 => n3319, A2 => n3330, ZN => n4023);
   U4867 : NAND2_X1 port map( A1 => n3319, A2 => n3330, ZN => n3933);
   U4868 : AOI21_X1 port map( B1 => n4023, B2 => n3933, A => n4131, ZN => n3324
                           );
   U4869 : AOI21_X1 port map( B1 => CtlToALU_port_alu_fun_0_port, B2 => n3319, 
                           A => IF_ALUxN137, ZN => n3322);
   U4870 : INV_X1 port map( A => n4060, ZN => n4123);
   U4871 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN137, B1 => IF_ALUxN136
                           , B2 => n4116, ZN => n3759);
   U4872 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN135, B1 => IF_ALUxN134
                           , B2 => n4116, ZN => n3667);
   U4873 : AOI22_X1 port map( A1 => n3725, A2 => n3759, B1 => n3667, B2 => 
                           n3856, ZN => n3825);
   U4874 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN133, B1 => IF_ALUxN132
                           , B2 => n4116, ZN => n3666);
   U4875 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN131, B1 => IF_ALUxN130
                           , B2 => n4116, ZN => n3549);
   U4876 : AOI22_X1 port map( A1 => n3725, A2 => n3666, B1 => n3549, B2 => 
                           n3856, ZN => n3531);
   U4877 : AOI22_X1 port map( A1 => n3761, A2 => n3825, B1 => n3531, B2 => 
                           n4141, ZN => n3321);
   U4878 : OAI211_X1 port map( C1 => n3322, C2 => n4123, A => n3321, B => n3882
                           , ZN => n3323);
   U4879 : AOI211_X1 port map( C1 => n4135, C2 => n3325, A => n3324, B => n3323
                           , ZN => n3326);
   U4880 : OAI211_X1 port map( C1 => n3328, C2 => n3851, A => n3327, B => n3326
                           , ZN => n3329);
   U4881 : INV_X1 port map( A => n3329, ZN => n3334);
   U4882 : NOR3_X1 port map( A1 => n3331, A2 => n4148, A3 => n3330, ZN => n3332
                           );
   U4883 : AOI21_X1 port map( B1 => n3640, B2 => C596xDATA2_25, A => n3332, ZN 
                           => n3333);
   U4884 : OAI21_X1 port map( B1 => n4078, B2 => n3334, A => n3333, ZN => 
                           IF_ALUxN963);
   U4885 : NAND2_X1 port map( A1 => ALUtoCtl_port_7_port, A2 => n4415, ZN => 
                           n3336);
   U4886 : OAI211_X1 port map( C1 => n3735, C2 => n4107, A => n3336, B => n3335
                           , ZN => n6445);
   U4887 : INV_X1 port map( A => n3743, ZN => n3781);
   U4888 : AOI22_X1 port map( A1 => n3860, A2 => n3338, B1 => n3337, B2 => 
                           n3856, ZN => n3591);
   U4889 : AOI22_X1 port map( A1 => n3725, A2 => n3340, B1 => n3339, B2 => 
                           n3856, ZN => n3592);
   U4890 : OAI221_X1 port map( B1 => n3490, B2 => n3591, C1 => n3726, C2 => 
                           n3592, A => n3866, ZN => n3349);
   U4891 : NAND2_X1 port map( A1 => n3781, A2 => n3349, ZN => n3678);
   U4892 : AOI22_X1 port map( A1 => n3860, A2 => n3342, B1 => n3341, B2 => 
                           n3856, ZN => n3413);
   U4893 : AOI22_X1 port map( A1 => n3860, A2 => n3344, B1 => n3343, B2 => 
                           n3856, ZN => n3421);
   U4894 : AOI22_X1 port map( A1 => n3490, A2 => n3413, B1 => n3421, B2 => 
                           n3875, ZN => n3594);
   U4895 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN119, B1 => IF_ALUxN120
                           , B2 => n4116, ZN => n3369);
   U4896 : AOI22_X1 port map( A1 => n4120, A2 => n3369, B1 => n3345, B2 => 
                           n3494, ZN => n3418);
   U4897 : AOI22_X1 port map( A1 => n3860, A2 => n3347, B1 => n3346, B2 => 
                           n3494, ZN => n3414);
   U4898 : OAI22_X1 port map( A1 => n3418, A2 => n4051, B1 => n3414, B2 => 
                           n4053, ZN => n3348);
   U4899 : AOI211_X1 port map( C1 => n3782, C2 => n3594, A => n4055, B => n3348
                           , ZN => n3360);
   U4900 : NAND2_X1 port map( A1 => n3860, A2 => n4115, ZN => n3590);
   U4901 : OAI21_X1 port map( B1 => n3590, B2 => n3625, A => n3349, ZN => n3350
                           );
   U4902 : INV_X1 port map( A => n3350, ZN => n3675);
   U4903 : INV_X1 port map( A => n4062, ZN => n3589);
   U4904 : OAI22_X1 port map( A1 => n4118, A2 => n3352, B1 => n3351, B2 => 
                           n3860, ZN => n3558);
   U4905 : AOI22_X1 port map( A1 => n3725, A2 => n3354, B1 => n3353, B2 => 
                           n3856, ZN => n3624);
   U4906 : INV_X1 port map( A => n3624, ZN => n3553);
   U4907 : OAI22_X1 port map( A1 => n3875, A2 => n3558, B1 => n3553, B2 => 
                           n3490, ZN => n3664);
   U4908 : INV_X1 port map( A => n3664, ZN => n3355);
   U4909 : AOI22_X1 port map( A1 => n4127, A2 => n3975, B1 => n3914, B2 => 
                           n3355, ZN => n3358);
   U4910 : NAND2_X1 port map( A1 => n3976, A2 => n3975, ZN => n3970);
   U4911 : OAI21_X1 port map( B1 => n3976, B2 => n3975, A => n3970, ZN => n3356
                           );
   U4912 : AOI22_X1 port map( A1 => n4060, A2 => IF_ALUxN119, B1 => n4073, B2 
                           => n3356, ZN => n3357);
   U4913 : OAI211_X1 port map( C1 => n3675, C2 => n3589, A => n3358, B => n3357
                           , ZN => n3359);
   U4914 : AOI211_X1 port map( C1 => n4063, C2 => n3678, A => n3360, B => n3359
                           , ZN => n3364);
   U4915 : NOR3_X1 port map( A1 => n3361, A2 => n3816, A3 => n3976, ZN => n3362
                           );
   U4916 : AOI21_X1 port map( B1 => n3640, B2 => C596xDATA2_7, A => n3362, ZN 
                           => n3363);
   U4917 : OAI21_X1 port map( B1 => n3364, B2 => n4154, A => n3363, ZN => 
                           IF_ALUxN945);
   U4918 : NAND2_X1 port map( A1 => ALUtoCtl_port_5_port, A2 => n4415, ZN => 
                           n3366);
   U4919 : OAI211_X1 port map( C1 => n3735, C2 => n4109, A => n3366, B => n3365
                           , ZN => n6447);
   U4920 : AOI22_X1 port map( A1 => n3490, A2 => n3368, B1 => n3367, B2 => 
                           n3875, ZN => n3606);
   U4921 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN117, B1 => IF_ALUxN118
                           , B2 => n4116, ZN => n3415);
   U4922 : AOI22_X1 port map( A1 => n3860, A2 => n3415, B1 => n3369, B2 => 
                           n3494, ZN => n3393);
   U4923 : OAI22_X1 port map( A1 => n3393, A2 => n4051, B1 => n3370, B2 => 
                           n4053, ZN => n3371);
   U4924 : AOI211_X1 port map( C1 => n4056, C2 => n3606, A => n4055, B => n3371
                           , ZN => n3384);
   U4925 : INV_X1 port map( A => n3967, ZN => n3385);
   U4926 : INV_X1 port map( A => n3397, ZN => n3571);
   U4927 : AOI22_X1 port map( A1 => n3490, A2 => n3372, B1 => n3571, B2 => 
                           n3875, ZN => n3604);
   U4928 : OAI22_X1 port map( A1 => n3385, A2 => n4079, B1 => n3604, B2 => 
                           n3671, ZN => n3383);
   U4929 : NOR2_X1 port map( A1 => n3385, A2 => IF_ALUxN117, ZN => n3962);
   U4930 : AOI21_X1 port map( B1 => n3385, B2 => IF_ALUxN117, A => n3962, ZN =>
                           n3373);
   U4931 : OAI22_X1 port map( A1 => n3968, A2 => n4123, B1 => n3373, B2 => 
                           n4131, ZN => n3382);
   U4932 : INV_X1 port map( A => n3374, ZN => n3376);
   U4933 : OAI211_X1 port map( C1 => n3875, C2 => n3376, A => n3375, B => n3491
                           , ZN => n3608);
   U4934 : AOI22_X1 port map( A1 => n3490, A2 => n3378, B1 => n3377, B2 => 
                           n3726, ZN => n3607);
   U4935 : NOR2_X1 port map( A1 => n3607, A2 => n3782, ZN => n3380);
   U4936 : AOI21_X1 port map( B1 => n3782, B2 => n3608, A => n3380, ZN => n3536
                           );
   U4937 : INV_X1 port map( A => n3625, ZN => n3785);
   U4938 : INV_X1 port map( A => n3379, ZN => n3832);
   U4939 : AOI21_X1 port map( B1 => n3785, B2 => n3832, A => n3380, ZN => n3535
                           );
   U4940 : OAI22_X1 port map( A1 => n3536, A2 => n3747, B1 => n3535, B2 => 
                           n3589, ZN => n3381);
   U4941 : NOR4_X1 port map( A1 => n3384, A2 => n3383, A3 => n3382, A4 => n3381
                           , ZN => n3388);
   U4942 : NOR3_X1 port map( A1 => n3385, A2 => n3968, A3 => n3816, ZN => n3386
                           );
   U4943 : AOI21_X1 port map( B1 => n3640, B2 => C596xDATA2_5, A => n3386, ZN 
                           => n3387);
   U4944 : OAI21_X1 port map( B1 => n3388, B2 => n4154, A => n3387, ZN => 
                           IF_ALUxN943);
   U4945 : NAND2_X1 port map( A1 => ALUtoCtl_port_1_port, A2 => n4415, ZN => 
                           n3390);
   U4946 : OAI211_X1 port map( C1 => n3735, C2 => n4113, A => n3390, B => n3389
                           , ZN => n6449);
   U4947 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN113, B1 => IF_ALUxN114
                           , B2 => n4116, ZN => n3391);
   U4948 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN115, B1 => IF_ALUxN116
                           , B2 => n4116, ZN => n3416);
   U4949 : AOI22_X1 port map( A1 => n3725, A2 => n3391, B1 => n3416, B2 => 
                           n3494, ZN => n3392);
   U4950 : OAI22_X1 port map( A1 => n3393, A2 => n4053, B1 => n4051, B2 => 
                           n3392, ZN => n3394);
   U4951 : AOI211_X1 port map( C1 => n4056, C2 => n3395, A => n4055, B => n3394
                           , ZN => n3406);
   U4952 : NAND2_X1 port map( A1 => n3860, A2 => IF_ALUxN113, ZN => n3955);
   U4953 : NOR2_X1 port map( A1 => n3725, A2 => IF_ALUxN113, ZN => n3958);
   U4954 : INV_X1 port map( A => n3958, ZN => n3396);
   U4955 : AOI21_X1 port map( B1 => n3955, B2 => n3396, A => n4131, ZN => n3405
                           );
   U4956 : AOI21_X1 port map( B1 => CtlToALU_port_alu_fun_0_port, B2 => n4118, 
                           A => IF_ALUxN113, ZN => n3398);
   U4957 : OAI22_X1 port map( A1 => n3398, A2 => n4123, B1 => n4117, B2 => 
                           n3397, ZN => n3404);
   U4958 : NAND2_X1 port map( A1 => n3954, A2 => n3399, ZN => n3401);
   U4959 : OAI21_X1 port map( B1 => n3954, B2 => n3400, A => n3401, ZN => n3575
                           );
   U4960 : OAI21_X1 port map( B1 => n3954, B2 => n3402, A => n3401, ZN => n3568
                           );
   U4961 : OAI22_X1 port map( A1 => n3747, A2 => n3575, B1 => n3589, B2 => 
                           n3568, ZN => n3403);
   U4962 : NOR4_X1 port map( A1 => n3406, A2 => n3405, A3 => n3404, A4 => n3403
                           , ZN => n3410);
   U4963 : NOR3_X1 port map( A1 => n3407, A2 => n3816, A3 => n3725, ZN => n3408
                           );
   U4964 : AOI21_X1 port map( B1 => n3640, B2 => C596xDATA2_1, A => n3408, ZN 
                           => n3409);
   U4965 : OAI21_X1 port map( B1 => n3410, B2 => n4154, A => n3409, ZN => 
                           IF_ALUxN939);
   U4966 : NAND2_X1 port map( A1 => ALUtoCtl_port_3_port, A2 => n4415, ZN => 
                           n3412);
   U4967 : OAI211_X1 port map( C1 => n3735, C2 => n4111, A => n3412, B => n3411
                           , ZN => n6451);
   U4968 : AOI22_X1 port map( A1 => n3490, A2 => n3414, B1 => n3413, B2 => 
                           n3875, ZN => n3628);
   U4969 : AOI22_X1 port map( A1 => n4120, A2 => n3416, B1 => n3415, B2 => 
                           n3494, ZN => n3417);
   U4970 : OAI22_X1 port map( A1 => n3418, A2 => n4053, B1 => n4051, B2 => 
                           n3417, ZN => n3419);
   U4971 : AOI211_X1 port map( C1 => n4056, C2 => n3628, A => n4055, B => n3419
                           , ZN => n3427);
   U4972 : AOI221_X1 port map( B1 => n3866, B2 => n3428, C1 => n3782, C2 => 
                           IF_ALUxN115, A => n4131, ZN => n3426);
   U4973 : AOI21_X1 port map( B1 => CtlToALU_port_alu_fun_0_port, B2 => n4056, 
                           A => IF_ALUxN115, ZN => n3420);
   U4974 : OAI22_X1 port map( A1 => n3420, A2 => n4123, B1 => n4117, B2 => 
                           n3624, ZN => n3425);
   U4975 : NAND2_X1 port map( A1 => n3490, A2 => n3591, ZN => n3422);
   U4976 : NAND2_X1 port map( A1 => n3422, A2 => n3491, ZN => n3629);
   U4977 : AOI22_X1 port map( A1 => n3490, A2 => n3421, B1 => n3592, B2 => 
                           n3726, ZN => n3627);
   U4978 : NAND2_X1 port map( A1 => n3954, A2 => n3627, ZN => n3423);
   U4979 : OAI21_X1 port map( B1 => n3954, B2 => n3629, A => n3423, ZN => n3559
                           );
   U4980 : OAI21_X1 port map( B1 => n3878, B2 => n3590, A => n3422, ZN => n3768
                           );
   U4981 : OAI21_X1 port map( B1 => n3954, B2 => n3768, A => n3423, ZN => n3547
                           );
   U4982 : OAI22_X1 port map( A1 => n3747, A2 => n3559, B1 => n3589, B2 => 
                           n3547, ZN => n3424);
   U4983 : NOR4_X1 port map( A1 => n3427, A2 => n3426, A3 => n3425, A4 => n3424
                           , ZN => n3431);
   U4984 : NOR3_X1 port map( A1 => n3428, A2 => n3866, A3 => n3816, ZN => n3429
                           );
   U4985 : AOI21_X1 port map( B1 => n3640, B2 => C596xDATA2_3, A => n3429, ZN 
                           => n3430);
   U4986 : OAI21_X1 port map( B1 => n3431, B2 => n4154, A => n3430, ZN => 
                           IF_ALUxN941);
   U4987 : NAND2_X1 port map( A1 => ALUtoCtl_port_2_port, A2 => n4415, ZN => 
                           n3433);
   U4988 : OAI211_X1 port map( C1 => n3735, C2 => n4112, A => n3433, B => n3432
                           , ZN => n6453);
   U4989 : NOR3_X1 port map( A1 => n3440, A2 => n3490, A3 => n3816, ZN => n3453
                           );
   U4990 : AOI22_X1 port map( A1 => n3490, A2 => n3435, B1 => n3434, B2 => 
                           n3726, ZN => n3804);
   U4991 : OAI221_X1 port map( B1 => n3860, B2 => n3489, C1 => n3494, C2 => 
                           n3495, A => n3490, ZN => n3437);
   U4992 : OAI21_X1 port map( B1 => n3490, B2 => n3436, A => n3437, ZN => n3439
                           );
   U4993 : INV_X1 port map( A => n3439, ZN => n3807);
   U4994 : AOI21_X1 port map( B1 => n3438, B2 => n3437, A => n3807, ZN => n3783
                           );
   U4995 : AOI22_X1 port map( A1 => n3954, A2 => n3804, B1 => n3783, B2 => 
                           n3782, ZN => n3511);
   U4996 : AOI22_X1 port map( A1 => n3954, A2 => n3804, B1 => n3439, B2 => 
                           n3782, ZN => n3520);
   U4997 : AOI22_X1 port map( A1 => n4063, A2 => n3511, B1 => n4062, B2 => 
                           n3520, ZN => n3451);
   U4998 : NAND2_X1 port map( A1 => n3440, A2 => n3726, ZN => n3959);
   U4999 : NAND2_X1 port map( A1 => n3490, A2 => IF_ALUxN114, ZN => n3956);
   U5000 : INV_X1 port map( A => n3441, ZN => n3784);
   U5001 : AOI22_X1 port map( A1 => n4127, A2 => n3726, B1 => n3761, B2 => 
                           n3784, ZN => n3442);
   U5002 : OAI221_X1 port map( B1 => n4131, B2 => n3959, C1 => n4131, C2 => 
                           n3956, A => n3442, ZN => n3449);
   U5003 : AOI22_X1 port map( A1 => n3490, A2 => n3444, B1 => n3443, B2 => 
                           n3726, ZN => n3805);
   U5004 : AOI22_X1 port map( A1 => n4045, A2 => IF_ALUxN114, B1 => IF_ALUxN115
                           , B2 => n3487, ZN => n4047);
   U5005 : AOI22_X1 port map( A1 => n3320, A2 => IF_ALUxN116, B1 => IF_ALUxN117
                           , B2 => n3487, ZN => n3482);
   U5006 : AOI22_X1 port map( A1 => n3725, A2 => n4047, B1 => n3482, B2 => 
                           n3494, ZN => n3445);
   U5007 : OAI22_X1 port map( A1 => n4053, A2 => n3446, B1 => n4051, B2 => 
                           n3445, ZN => n3447);
   U5008 : AOI211_X1 port map( C1 => n3805, C2 => n4056, A => n4055, B => n3447
                           , ZN => n3448);
   U5009 : AOI211_X1 port map( C1 => n4060, C2 => IF_ALUxN114, A => n3449, B =>
                           n3448, ZN => n3450);
   U5010 : AOI21_X1 port map( B1 => n3451, B2 => n3450, A => n4078, ZN => n3452
                           );
   U5011 : AOI211_X1 port map( C1 => n4152, C2 => C596xDATA2_2, A => n3453, B 
                           => n3452, ZN => n3454);
   U5012 : INV_X1 port map( A => n3454, ZN => IF_ALUxN940);
   U5013 : NAND2_X1 port map( A1 => ALUtoCtl_port_14_port, A2 => n4413, ZN => 
                           n3456);
   U5014 : OAI211_X1 port map( C1 => n3735, C2 => n4100, A => n3456, B => n3455
                           , ZN => n6455);
   U5015 : AOI221_X1 port map( B1 => n3458, B2 => n3866, C1 => n3457, C2 => 
                           n4056, A => n4055, ZN => n3468);
   U5016 : INV_X1 port map( A => n3942, ZN => n3469);
   U5017 : NAND2_X1 port map( A1 => n3469, A2 => IF_ALUxN126, ZN => n3459);
   U5018 : NAND2_X1 port map( A1 => n3941, A2 => n3942, ZN => n3945);
   U5019 : AOI21_X1 port map( B1 => n3459, B2 => n3945, A => n4131, ZN => n3467
                           );
   U5020 : AOI21_X1 port map( B1 => CtlToALU_port_alu_fun_0_port, B2 => n3942, 
                           A => IF_ALUxN126, ZN => n3462);
   U5021 : OAI22_X1 port map( A1 => n3462, A2 => n4123, B1 => n3461, B2 => 
                           n3460, ZN => n3466);
   U5022 : OAI22_X1 port map( A1 => n3464, A2 => n3747, B1 => n3862, B2 => 
                           n3463, ZN => n3465);
   U5023 : NOR4_X1 port map( A1 => n3468, A2 => n3467, A3 => n3466, A4 => n3465
                           , ZN => n3472);
   U5024 : NOR3_X1 port map( A1 => n3469, A2 => n3941, A3 => n3816, ZN => n3470
                           );
   U5025 : AOI21_X1 port map( B1 => n3640, B2 => C596xDATA2_14, A => n3470, ZN 
                           => n3471);
   U5026 : OAI21_X1 port map( B1 => n3472, B2 => n4154, A => n3471, ZN => 
                           IF_ALUxN952);
   U5027 : CLKBUF_X1 port map( A => n3735, Z => n3925);
   U5028 : NAND2_X1 port map( A1 => ALUtoCtl_port_4_port, A2 => n4415, ZN => 
                           n3474);
   U5029 : OAI211_X1 port map( C1 => n3925, C2 => n4110, A => n3474, B => n3473
                           , ZN => n6457);
   U5030 : AOI22_X1 port map( A1 => n4120, A2 => n3476, B1 => n3475, B2 => 
                           n3494, ZN => n3646);
   U5031 : AOI22_X1 port map( A1 => n4120, A2 => n3478, B1 => n3477, B2 => 
                           n3494, ZN => n3649);
   U5032 : AOI22_X1 port map( A1 => n3490, A2 => n3646, B1 => n3649, B2 => 
                           n3875, ZN => n3737);
   U5033 : AOI22_X1 port map( A1 => n4120, A2 => n3480, B1 => n3479, B2 => 
                           n4118, ZN => n3647);
   U5034 : AOI22_X1 port map( A1 => n4120, A2 => n3482, B1 => n3481, B2 => 
                           n3494, ZN => n4052);
   U5035 : OAI22_X1 port map( A1 => n4053, A2 => n3647, B1 => n4052, B2 => 
                           n4051, ZN => n3483);
   U5036 : AOI211_X1 port map( C1 => n3737, C2 => n4056, A => n4055, B => n3483
                           , ZN => n3502);
   U5037 : OAI22_X1 port map( A1 => n4118, A2 => n3485, B1 => n3484, B2 => 
                           n3860, ZN => n3652);
   U5038 : NAND3_X1 port map( A1 => n4045, A2 => n3860, A3 => IF_ALUxN112, ZN 
                           => n4066);
   U5039 : OAI22_X1 port map( A1 => n3875, A2 => n3652, B1 => n4066, B2 => 
                           n3490, ZN => n3745);
   U5040 : INV_X1 port map( A => n3745, ZN => n3712);
   U5041 : OAI22_X1 port map( A1 => n3953, A2 => n4079, B1 => n3712, B2 => 
                           n3671, ZN => n3501);
   U5042 : NOR2_X1 port map( A1 => n3953, A2 => IF_ALUxN116, ZN => n3961);
   U5043 : AOI21_X1 port map( B1 => n3953, B2 => IF_ALUxN116, A => n3961, ZN =>
                           n3486);
   U5044 : OAI22_X1 port map( A1 => n3503, A2 => n4123, B1 => n3486, B2 => 
                           n4131, ZN => n3500);
   U5045 : OAI221_X1 port map( B1 => n3320, B2 => n4144, C1 => n3487, C2 => 
                           IF_ALUxN142, A => n4118, ZN => n3488);
   U5046 : OAI21_X1 port map( B1 => n4118, B2 => n3489, A => n3488, ZN => n3855
                           );
   U5047 : NAND2_X1 port map( A1 => n3490, A2 => n3855, ZN => n3497);
   U5048 : NAND2_X1 port map( A1 => n3491, A2 => n3497, ZN => n3744);
   U5049 : AOI22_X1 port map( A1 => n4120, A2 => n3493, B1 => n3492, B2 => 
                           n3494, ZN => n3648);
   U5050 : AOI22_X1 port map( A1 => n4120, A2 => n3496, B1 => n3495, B2 => 
                           n3494, ZN => n3645);
   U5051 : AOI22_X1 port map( A1 => n3878, A2 => n3648, B1 => n3645, B2 => 
                           n3875, ZN => n3736);
   U5052 : NOR2_X1 port map( A1 => n3736, A2 => n3782, ZN => n3498);
   U5053 : AOI21_X1 port map( B1 => n3782, B2 => n3744, A => n3498, ZN => n3715
                           );
   U5054 : INV_X1 port map( A => n3497, ZN => n3738);
   U5055 : AOI21_X1 port map( B1 => n3738, B2 => n4056, A => n3498, ZN => n3714
                           );
   U5056 : OAI22_X1 port map( A1 => n3715, A2 => n3747, B1 => n3714, B2 => 
                           n3589, ZN => n3499);
   U5057 : NOR4_X1 port map( A1 => n3502, A2 => n3501, A3 => n3500, A4 => n3499
                           , ZN => n3506);
   U5058 : NOR3_X1 port map( A1 => n3953, A2 => n3503, A3 => n4148, ZN => n3504
                           );
   U5059 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_4, A => n3504, ZN 
                           => n3505);
   U5060 : OAI21_X1 port map( B1 => n3506, B2 => n4154, A => n3505, ZN => 
                           IF_ALUxN942);
   U5061 : NAND2_X1 port map( A1 => ALUtoCtl_port_18_port, A2 => n4415, ZN => 
                           n3508);
   U5062 : OAI211_X1 port map( C1 => n3735, C2 => n4096, A => n3508, B => n3507
                           , ZN => n6459);
   U5063 : INV_X1 port map( A => n3996, ZN => n3514);
   U5064 : NOR3_X1 port map( A1 => n3997, A2 => n3514, A3 => n3816, ZN => n3524
                           );
   U5065 : AOI22_X1 port map( A1 => n3878, A2 => n3510, B1 => n3509, B2 => 
                           n3875, ZN => n3786);
   U5066 : AOI22_X1 port map( A1 => n3891, A2 => n3511, B1 => n3912, B2 => 
                           n3786, ZN => n3522);
   U5067 : AOI22_X1 port map( A1 => n4060, A2 => IF_ALUxN130, B1 => n4127, B2 
                           => n3996, ZN => n3518);
   U5068 : AOI22_X1 port map( A1 => n3878, A2 => n3513, B1 => n3512, B2 => 
                           n3726, ZN => n3787);
   U5069 : NOR2_X1 port map( A1 => n4056, A2 => n3894, ZN => n3689);
   U5070 : INV_X1 port map( A => n3689, ZN => n3711);
   U5071 : NOR2_X1 port map( A1 => n3726, A2 => n3711, ZN => n3909);
   U5072 : AOI22_X1 port map( A1 => n3914, A2 => n3787, B1 => n3909, B2 => 
                           n3784, ZN => n3517);
   U5073 : NOR2_X1 port map( A1 => n3997, A2 => n3996, ZN => n3515);
   U5074 : NOR2_X1 port map( A1 => n3514, A2 => IF_ALUxN130, ZN => n4006);
   U5075 : OAI21_X1 port map( B1 => n3515, B2 => n4006, A => n4073, ZN => n3516
                           );
   U5076 : NAND4_X1 port map( A1 => n3518, A2 => n3517, A3 => n3882, A4 => 
                           n3516, ZN => n3519);
   U5077 : AOI21_X1 port map( B1 => n3696, B2 => n3520, A => n3519, ZN => n3521
                           );
   U5078 : AOI21_X1 port map( B1 => n3522, B2 => n3521, A => n4078, ZN => n3523
                           );
   U5079 : AOI211_X1 port map( C1 => n4152, C2 => C596xDATA2_18, A => n3524, B 
                           => n3523, ZN => n3525);
   U5080 : INV_X1 port map( A => n3525, ZN => IF_ALUxN956);
   U5081 : NAND2_X1 port map( A1 => ALUtoCtl_port_21_port, A2 => n4415, ZN => 
                           n3527);
   U5082 : OAI211_X1 port map( C1 => n3735, C2 => n4093, A => n3527, B => n3526
                           , ZN => n6461);
   U5083 : AOI22_X1 port map( A1 => n3878, A2 => n3529, B1 => n3528, B2 => 
                           n3726, ZN => n3605);
   U5084 : INV_X1 port map( A => n3912, ZN => n4137);
   U5085 : OAI22_X1 port map( A1 => n3605, A2 => n4137, B1 => n3604, B2 => 
                           n3711, ZN => n3539);
   U5086 : AOI22_X1 port map( A1 => n3878, A2 => n3531, B1 => n3530, B2 => 
                           n3875, ZN => n3827);
   U5087 : AOI22_X1 port map( A1 => n4060, A2 => IF_ALUxN133, B1 => n4127, B2 
                           => n3532, ZN => n3534);
   U5088 : NOR2_X1 port map( A1 => n3540, A2 => n3532, ZN => n4015);
   U5089 : INV_X1 port map( A => n3532, ZN => n3541);
   U5090 : NOR2_X1 port map( A1 => n3541, A2 => IF_ALUxN133, ZN => n3940);
   U5091 : OAI21_X1 port map( B1 => n4015, B2 => n3940, A => n4073, ZN => n3533
                           );
   U5092 : OAI211_X1 port map( C1 => n3827, C2 => n3671, A => n3534, B => n3533
                           , ZN => n3538);
   U5093 : OAI22_X1 port map( A1 => n3536, A2 => n3851, B1 => n3535, B2 => 
                           n3713, ZN => n3537);
   U5094 : NOR4_X1 port map( A1 => n3908, A2 => n3539, A3 => n3538, A4 => n3537
                           , ZN => n3544);
   U5095 : NOR3_X1 port map( A1 => n3541, A2 => n3540, A3 => n4148, ZN => n3542
                           );
   U5096 : AOI21_X1 port map( B1 => n3640, B2 => C596xDATA2_21, A => n3542, ZN 
                           => n3543);
   U5097 : OAI21_X1 port map( B1 => n3544, B2 => n4078, A => n3543, ZN => 
                           IF_ALUxN959);
   U5098 : NAND2_X1 port map( A1 => ALUtoCtl_port_19_port, A2 => n4415, ZN => 
                           n3546);
   U5099 : OAI211_X1 port map( C1 => n3735, C2 => n4095, A => n3546, B => n3545
                           , ZN => n6463);
   U5100 : INV_X1 port map( A => n3547, ZN => n3562);
   U5101 : AOI22_X1 port map( A1 => n3860, A2 => n3549, B1 => n3548, B2 => 
                           n3856, ZN => n3668);
   U5102 : AOI22_X1 port map( A1 => n3725, A2 => n3551, B1 => n3550, B2 => 
                           n3494, ZN => n3587);
   U5103 : AOI22_X1 port map( A1 => n3878, A2 => n3668, B1 => n3587, B2 => 
                           n3726, ZN => n3767);
   U5104 : INV_X1 port map( A => n4007, ZN => n3994);
   U5105 : OAI22_X1 port map( A1 => n4008, A2 => n4123, B1 => n3994, B2 => 
                           n4079, ZN => n3552);
   U5106 : AOI211_X1 port map( C1 => n3553, C2 => n3909, A => n3908, B => n3552
                           , ZN => n3555);
   U5107 : OAI221_X1 port map( B1 => n4008, B2 => n3994, C1 => IF_ALUxN131, C2 
                           => n4007, A => n4073, ZN => n3554);
   U5108 : OAI211_X1 port map( C1 => n3767, C2 => n3671, A => n3555, B => n3554
                           , ZN => n3561);
   U5109 : AOI22_X1 port map( A1 => n3860, A2 => n3557, B1 => n3556, B2 => 
                           n3856, ZN => n3586);
   U5110 : AOI22_X1 port map( A1 => n3878, A2 => n3586, B1 => n3558, B2 => 
                           n3875, ZN => n3626);
   U5111 : OAI22_X1 port map( A1 => n3626, A2 => n4137, B1 => n3851, B2 => 
                           n3559, ZN => n3560);
   U5112 : AOI211_X1 port map( C1 => n3696, C2 => n3562, A => n3561, B => n3560
                           , ZN => n3565);
   U5113 : NOR3_X1 port map( A1 => n3994, A2 => n4008, A3 => n3816, ZN => n3563
                           );
   U5114 : AOI21_X1 port map( B1 => n3640, B2 => C596xDATA2_19, A => n3563, ZN 
                           => n3564);
   U5115 : OAI21_X1 port map( B1 => n3565, B2 => n4078, A => n3564, ZN => 
                           IF_ALUxN957);
   U5116 : NAND2_X1 port map( A1 => ALUtoCtl_port_17_port, A2 => n4415, ZN => 
                           n3567);
   U5117 : OAI211_X1 port map( C1 => n3735, C2 => n4097, A => n3567, B => n3566
                           , ZN => n6465);
   U5118 : INV_X1 port map( A => n3568, ZN => n3579);
   U5119 : NAND2_X1 port map( A1 => n4002, A2 => n4001, ZN => n3569);
   U5120 : INV_X1 port map( A => n4001, ZN => n3580);
   U5121 : NAND2_X1 port map( A1 => n3580, A2 => IF_ALUxN129, ZN => n3995);
   U5122 : AOI21_X1 port map( B1 => n3569, B2 => n3995, A => n4131, ZN => n3570
                           );
   U5123 : AOI211_X1 port map( C1 => n3571, C2 => n3909, A => n3908, B => n3570
                           , ZN => n3573);
   U5124 : OAI221_X1 port map( B1 => IF_ALUxN129, B2 => 
                           CtlToALU_port_alu_fun_0_port, C1 => IF_ALUxN129, C2 
                           => n4001, A => n4060, ZN => n3572);
   U5125 : OAI211_X1 port map( C1 => n3574, C2 => n3671, A => n3573, B => n3572
                           , ZN => n3578);
   U5126 : OAI22_X1 port map( A1 => n3576, A2 => n4137, B1 => n3851, B2 => 
                           n3575, ZN => n3577);
   U5127 : AOI211_X1 port map( C1 => n3696, C2 => n3579, A => n3578, B => n3577
                           , ZN => n3583);
   U5128 : NOR3_X1 port map( A1 => n3580, A2 => n4002, A3 => n3816, ZN => n3581
                           );
   U5129 : AOI21_X1 port map( B1 => n3640, B2 => C596xDATA2_17, A => n3581, ZN 
                           => n3582);
   U5130 : OAI21_X1 port map( B1 => n3583, B2 => n4078, A => n3582, ZN => 
                           IF_ALUxN955);
   U5131 : NAND2_X1 port map( A1 => ALUtoCtl_port_15_port, A2 => n4415, ZN => 
                           n3585);
   U5132 : OAI211_X1 port map( C1 => n3735, C2 => n4099, A => n3585, B => n3584
                           , ZN => n6467);
   U5133 : INV_X1 port map( A => n3944, ZN => n3948);
   U5134 : NOR3_X1 port map( A1 => n3948, A2 => n3943, A3 => n3816, ZN => n3600
                           );
   U5135 : AOI22_X1 port map( A1 => n3878, A2 => n3587, B1 => n3586, B2 => 
                           n3875, ZN => n3665);
   U5136 : AOI22_X1 port map( A1 => n3866, A2 => n3665, B1 => n3664, B2 => 
                           n3782, ZN => n4134);
   U5137 : OAI22_X1 port map( A1 => n3943, A2 => n4123, B1 => n3948, B2 => 
                           n4079, ZN => n3588);
   U5138 : AOI211_X1 port map( C1 => n4134, C2 => n3636, A => n3908, B => n3588
                           , ZN => n3598);
   U5139 : NOR2_X1 port map( A1 => n3589, A2 => n4051, ZN => n3609);
   U5140 : INV_X1 port map( A => n3590, ZN => n4126);
   U5141 : AOI22_X1 port map( A1 => n3878, A2 => n3592, B1 => n3591, B2 => 
                           n3726, ZN => n3593);
   U5142 : AOI221_X1 port map( B1 => n3954, B2 => n3594, C1 => n3782, C2 => 
                           n3593, A => n4055, ZN => n3596);
   U5143 : AOI221_X1 port map( B1 => n3943, B2 => n3948, C1 => IF_ALUxN127, C2 
                           => n3944, A => n4131, ZN => n3595);
   U5144 : AOI211_X1 port map( C1 => n3609, C2 => n4126, A => n3596, B => n3595
                           , ZN => n3597);
   U5145 : AOI21_X1 port map( B1 => n3598, B2 => n3597, A => n4078, ZN => n3599
                           );
   U5146 : AOI211_X1 port map( C1 => n4152, C2 => C596xDATA2_15, A => n3600, B 
                           => n3599, ZN => n3601);
   U5147 : INV_X1 port map( A => n3601, ZN => IF_ALUxN953);
   U5148 : NAND2_X1 port map( A1 => ALUtoCtl_port_13_port, A2 => n4415, ZN => 
                           n3603);
   U5149 : OAI211_X1 port map( C1 => n3925, C2 => n4101, A => n3603, B => n3602
                           , ZN => n6469);
   U5150 : AOI22_X1 port map( A1 => n3954, A2 => n3605, B1 => n3604, B2 => 
                           n3782, ZN => n3838);
   U5151 : AOI221_X1 port map( B1 => n3607, B2 => n3782, C1 => n3606, C2 => 
                           n3866, A => n4055, ZN => n3616);
   U5152 : AOI21_X1 port map( B1 => n3954, B2 => n3608, A => n3743, ZN => n3835
                           );
   U5153 : AOI22_X1 port map( A1 => n4127, A2 => n3610, B1 => n3609, B2 => 
                           n3832, ZN => n3614);
   U5154 : NOR2_X1 port map( A1 => n3617, A2 => n3610, ZN => n3980);
   U5155 : INV_X1 port map( A => n3980, ZN => n3611);
   U5156 : NAND2_X1 port map( A1 => n3617, A2 => n3610, ZN => n3946);
   U5157 : AOI21_X1 port map( B1 => n3611, B2 => n3946, A => n4131, ZN => n3612
                           );
   U5158 : AOI21_X1 port map( B1 => n4060, B2 => IF_ALUxN125, A => n3612, ZN =>
                           n3613);
   U5159 : OAI211_X1 port map( C1 => n3835, C2 => n3747, A => n3614, B => n3613
                           , ZN => n3615);
   U5160 : AOI211_X1 port map( C1 => n3838, C2 => n3636, A => n3616, B => n3615
                           , ZN => n3621);
   U5161 : NOR3_X1 port map( A1 => n3618, A2 => n4148, A3 => n3617, ZN => n3619
                           );
   U5162 : AOI21_X1 port map( B1 => n3640, B2 => C596xDATA2_13, A => n3619, ZN 
                           => n3620);
   U5163 : OAI21_X1 port map( B1 => n3621, B2 => n4078, A => n3620, ZN => 
                           IF_ALUxN951);
   U5164 : NAND2_X1 port map( A1 => ALUtoCtl_port_11_port, A2 => n4415, ZN => 
                           n3623);
   U5165 : OAI211_X1 port map( C1 => n3735, C2 => n4103, A => n3623, B => n3622
                           , ZN => n6471);
   U5166 : OAI22_X1 port map( A1 => n3626, A2 => n3782, B1 => n3625, B2 => 
                           n3624, ZN => n3774);
   U5167 : AOI221_X1 port map( B1 => n3866, B2 => n3628, C1 => n3782, C2 => 
                           n3627, A => n4055, ZN => n3635);
   U5168 : AOI21_X1 port map( B1 => n3954, B2 => n3629, A => n3743, ZN => n3771
                           );
   U5169 : INV_X1 port map( A => n3631, ZN => n3637);
   U5170 : OAI21_X1 port map( B1 => n3637, B2 => n6201, A => n3638, ZN => n3630
                           );
   U5171 : AOI22_X1 port map( A1 => n4060, A2 => n3630, B1 => n3806, B2 => 
                           n3768, ZN => n3633);
   U5172 : NOR2_X1 port map( A1 => n3637, A2 => IF_ALUxN123, ZN => n3993);
   U5173 : NOR2_X1 port map( A1 => n3638, A2 => n3631, ZN => n3978);
   U5174 : OAI21_X1 port map( B1 => n3993, B2 => n3978, A => n4073, ZN => n3632
                           );
   U5175 : OAI211_X1 port map( C1 => n3771, C2 => n3747, A => n3633, B => n3632
                           , ZN => n3634);
   U5176 : AOI211_X1 port map( C1 => n3636, C2 => n3774, A => n3635, B => n3634
                           , ZN => n3642);
   U5177 : NOR3_X1 port map( A1 => n3638, A2 => n3637, A3 => n3816, ZN => n3639
                           );
   U5178 : AOI21_X1 port map( B1 => n3640, B2 => C596xDATA2_11, A => n3639, ZN 
                           => n3641);
   U5179 : OAI21_X1 port map( B1 => n3642, B2 => n4078, A => n3641, ZN => 
                           IF_ALUxN949);
   U5180 : NAND2_X1 port map( A1 => ALUtoCtl_port_8_port, A2 => n4415, ZN => 
                           n3644);
   U5181 : OAI211_X1 port map( C1 => n3925, C2 => n4106, A => n3644, B => n3643
                           , ZN => n6473);
   U5182 : AOI22_X1 port map( A1 => n3878, A2 => n3645, B1 => n3855, B2 => 
                           n3726, ZN => n3903);
   U5183 : OAI21_X1 port map( B1 => n3903, B2 => n3782, A => n3781, ZN => n3890
                           );
   U5184 : AOI22_X1 port map( A1 => n3878, A2 => n3647, B1 => n3646, B2 => 
                           n3726, ZN => n4057);
   U5185 : AOI22_X1 port map( A1 => n3878, A2 => n3649, B1 => n3648, B2 => 
                           n3726, ZN => n3904);
   U5186 : AOI221_X1 port map( B1 => n4057, B2 => n3866, C1 => n3904, C2 => 
                           n4056, A => n4055, ZN => n3657);
   U5187 : AOI22_X1 port map( A1 => n3860, A2 => n3651, B1 => n3650, B2 => 
                           n3856, ZN => n3727);
   U5188 : AOI22_X1 port map( A1 => n3490, A2 => n3727, B1 => n3652, B2 => 
                           n3726, ZN => n3911);
   U5189 : INV_X1 port map( A => n4066, ZN => n3910);
   U5190 : AOI22_X1 port map( A1 => n3954, A2 => n3911, B1 => n3910, B2 => 
                           n3785, ZN => n3895);
   U5191 : INV_X1 port map( A => n3903, ZN => n3879);
   U5192 : AOI22_X1 port map( A1 => n4060, A2 => IF_ALUxN120, B1 => n3806, B2 
                           => n3879, ZN => n3655);
   U5193 : INV_X1 port map( A => n3951, ZN => n3658);
   U5194 : NAND2_X1 port map( A1 => n3658, A2 => IF_ALUxN120, ZN => n3973);
   U5195 : OAI21_X1 port map( B1 => n3658, B2 => IF_ALUxN120, A => n3973, ZN =>
                           n3653);
   U5196 : AOI22_X1 port map( A1 => n4127, A2 => n3951, B1 => n4073, B2 => 
                           n3653, ZN => n3654);
   U5197 : OAI211_X1 port map( C1 => n3895, C2 => n3862, A => n3655, B => n3654
                           , ZN => n3656);
   U5198 : AOI211_X1 port map( C1 => n4063, C2 => n3890, A => n3657, B => n3656
                           , ZN => n3661);
   U5199 : NOR3_X1 port map( A1 => n3952, A2 => n3658, A3 => n3816, ZN => n3659
                           );
   U5200 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_8, A => n3659, ZN 
                           => n3660);
   U5201 : OAI21_X1 port map( B1 => n3661, B2 => n4078, A => n3660, ZN => 
                           IF_ALUxN946);
   U5202 : NAND2_X1 port map( A1 => ALUtoCtl_port_23_port, A2 => n4413, ZN => 
                           n3663);
   U5203 : OAI211_X1 port map( C1 => n3735, C2 => n4091, A => n3663, B => n3662
                           , ZN => n6475);
   U5204 : OAI22_X1 port map( A1 => n3665, A2 => n4137, B1 => n3664, B2 => 
                           n3711, ZN => n3677);
   U5205 : NOR2_X1 port map( A1 => n3679, A2 => n3669, ZN => n3935);
   U5206 : NAND2_X1 port map( A1 => n3679, A2 => n3669, ZN => n3937);
   U5207 : INV_X1 port map( A => n3937, ZN => n3673);
   U5208 : AOI22_X1 port map( A1 => n3860, A2 => n3667, B1 => n3666, B2 => 
                           n3856, ZN => n3760);
   U5209 : AOI22_X1 port map( A1 => n3878, A2 => n3760, B1 => n3668, B2 => 
                           n3875, ZN => n4138);
   U5210 : AOI21_X1 port map( B1 => CtlToALU_port_alu_fun_0_port, B2 => n3669, 
                           A => IF_ALUxN135, ZN => n3670);
   U5211 : OAI22_X1 port map( A1 => n4138, A2 => n3671, B1 => n3670, B2 => 
                           n4123, ZN => n3672);
   U5212 : AOI221_X1 port map( B1 => n3935, B2 => n4073, C1 => n3673, C2 => 
                           n4073, A => n3672, ZN => n3674);
   U5213 : OAI211_X1 port map( C1 => n3675, C2 => n3713, A => n3674, B => n3882
                           , ZN => n3676);
   U5214 : AOI211_X1 port map( C1 => n3891, C2 => n3678, A => n3677, B => n3676
                           , ZN => n3683);
   U5215 : NOR3_X1 port map( A1 => n3680, A2 => n3816, A3 => n3679, ZN => n3681
                           );
   U5216 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_23, A => n3681, ZN 
                           => n3682);
   U5217 : OAI21_X1 port map( B1 => n3683, B2 => n4078, A => n3682, ZN => 
                           IF_ALUxN961);
   U5218 : NAND2_X1 port map( A1 => ALUtoCtl_port_22_port, A2 => n4413, ZN => 
                           n3685);
   U5219 : OAI211_X1 port map( C1 => n3735, C2 => n4092, A => n3685, B => n3684
                           , ZN => n6477);
   U5220 : AOI22_X1 port map( A1 => n3914, A2 => n3687, B1 => n3912, B2 => 
                           n3686, ZN => n3698);
   U5221 : NAND2_X1 port map( A1 => n3701, A2 => n3688, ZN => n3936);
   U5222 : INV_X1 port map( A => n3688, ZN => n3934);
   U5223 : NAND2_X1 port map( A1 => n3934, A2 => IF_ALUxN134, ZN => n3693);
   U5224 : OAI21_X1 port map( B1 => n3934, B2 => n6201, A => n3701, ZN => n3691
                           );
   U5225 : AOI22_X1 port map( A1 => n4060, A2 => n3691, B1 => n3690, B2 => 
                           n3689, ZN => n3692);
   U5226 : OAI221_X1 port map( B1 => n4131, B2 => n3936, C1 => n4131, C2 => 
                           n3693, A => n3692, ZN => n3694);
   U5227 : AOI211_X1 port map( C1 => n3696, C2 => n3695, A => n3908, B => n3694
                           , ZN => n3697);
   U5228 : OAI211_X1 port map( C1 => n3699, C2 => n3851, A => n3698, B => n3697
                           , ZN => n3700);
   U5229 : INV_X1 port map( A => n3700, ZN => n3704);
   U5230 : NOR3_X1 port map( A1 => n3934, A2 => n3701, A3 => n3816, ZN => n3702
                           );
   U5231 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_22, A => n3702, ZN 
                           => n3703);
   U5232 : OAI21_X1 port map( B1 => n4078, B2 => n3704, A => n3703, ZN => 
                           IF_ALUxN960);
   U5233 : NAND2_X1 port map( A1 => ALUtoCtl_port_20_port, A2 => n4413, ZN => 
                           n3706);
   U5234 : OAI211_X1 port map( C1 => n3735, C2 => n4094, A => n3706, B => n3705
                           , ZN => n6479);
   U5235 : INV_X1 port map( A => n3709, ZN => n4016);
   U5236 : NOR3_X1 port map( A1 => n3707, A2 => n4016, A3 => n3816, ZN => n3731
                           );
   U5237 : NAND2_X1 port map( A1 => n3707, A2 => n3709, ZN => n4009);
   U5238 : NAND2_X1 port map( A1 => n4016, A2 => IF_ALUxN132, ZN => n3708);
   U5239 : AOI21_X1 port map( B1 => n4009, B2 => n3708, A => n4131, ZN => n3718
                           );
   U5240 : AOI21_X1 port map( B1 => CtlToALU_port_alu_fun_0_port, B2 => n3709, 
                           A => IF_ALUxN132, ZN => n3710);
   U5241 : OAI22_X1 port map( A1 => n3712, A2 => n3711, B1 => n3710, B2 => 
                           n4123, ZN => n3717);
   U5242 : OAI22_X1 port map( A1 => n3715, A2 => n3851, B1 => n3714, B2 => 
                           n3713, ZN => n3716);
   U5243 : NOR4_X1 port map( A1 => n3908, A2 => n3718, A3 => n3717, A4 => n3716
                           , ZN => n3729);
   U5244 : AOI22_X1 port map( A1 => n4120, A2 => n3720, B1 => n3719, B2 => 
                           n3856, ZN => n3887);
   U5245 : AOI22_X1 port map( A1 => n4120, A2 => n3722, B1 => n3721, B2 => 
                           n3856, ZN => n3877);
   U5246 : AOI22_X1 port map( A1 => n3878, A2 => n3887, B1 => n3877, B2 => 
                           n3726, ZN => n3867);
   U5247 : AOI22_X1 port map( A1 => n3725, A2 => n3724, B1 => n3723, B2 => 
                           n3856, ZN => n3876);
   U5248 : AOI22_X1 port map( A1 => n3878, A2 => n3876, B1 => n3727, B2 => 
                           n3726, ZN => n3746);
   U5249 : AOI22_X1 port map( A1 => n3914, A2 => n3867, B1 => n3912, B2 => 
                           n3746, ZN => n3728);
   U5250 : AOI21_X1 port map( B1 => n3729, B2 => n3728, A => n4078, ZN => n3730
                           );
   U5251 : AOI211_X1 port map( C1 => n4152, C2 => C596xDATA2_20, A => n3731, B 
                           => n3730, ZN => n3732);
   U5252 : INV_X1 port map( A => n3732, ZN => IF_ALUxN958);
   U5253 : NAND2_X1 port map( A1 => ALUtoCtl_port_12_port, A2 => n4413, ZN => 
                           n3734);
   U5254 : OAI211_X1 port map( C1 => n3735, C2 => n4102, A => n3734, B => n3733
                           , ZN => n6481);
   U5255 : AOI221_X1 port map( B1 => n3737, B2 => n3866, C1 => n3736, C2 => 
                           n4056, A => n4055, ZN => n3750);
   U5256 : AOI22_X1 port map( A1 => n4127, A2 => n3739, B1 => n3806, B2 => 
                           n3738, ZN => n3742);
   U5257 : NOR2_X1 port map( A1 => n3751, A2 => n3739, ZN => n3979);
   U5258 : NAND2_X1 port map( A1 => n3751, A2 => n3739, ZN => n3947);
   U5259 : INV_X1 port map( A => n3947, ZN => n3740);
   U5260 : OAI21_X1 port map( B1 => n3979, B2 => n3740, A => n4073, ZN => n3741
                           );
   U5261 : OAI211_X1 port map( C1 => n3751, C2 => n4123, A => n3742, B => n3741
                           , ZN => n3749);
   U5262 : AOI21_X1 port map( B1 => n3866, B2 => n3744, A => n3743, ZN => n3852
                           );
   U5263 : AOI22_X1 port map( A1 => n3954, A2 => n3746, B1 => n3745, B2 => 
                           n3782, ZN => n3850);
   U5264 : OAI22_X1 port map( A1 => n3852, A2 => n3747, B1 => n3850, B2 => 
                           n3862, ZN => n3748);
   U5265 : NOR3_X1 port map( A1 => n3750, A2 => n3749, A3 => n3748, ZN => n3755
                           );
   U5266 : NOR3_X1 port map( A1 => n3752, A2 => n3816, A3 => n3751, ZN => n3753
                           );
   U5267 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_12, A => n3753, ZN 
                           => n3754);
   U5268 : OAI21_X1 port map( B1 => n3755, B2 => n4078, A => n3754, ZN => 
                           IF_ALUxN950);
   U5269 : NAND2_X1 port map( A1 => ALUtoCtl_port_27_port, A2 => n4413, ZN => 
                           n3757);
   U5270 : OAI211_X1 port map( C1 => n3925, C2 => n4087, A => n3757, B => n3756
                           , ZN => n6483);
   U5271 : AOI22_X1 port map( A1 => n4060, A2 => IF_ALUxN139, B1 => n4127, B2 
                           => n3762, ZN => n3766);
   U5272 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN139, B1 => IF_ALUxN138
                           , B2 => n4116, ZN => n3823);
   U5273 : AOI22_X1 port map( A1 => n4120, A2 => n3823, B1 => n3759, B2 => 
                           n4118, ZN => n4142);
   U5274 : AOI22_X1 port map( A1 => n3761, A2 => n4142, B1 => n3760, B2 => 
                           n4141, ZN => n3765);
   U5275 : INV_X1 port map( A => n3762, ZN => n4029);
   U5276 : NOR2_X1 port map( A1 => n4029, A2 => IF_ALUxN139, ZN => n4031);
   U5277 : NOR2_X1 port map( A1 => n3775, A2 => n3762, ZN => n3763);
   U5278 : OAI21_X1 port map( B1 => n4031, B2 => n3763, A => n4073, ZN => n3764
                           );
   U5279 : NAND4_X1 port map( A1 => n3766, A2 => n3765, A3 => n3882, A4 => 
                           n3764, ZN => n3773);
   U5280 : INV_X1 port map( A => n3767, ZN => n3769);
   U5281 : AOI22_X1 port map( A1 => n3912, A2 => n3769, B1 => n3880, B2 => 
                           n3768, ZN => n3770);
   U5282 : OAI21_X1 port map( B1 => n3771, B2 => n3851, A => n3770, ZN => n3772
                           );
   U5283 : AOI211_X1 port map( C1 => n4135, C2 => n3774, A => n3773, B => n3772
                           , ZN => n3778);
   U5284 : NOR3_X1 port map( A1 => n4029, A2 => n3775, A3 => n3816, ZN => n3776
                           );
   U5285 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_27, A => n3776, ZN 
                           => n3777);
   U5286 : OAI21_X1 port map( B1 => n3778, B2 => n4078, A => n3777, ZN => 
                           IF_ALUxN965);
   U5287 : NAND2_X1 port map( A1 => ALUtoCtl_port_26_port, A2 => n4413, ZN => 
                           n3780);
   U5288 : OAI211_X1 port map( C1 => n3925, C2 => n4088, A => n3780, B => n3779
                           , ZN => n6485);
   U5289 : OAI21_X1 port map( B1 => n3783, B2 => n3782, A => n3781, ZN => n3815
                           );
   U5290 : AOI22_X1 port map( A1 => n3954, A2 => n3786, B1 => n3785, B2 => 
                           n3784, ZN => n3812);
   U5291 : AOI22_X1 port map( A1 => n3807, A2 => n3880, B1 => n3912, B2 => 
                           n3787, ZN => n3795);
   U5292 : NAND2_X1 port map( A1 => n3798, A2 => n3788, ZN => n4028);
   U5293 : INV_X1 port map( A => n3788, ZN => n3797);
   U5294 : NAND2_X1 port map( A1 => n3797, A2 => IF_ALUxN138, ZN => n4024);
   U5295 : AOI21_X1 port map( B1 => n4028, B2 => n4024, A => n4131, ZN => n3793
                           );
   U5296 : OAI22_X1 port map( A1 => n3798, A2 => n4123, B1 => n3797, B2 => 
                           n4079, ZN => n3792);
   U5297 : OAI22_X1 port map( A1 => n3790, A2 => n3886, B1 => n3789, B2 => 
                           n4117, ZN => n3791);
   U5298 : NOR4_X1 port map( A1 => n3908, A2 => n3793, A3 => n3792, A4 => n3791
                           , ZN => n3794);
   U5299 : OAI211_X1 port map( C1 => n3812, C2 => n3894, A => n3795, B => n3794
                           , ZN => n3796);
   U5300 : AOI21_X1 port map( B1 => n3891, B2 => n3815, A => n3796, ZN => n3801
                           );
   U5301 : NOR3_X1 port map( A1 => n3798, A2 => n3797, A3 => n3816, ZN => n3799
                           );
   U5302 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_26, A => n3799, ZN 
                           => n3800);
   U5303 : OAI21_X1 port map( B1 => n3801, B2 => n4078, A => n3800, ZN => 
                           IF_ALUxN964);
   U5304 : NAND2_X1 port map( A1 => ALUtoCtl_port_10_port, A2 => n4413, ZN => 
                           n3803);
   U5305 : OAI211_X1 port map( C1 => n3925, C2 => n4104, A => n3803, B => n3802
                           , ZN => n6487);
   U5306 : AOI221_X1 port map( B1 => n3805, B2 => n3866, C1 => n3804, C2 => 
                           n4056, A => n4055, ZN => n3814);
   U5307 : INV_X1 port map( A => n3982, ZN => n3817);
   U5308 : OAI21_X1 port map( B1 => n3817, B2 => n6201, A => n3983, ZN => n3808
                           );
   U5309 : AOI22_X1 port map( A1 => n4060, A2 => n3808, B1 => n3807, B2 => 
                           n3806, ZN => n3811);
   U5310 : NOR2_X1 port map( A1 => n3817, A2 => IF_ALUxN122, ZN => n3992);
   U5311 : NOR2_X1 port map( A1 => n3983, A2 => n3982, ZN => n3809);
   U5312 : OAI21_X1 port map( B1 => n3992, B2 => n3809, A => n4073, ZN => n3810
                           );
   U5313 : OAI211_X1 port map( C1 => n3812, C2 => n3862, A => n3811, B => n3810
                           , ZN => n3813);
   U5314 : AOI211_X1 port map( C1 => n4063, C2 => n3815, A => n3814, B => n3813
                           , ZN => n3820);
   U5315 : NOR3_X1 port map( A1 => n3983, A2 => n3817, A3 => n3816, ZN => n3818
                           );
   U5316 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_10, A => n3818, ZN 
                           => n3819);
   U5317 : OAI21_X1 port map( B1 => n3820, B2 => n4154, A => n3819, ZN => 
                           IF_ALUxN948);
   U5318 : NAND2_X1 port map( A1 => ALUtoCtl_port_29_port, A2 => n4413, ZN => 
                           n3822);
   U5319 : OAI211_X1 port map( C1 => n3925, C2 => n4085, A => n3822, B => n3821
                           , ZN => n6489);
   U5320 : AOI22_X1 port map( A1 => n3758, A2 => IF_ALUxN141, B1 => IF_ALUxN140
                           , B2 => n4116, ZN => n4119);
   U5321 : AOI22_X1 port map( A1 => n4120, A2 => n4119, B1 => n3823, B2 => 
                           n4118, ZN => n3824);
   U5322 : OAI22_X1 port map( A1 => n3825, A2 => n4053, B1 => n4051, B2 => 
                           n3824, ZN => n3826);
   U5323 : AOI211_X1 port map( C1 => n3827, C2 => n4056, A => n3862, B => n3826
                           , ZN => n3837);
   U5324 : AOI22_X1 port map( A1 => n4060, A2 => IF_ALUxN141, B1 => n4127, B2 
                           => n3829, ZN => n3834);
   U5325 : INV_X1 port map( A => n3828, ZN => n4125);
   U5326 : NOR2_X1 port map( A1 => n3839, A2 => n3829, ZN => n4034);
   U5327 : INV_X1 port map( A => n4034, ZN => n3830);
   U5328 : NAND2_X1 port map( A1 => n3839, A2 => n3829, ZN => n4036);
   U5329 : AOI21_X1 port map( B1 => n3830, B2 => n4036, A => n4131, ZN => n3831
                           );
   U5330 : AOI211_X1 port map( C1 => n4125, C2 => n3832, A => n3831, B => n3908
                           , ZN => n3833);
   U5331 : OAI211_X1 port map( C1 => n3835, C2 => n3851, A => n3834, B => n3833
                           , ZN => n3836);
   U5332 : AOI211_X1 port map( C1 => n4135, C2 => n3838, A => n3837, B => n3836
                           , ZN => n3843);
   U5333 : NOR3_X1 port map( A1 => n3840, A2 => n4148, A3 => n3839, ZN => n3841
                           );
   U5334 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_29, A => n3841, ZN 
                           => n3842);
   U5335 : OAI21_X1 port map( B1 => n3843, B2 => n4154, A => n3842, ZN => 
                           IF_ALUxN967);
   U5336 : NAND2_X1 port map( A1 => ALUtoCtl_port_28_port, A2 => n4413, ZN => 
                           n3845);
   U5337 : OAI211_X1 port map( C1 => n3925, C2 => n4086, A => n3845, B => n3844
                           , ZN => n6491);
   U5338 : NOR3_X1 port map( A1 => n3846, A2 => n4148, A3 => n4033, ZN => n3871
                           );
   U5339 : AOI21_X1 port map( B1 => CtlToALU_port_alu_fun_0_port, B2 => n4032, 
                           A => IF_ALUxN140, ZN => n3849);
   U5340 : AND2_X1 port map( A1 => n4032, A2 => n4033, ZN => n3847);
   U5341 : NOR2_X1 port map( A1 => n4033, A2 => n4032, ZN => n4035);
   U5342 : OAI21_X1 port map( B1 => n3847, B2 => n4035, A => n4073, ZN => n3848
                           );
   U5343 : OAI211_X1 port map( C1 => n3849, C2 => n4123, A => n3882, B => n3848
                           , ZN => n3854);
   U5344 : OAI22_X1 port map( A1 => n3852, A2 => n3851, B1 => n3850, B2 => 
                           n3894, ZN => n3853);
   U5345 : AOI211_X1 port map( C1 => n4125, C2 => n3855, A => n3854, B => n3853
                           , ZN => n3869);
   U5346 : AOI22_X1 port map( A1 => n4120, A2 => n3858, B1 => n3857, B2 => 
                           n3856, ZN => n3885);
   U5347 : AOI221_X1 port map( B1 => n3861, B2 => n3860, C1 => n3859, C2 => 
                           n4118, A => n4051, ZN => n3863);
   U5348 : AOI211_X1 port map( C1 => n3864, C2 => n3885, A => n3863, B => n3862
                           , ZN => n3865);
   U5349 : OAI21_X1 port map( B1 => n3867, B2 => n3866, A => n3865, ZN => n3868
                           );
   U5350 : AOI21_X1 port map( B1 => n3869, B2 => n3868, A => n4154, ZN => n3870
                           );
   U5351 : AOI211_X1 port map( C1 => n4152, C2 => C596xDATA2_28, A => n3871, B 
                           => n3870, ZN => n3872);
   U5352 : INV_X1 port map( A => n3872, ZN => IF_ALUxN966);
   U5353 : NAND2_X1 port map( A1 => ALUtoCtl_port_24_port, A2 => n4413, ZN => 
                           n3874);
   U5354 : OAI211_X1 port map( C1 => n3925, C2 => n4090, A => n3874, B => n3873
                           , ZN => n6493);
   U5355 : AOI22_X1 port map( A1 => n3878, A2 => n3877, B1 => n3876, B2 => 
                           n3875, ZN => n3913);
   U5356 : AOI22_X1 port map( A1 => n3912, A2 => n3913, B1 => n3880, B2 => 
                           n3879, ZN => n3893);
   U5357 : NOR2_X1 port map( A1 => n4020, A2 => IF_ALUxN136, ZN => n3938);
   U5358 : AOI21_X1 port map( B1 => n4020, B2 => IF_ALUxN136, A => n3938, ZN =>
                           n3884);
   U5359 : AOI22_X1 port map( A1 => n4060, A2 => IF_ALUxN136, B1 => n4127, B2 
                           => n3881, ZN => n3883);
   U5360 : OAI211_X1 port map( C1 => n3884, C2 => n4131, A => n3883, B => n3882
                           , ZN => n3889);
   U5361 : OAI22_X1 port map( A1 => n3887, A2 => n3886, B1 => n3885, B2 => 
                           n4117, ZN => n3888);
   U5362 : AOI211_X1 port map( C1 => n3891, C2 => n3890, A => n3889, B => n3888
                           , ZN => n3892);
   U5363 : OAI211_X1 port map( C1 => n3895, C2 => n3894, A => n3893, B => n3892
                           , ZN => n3896);
   U5364 : INV_X1 port map( A => n3896, ZN => n3900);
   U5365 : NOR3_X1 port map( A1 => n4020, A2 => n4148, A3 => n3897, ZN => n3898
                           );
   U5366 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_24, A => n3898, ZN 
                           => n3899);
   U5367 : OAI21_X1 port map( B1 => n4078, B2 => n3900, A => n3899, ZN => 
                           IF_ALUxN962);
   U5368 : NAND2_X1 port map( A1 => ALUtoCtl_port_16_port, A2 => n4413, ZN => 
                           n3902);
   U5369 : OAI211_X1 port map( C1 => n3925, C2 => n4098, A => n3902, B => n3901
                           , ZN => n6495);
   U5370 : AOI22_X1 port map( A1 => n3954, A2 => n3904, B1 => n3903, B2 => 
                           n4056, ZN => n4061);
   U5371 : INV_X1 port map( A => n4061, ZN => n3917);
   U5372 : NOR2_X1 port map( A1 => n4004, A2 => n4003, ZN => n3998);
   U5373 : AOI21_X1 port map( B1 => n4004, B2 => n4003, A => n3998, ZN => n3906
                           );
   U5374 : AOI21_X1 port map( B1 => CtlToALU_port_alu_fun_0_port, B2 => n4003, 
                           A => IF_ALUxN128, ZN => n3905);
   U5375 : OAI22_X1 port map( A1 => n3906, A2 => n4131, B1 => n3905, B2 => 
                           n4123, ZN => n3907);
   U5376 : AOI211_X1 port map( C1 => n3910, C2 => n3909, A => n3908, B => n3907
                           , ZN => n3916);
   U5377 : AOI22_X1 port map( A1 => n3914, A2 => n3913, B1 => n3912, B2 => 
                           n3911, ZN => n3915);
   U5378 : OAI211_X1 port map( C1 => n4055, C2 => n3917, A => n3916, B => n3915
                           , ZN => n3918);
   U5379 : INV_X1 port map( A => n3918, ZN => n3922);
   U5380 : NOR3_X1 port map( A1 => n3919, A2 => n4148, A3 => n4004, ZN => n3920
                           );
   U5381 : AOI21_X1 port map( B1 => n4152, B2 => C596xDATA2_16, A => n3920, ZN 
                           => n3921);
   U5382 : OAI21_X1 port map( B1 => n4078, B2 => n3922, A => n3921, ZN => 
                           IF_ALUxN954);
   U5383 : NAND2_X1 port map( A1 => ALUtoCtl_port_0_port, A2 => n4413, ZN => 
                           n3924);
   U5384 : OAI211_X1 port map( C1 => n3925, C2 => n4114, A => n3924, B => n3923
                           , ZN => n6497);
   U5385 : NOR2_X1 port map( A1 => n3926, A2 => n4148, ZN => n4083);
   U5386 : NOR2_X1 port map( A1 => n4116, A2 => IF_ALUxN112, ZN => n4081);
   U5387 : NOR2_X1 port map( A1 => n4131, A2 => n3927, ZN => n4076);
   U5388 : NOR2_X1 port map( A1 => n4045, A2 => IF_ALUxN112, ZN => n3957);
   U5389 : INV_X1 port map( A => n3957, ZN => n4075);
   U5390 : NAND2_X1 port map( A1 => n3929, A2 => n3928, ZN => n4071);
   U5391 : AOI222_X1 port map( A1 => n3932, A2 => 
                           CtlToALU_port_reg2_contents_31_port, B1 => n3931, B2
                           => CtlToALU_port_pc_reg_31_port, C1 => n3930, C2 => 
                           CtlToALU_port_imm_31_port, ZN => n4149);
   U5392 : INV_X1 port map( A => n4149, ZN => n4143);
   U5393 : NOR2_X1 port map( A1 => n4147, A2 => n4143, ZN => n4124);
   U5394 : INV_X1 port map( A => n3933, ZN => n4026);
   U5395 : AOI21_X1 port map( B1 => n3934, B2 => IF_ALUxN134, A => n3935, ZN =>
                           n4013);
   U5396 : AOI21_X1 port map( B1 => n3937, B2 => n3936, A => n3935, ZN => n3939
                           );
   U5397 : AOI211_X1 port map( C1 => n4013, C2 => n3940, A => n3939, B => n3938
                           , ZN => n4022);
   U5398 : OAI22_X1 port map( A1 => n3944, A2 => n3943, B1 => n3942, B2 => 
                           n3941, ZN => n3977);
   U5399 : INV_X1 port map( A => n3977, ZN => n3990);
   U5400 : OAI211_X1 port map( C1 => n3980, C2 => n3947, A => n3946, B => n3945
                           , ZN => n3989);
   U5401 : NOR2_X1 port map( A1 => n3948, A2 => IF_ALUxN127, ZN => n3988);
   U5402 : AOI22_X1 port map( A1 => n3952, A2 => n3951, B1 => n3950, B2 => 
                           n3949, ZN => n3986);
   U5403 : AOI22_X1 port map( A1 => n3954, A2 => IF_ALUxN115, B1 => n3953, B2 
                           => IF_ALUxN116, ZN => n3964);
   U5404 : OAI211_X1 port map( C1 => n3958, C2 => n3957, A => n3956, B => n3955
                           , ZN => n3960);
   U5405 : OAI211_X1 port map( C1 => n3954, C2 => IF_ALUxN115, A => n3960, B =>
                           n3959, ZN => n3963);
   U5406 : AOI211_X1 port map( C1 => n3964, C2 => n3963, A => n3962, B => n3961
                           , ZN => n3972);
   U5407 : OAI22_X1 port map( A1 => n3968, A2 => n3967, B1 => n3966, B2 => 
                           n3965, ZN => n3971);
   U5408 : OAI211_X1 port map( C1 => n3972, C2 => n3971, A => n3970, B => n3969
                           , ZN => n3974);
   U5409 : OAI211_X1 port map( C1 => n3976, C2 => n3975, A => n3974, B => n3973
                           , ZN => n3985);
   U5410 : NOR4_X1 port map( A1 => n3980, A2 => n3979, A3 => n3978, A4 => n3977
                           , ZN => n3991);
   U5411 : OAI211_X1 port map( C1 => n3983, C2 => n3982, A => n3991, B => n3981
                           , ZN => n3984);
   U5412 : AOI21_X1 port map( B1 => n3986, B2 => n3985, A => n3984, ZN => n3987
                           );
   U5413 : AOI211_X1 port map( C1 => n3990, C2 => n3989, A => n3988, B => n3987
                           , ZN => n4000);
   U5414 : OAI21_X1 port map( B1 => n3993, B2 => n3992, A => n3991, ZN => n3999
                           );
   U5415 : NAND2_X1 port map( A1 => n3994, A2 => IF_ALUxN131, ZN => n4005);
   U5416 : OAI211_X1 port map( C1 => n3997, C2 => n3996, A => n3995, B => n4005
                           , ZN => n4011);
   U5417 : AOI211_X1 port map( C1 => n4000, C2 => n3999, A => n3998, B => n4011
                           , ZN => n4019);
   U5418 : AOI22_X1 port map( A1 => n4004, A2 => n4003, B1 => n4002, B2 => 
                           n4001, ZN => n4012);
   U5419 : AOI22_X1 port map( A1 => n4008, A2 => n4007, B1 => n4006, B2 => 
                           n4005, ZN => n4010);
   U5420 : OAI211_X1 port map( C1 => n4012, C2 => n4011, A => n4010, B => n4009
                           , ZN => n4018);
   U5421 : INV_X1 port map( A => n4013, ZN => n4014);
   U5422 : AOI211_X1 port map( C1 => n4016, C2 => IF_ALUxN132, A => n4015, B =>
                           n4014, ZN => n4017);
   U5423 : OAI21_X1 port map( B1 => n4019, B2 => n4018, A => n4017, ZN => n4021
                           );
   U5424 : AOI22_X1 port map( A1 => n4022, A2 => n4021, B1 => n4020, B2 => 
                           IF_ALUxN136, ZN => n4025);
   U5425 : OAI211_X1 port map( C1 => n4026, C2 => n4025, A => n4024, B => n4023
                           , ZN => n4027);
   U5426 : AOI22_X1 port map( A1 => n4029, A2 => IF_ALUxN139, B1 => n4028, B2 
                           => n4027, ZN => n4030);
   U5427 : AOI211_X1 port map( C1 => n4033, C2 => n4032, A => n4031, B => n4030
                           , ZN => n4037);
   U5428 : AOI221_X1 port map( B1 => n4037, B2 => n4036, C1 => n4035, C2 => 
                           n4036, A => n4034, ZN => n4039);
   U5429 : AOI22_X1 port map( A1 => n4041, A2 => n4040, B1 => n4039, B2 => 
                           n4038, ZN => n4044);
   U5430 : INV_X1 port map( A => n4044, ZN => n4042);
   U5431 : NAND2_X1 port map( A1 => n4147, A2 => n4143, ZN => n4130);
   U5432 : OAI21_X1 port map( B1 => n4124, B2 => n4042, A => n4130, ZN => n4070
                           );
   U5433 : NOR3_X1 port map( A1 => CtlToALU_port_alu_fun_0_port, A2 => n6246, 
                           A3 => n4043, ZN => n4058);
   U5434 : OAI211_X1 port map( C1 => n4124, C2 => n4044, A => n4058, B => n4130
                           , ZN => n4068);
   U5435 : NOR2_X1 port map( A1 => n4045, A2 => IF_ALUxN113, ZN => n4046);
   U5436 : NOR2_X1 port map( A1 => n4046, A2 => n4081, ZN => n4049);
   U5437 : INV_X1 port map( A => n4047, ZN => n4048);
   U5438 : MUX2_X1 port map( A => n4049, B => n4048, S => n4118, Z => n4050);
   U5439 : OAI22_X1 port map( A1 => n4053, A2 => n4052, B1 => n4051, B2 => 
                           n4050, ZN => n4054);
   U5440 : AOI211_X1 port map( C1 => n4057, C2 => n4056, A => n4055, B => n4054
                           , ZN => n4059);
   U5441 : AOI211_X1 port map( C1 => n4060, C2 => IF_ALUxN112, A => n4059, B =>
                           n4058, ZN => n4065);
   U5442 : OAI21_X1 port map( B1 => n4063, B2 => n4062, A => n4061, ZN => n4064
                           );
   U5443 : OAI211_X1 port map( C1 => n4117, C2 => n4066, A => n4065, B => n4064
                           , ZN => n4067);
   U5444 : NAND3_X1 port map( A1 => n4071, A2 => n4068, A3 => n4067, ZN => 
                           n4069);
   U5445 : OAI21_X1 port map( B1 => n4071, B2 => n4070, A => n4069, ZN => n4072
                           );
   U5446 : NOR2_X1 port map( A1 => n4073, A2 => n4072, ZN => n4074);
   U5447 : AOI21_X1 port map( B1 => n4076, B2 => n4075, A => n4074, ZN => n4077
                           );
   U5448 : INV_X1 port map( A => n4077, ZN => n4080);
   U5449 : AOI221_X1 port map( B1 => n4081, B2 => n4127, C1 => n4080, C2 => 
                           n4079, A => n4078, ZN => n4082);
   U5450 : AOI211_X1 port map( C1 => n4152, C2 => C596xDATA2_0, A => n4083, B 
                           => n4082, ZN => n4084);
   U5451 : INV_X1 port map( A => n4084, ZN => IF_ALUxN938);
   U5452 : NOR2_X1 port map( A1 => rst, A2 => n4085, ZN => IF_CPathxN2271);
   U5453 : NOR2_X1 port map( A1 => rst, A2 => n4086, ZN => IF_CPathxN2270);
   U5454 : NOR2_X1 port map( A1 => rst, A2 => n4087, ZN => IF_CPathxN2269);
   U5455 : NOR2_X1 port map( A1 => rst, A2 => n4088, ZN => IF_CPathxN2268);
   U5456 : NOR2_X1 port map( A1 => rst, A2 => n4089, ZN => IF_CPathxN2267);
   U5457 : NOR2_X1 port map( A1 => rst, A2 => n4090, ZN => IF_CPathxN2266);
   U5458 : NOR2_X1 port map( A1 => rst, A2 => n4091, ZN => IF_CPathxN2265);
   U5459 : NOR2_X1 port map( A1 => rst, A2 => n4092, ZN => IF_CPathxN2264);
   U5460 : NOR2_X1 port map( A1 => rst, A2 => n4093, ZN => IF_CPathxN2263);
   U5461 : NOR2_X1 port map( A1 => rst, A2 => n4094, ZN => IF_CPathxN2262);
   U5462 : NOR2_X1 port map( A1 => rst, A2 => n4095, ZN => IF_CPathxN2261);
   U5463 : NOR2_X1 port map( A1 => rst, A2 => n4096, ZN => IF_CPathxN2260);
   U5464 : NOR2_X1 port map( A1 => rst, A2 => n4097, ZN => IF_CPathxN2259);
   U5465 : NOR2_X1 port map( A1 => rst, A2 => n4098, ZN => IF_CPathxN2258);
   U5466 : NOR2_X1 port map( A1 => rst, A2 => n4099, ZN => IF_CPathxN2257);
   U5467 : NOR2_X1 port map( A1 => rst, A2 => n4100, ZN => IF_CPathxN2256);
   U5468 : NOR2_X1 port map( A1 => rst, A2 => n4101, ZN => IF_CPathxN2255);
   U5469 : NOR2_X1 port map( A1 => rst, A2 => n4102, ZN => IF_CPathxN2254);
   U5470 : NOR2_X1 port map( A1 => rst, A2 => n4103, ZN => IF_CPathxN2253);
   U5471 : NOR2_X1 port map( A1 => rst, A2 => n4104, ZN => IF_CPathxN2252);
   U5472 : NOR2_X1 port map( A1 => rst, A2 => n4105, ZN => IF_CPathxN2251);
   U5473 : NOR2_X1 port map( A1 => rst, A2 => n4106, ZN => IF_CPathxN2250);
   U5474 : NOR2_X1 port map( A1 => rst, A2 => n4107, ZN => IF_CPathxN2249);
   U5475 : NOR2_X1 port map( A1 => rst, A2 => n4108, ZN => IF_CPathxN2248);
   U5476 : NOR2_X1 port map( A1 => rst, A2 => n4109, ZN => IF_CPathxN2247);
   U5477 : NOR2_X1 port map( A1 => rst, A2 => n4110, ZN => IF_CPathxN2246);
   U5478 : NOR2_X1 port map( A1 => rst, A2 => n4111, ZN => IF_CPathxN2245);
   U5479 : NOR2_X1 port map( A1 => rst, A2 => n4112, ZN => IF_CPathxN2244);
   U5480 : NOR2_X1 port map( A1 => rst, A2 => n4113, ZN => IF_CPathxN2243);
   U5481 : NOR2_X1 port map( A1 => rst, A2 => n4114, ZN => IF_CPathxN2242);
   U5482 : AOI21_X1 port map( B1 => n4116, B2 => IF_ALUxN142, A => n4115, ZN =>
                           n4121);
   U5483 : AOI221_X1 port map( B1 => n4121, B2 => n4120, C1 => n4119, C2 => 
                           n4118, A => n4117, ZN => n4140);
   U5484 : AOI21_X1 port map( B1 => n4123, B2 => n4122, A => n4147, ZN => n4133
                           );
   U5485 : INV_X1 port map( A => n4124, ZN => n4129);
   U5486 : AOI22_X1 port map( A1 => n4127, A2 => n4143, B1 => n4126, B2 => 
                           n4125, ZN => n4128);
   U5487 : OAI221_X1 port map( B1 => n4131, B2 => n4130, C1 => n4131, C2 => 
                           n4129, A => n4128, ZN => n4132);
   U5488 : AOI211_X1 port map( C1 => n4135, C2 => n4134, A => n4133, B => n4132
                           , ZN => n4136);
   U5489 : OAI21_X1 port map( B1 => n4138, B2 => n4137, A => n4136, ZN => n4139
                           );
   U5490 : AOI211_X1 port map( C1 => n4142, C2 => n4141, A => n4140, B => n4139
                           , ZN => n4155);
   U5491 : XOR2_X1 port map( A => n6378, B => n4143, Z => n4145);
   U5492 : XOR2_X1 port map( A => n4145, B => n4144, Z => n4146);
   U5493 : XOR2_X1 port map( A => DP_OP_1698J95_122_4028xn2, B => n4146, Z => 
                           n4151);
   U5494 : NOR3_X1 port map( A1 => n4149, A2 => n4148, A3 => n4147, ZN => n4150
                           );
   U5495 : AOI21_X1 port map( B1 => n4152, B2 => n4151, A => n4150, ZN => n4153
                           );
   U5496 : OAI21_X1 port map( B1 => n4155, B2 => n4154, A => n4153, ZN => 
                           IF_ALUxN969);
   U5497 : AOI22_X1 port map( A1 => n4277, A2 => IF_CPathxN2162, B1 => n4210, 
                           B2 => IF_CPathxDecToCtl_data_signal_imm_4_port, ZN 
                           => n4156);
   U5498 : INV_X1 port map( A => n4156, ZN => n6670);
   U5499 : AOI22_X1 port map( A1 => n4277, A2 => IF_CPathxN2160, B1 => n4210, 
                           B2 => IF_CPathxDecToCtl_data_signal_imm_2_port, ZN 
                           => n4157);
   U5500 : INV_X1 port map( A => n4157, ZN => n6672);
   U5501 : AOI22_X1 port map( A1 => n4277, A2 => IF_CPathxN2159, B1 => n4210, 
                           B2 => IF_CPathxDecToCtl_data_signal_imm_1_port, ZN 
                           => n4158);
   U5502 : INV_X1 port map( A => n4158, ZN => n6673);
   U5503 : AOI22_X1 port map( A1 => n4277, A2 => IF_CPathxN2158, B1 => n4210, 
                           B2 => IF_CPathxDecToCtl_data_signal_imm_0_port, ZN 
                           => n4159);
   U5504 : INV_X1 port map( A => n4159, ZN => n6674);
   U5505 : NOR2_X1 port map( A1 => rst, A2 => n6274, ZN => IF_DecoderxN602);
   U5506 : AND2_X1 port map( A1 => CtlToDec_port_5_port, A2 => n6234, ZN => 
                           n4562);
   U5507 : NAND2_X1 port map( A1 => CtlToDec_port_6_port, A2 => n4562, ZN => 
                           n4565);
   U5508 : NOR2_X1 port map( A1 => n6229, A2 => n4565, ZN => n4595);
   U5509 : NAND2_X1 port map( A1 => n4595, A2 => IF_DecoderxN602, ZN => n4173);
   U5510 : NOR3_X1 port map( A1 => rst, A2 => CtlToDec_port_5_port, A3 => 
                           CtlToDec_port_2_port, ZN => n4162);
   U5511 : NAND3_X1 port map( A1 => n4571, A2 => n6229, A3 => n4562, ZN => 
                           n4163);
   U5512 : INV_X1 port map( A => n4163, ZN => n4160);
   U5513 : AOI22_X1 port map( A1 => n4162, A2 => CtlToDec_port_20_port, B1 => 
                           CtlToDec_port_7_port, B2 => n4160, ZN => n4161);
   U5514 : AOI221_X1 port map( B1 => CtlToDec_port_6_port, B2 => n4173, C1 => 
                           n4161, C2 => n4173, A => CtlToDec_port_3_port, ZN =>
                           n6719);
   U5515 : INV_X1 port map( A => n4162, ZN => n4648);
   U5516 : NOR2_X1 port map( A1 => rst, A2 => n6229, ZN => n4176);
   U5517 : NAND2_X1 port map( A1 => n4562, A2 => n4176, ZN => n4167);
   U5518 : AND2_X1 port map( A1 => n4648, A2 => n4167, ZN => n4164);
   U5519 : OAI22_X1 port map( A1 => n4164, A2 => n6210, B1 => n4163, B2 => 
                           n6319, ZN => n6718);
   U5520 : OAI22_X1 port map( A1 => n4164, A2 => n6211, B1 => n4163, B2 => 
                           n6320, ZN => n6717);
   U5521 : OAI22_X1 port map( A1 => n4164, A2 => n6212, B1 => n4163, B2 => 
                           n6321, ZN => n6716);
   U5522 : OAI22_X1 port map( A1 => n4164, A2 => n6213, B1 => n4163, B2 => 
                           n6322, ZN => n6715);
   U5523 : NAND2_X1 port map( A1 => n6208, A2 => n6261, ZN => n4617);
   U5524 : NOR2_X1 port map( A1 => n4617, A2 => n6259, ZN => n4613);
   U5525 : AOI221_X1 port map( B1 => CtlToDec_port_5_port, B2 => 
                           CtlToDec_port_4_port, C1 => n4613, C2 => 
                           CtlToDec_port_4_port, A => rst, ZN => n4168);
   U5526 : OAI21_X1 port map( B1 => n4562, B2 => n6229, A => n4168, ZN => n4180
                           );
   U5527 : NOR2_X1 port map( A1 => n6264, A2 => n4180, ZN => n6714);
   U5528 : NOR2_X1 port map( A1 => n6273, A2 => n4180, ZN => n6713);
   U5529 : NOR2_X1 port map( A1 => n6271, A2 => n4180, ZN => n6712);
   U5530 : NOR2_X1 port map( A1 => n6272, A2 => n4180, ZN => n6711);
   U5531 : NOR2_X1 port map( A1 => n6270, A2 => n4180, ZN => n6710);
   U5532 : NOR2_X1 port map( A1 => CtlToDec_port_13_port, A2 => n6261, ZN => 
                           n4628);
   U5533 : NOR4_X1 port map( A1 => CtlToDec_port_26_port, A2 => 
                           CtlToDec_port_28_port, A3 => CtlToDec_port_27_port, 
                           A4 => CtlToDec_port_29_port, ZN => n4165);
   U5534 : NAND3_X1 port map( A1 => n4165, A2 => n6264, A3 => n6209, ZN => 
                           n4582);
   U5535 : INV_X1 port map( A => n4582, ZN => n4578);
   U5536 : NAND3_X1 port map( A1 => n4628, A2 => CtlToDec_port_12_port, A3 => 
                           n4578, ZN => n4638);
   U5537 : INV_X1 port map( A => n4638, ZN => n4166);
   U5538 : AOI211_X1 port map( C1 => CtlToDec_port_4_port, C2 => n4166, A => 
                           n6260, B => n4180, ZN => n6709);
   U5539 : NOR2_X1 port map( A1 => n6209, A2 => n4167, ZN => n4171);
   U5540 : NAND2_X1 port map( A1 => CtlToDec_port_31_port, A2 => n4168, ZN => 
                           n4169);
   U5541 : NAND2_X1 port map( A1 => CtlToDec_port_7_port, A2 => n6178, ZN => 
                           n4640);
   U5542 : OAI22_X1 port map( A1 => CtlToDec_port_6_port, A2 => n4169, B1 => 
                           n4640, B2 => n4565, ZN => n4170);
   U5543 : AOI22_X1 port map( A1 => CtlToDec_port_6_port, A2 => n4171, B1 => 
                           n6229, B2 => n4170, ZN => n4172);
   U5544 : AOI22_X1 port map( A1 => CtlToDec_port_3_port, A2 => n4173, B1 => 
                           n4172, B2 => n6231, ZN => n6708);
   U5545 : OAI221_X1 port map( B1 => CtlToDec_port_3_port, B2 => 
                           CtlToDec_port_4_port, C1 => n6231, C2 => n4562, A =>
                           n4176, ZN => n4175);
   U5546 : NOR2_X1 port map( A1 => n6209, A2 => n4180, ZN => n4177);
   U5547 : NAND2_X1 port map( A1 => n4177, A2 => n6231, ZN => n4174);
   U5548 : OAI21_X1 port map( B1 => n6259, B2 => n4175, A => n4174, ZN => n6707
                           );
   U5549 : OAI21_X1 port map( B1 => n6208, B2 => n4175, A => n4174, ZN => n6706
                           );
   U5550 : OAI21_X1 port map( B1 => n6261, B2 => n4175, A => n4174, ZN => n6705
                           );
   U5551 : OAI21_X1 port map( B1 => n4175, B2 => n6324, A => n4174, ZN => n6704
                           );
   U5552 : OAI21_X1 port map( B1 => n4175, B2 => n6325, A => n4174, ZN => n6703
                           );
   U5553 : OAI21_X1 port map( B1 => n4175, B2 => n6326, A => n4174, ZN => n6702
                           );
   U5554 : OAI21_X1 port map( B1 => n4175, B2 => n6327, A => n4174, ZN => n6701
                           );
   U5555 : OAI21_X1 port map( B1 => n4175, B2 => n6328, A => n4174, ZN => n6700
                           );
   U5556 : NAND2_X1 port map( A1 => CtlToDec_port_4_port, A2 => n4176, ZN => 
                           n4179);
   U5557 : INV_X1 port map( A => n4177, ZN => n4178);
   U5558 : OAI21_X1 port map( B1 => n6274, B2 => n4179, A => n4178, ZN => n6699
                           );
   U5559 : OAI21_X1 port map( B1 => n4179, B2 => n6210, A => n4178, ZN => n6698
                           );
   U5560 : OAI21_X1 port map( B1 => n4179, B2 => n6211, A => n4178, ZN => n6697
                           );
   U5561 : OAI21_X1 port map( B1 => n4179, B2 => n6212, A => n4178, ZN => n6696
                           );
   U5562 : OAI21_X1 port map( B1 => n4179, B2 => n6213, A => n4178, ZN => n6695
                           );
   U5563 : OAI21_X1 port map( B1 => n6264, B2 => n4179, A => n4178, ZN => n6694
                           );
   U5564 : OAI21_X1 port map( B1 => n6273, B2 => n4179, A => n4178, ZN => n6693
                           );
   U5565 : OAI21_X1 port map( B1 => n6271, B2 => n4179, A => n4178, ZN => n6692
                           );
   U5566 : OAI21_X1 port map( B1 => n6272, B2 => n4179, A => n4178, ZN => n6691
                           );
   U5567 : OAI21_X1 port map( B1 => n6270, B2 => n4179, A => n4178, ZN => n6690
                           );
   U5568 : OAI21_X1 port map( B1 => n6260, B2 => n4179, A => n4178, ZN => n6689
                           );
   U5569 : AOI21_X1 port map( B1 => n4180, B2 => n4179, A => n6209, ZN => n6688
                           );
   U5570 : NAND2_X1 port map( A1 => n4571, A2 => n6228, ZN => n6185);
   U5571 : AOI21_X1 port map( B1 => n6185, B2 => n4268, A => 
                           IF_CPathxsection_0_port, ZN => n6687);
   U5572 : INV_X1 port map( A => n4188, ZN => n4549);
   U5573 : NAND2_X1 port map( A1 => n4181, A2 => n4549, ZN => n4207);
   U5574 : OAI21_X1 port map( B1 => n4549, B2 => n4282, A => n4207, ZN => n6686
                           );
   U5575 : NOR2_X1 port map( A1 => n6196, A2 => IF_CPathxsection_3_port, ZN => 
                           n4445);
   U5576 : NOR2_X1 port map( A1 => IF_CPathxsection_2_port, A2 => n6228, ZN => 
                           n4554);
   U5577 : NOR2_X1 port map( A1 => n4445, A2 => n4554, ZN => n4416);
   U5578 : NOR2_X1 port map( A1 => rst, A2 => n4416, ZN => n6546);
   U5579 : NOR3_X1 port map( A1 => n6197, A2 => n6230, A3 => 
                           DecToCtl_port_encType_1_port, ZN => n4464);
   U5580 : NAND2_X1 port map( A1 => n4571, A2 => n4464, ZN => n4406);
   U5581 : NAND2_X1 port map( A1 => n2953, A2 => DecToCtl_port_instrType_0_port
                           , ZN => n4247);
   U5582 : AOI211_X1 port map( C1 => DecToCtl_port_instrType_2_port, C2 => 
                           n4247, A => DecToCtl_port_instrType_3_port, B => 
                           n6191, ZN => n4183);
   U5583 : NOR2_X1 port map( A1 => n6195, A2 => n6232, ZN => n4254);
   U5584 : NAND2_X1 port map( A1 => DecToCtl_port_instrType_3_port, A2 => 
                           DecToCtl_port_instrType_1_port, ZN => n4267);
   U5585 : AOI22_X1 port map( A1 => DecToCtl_port_instrType_3_port, A2 => 
                           DecToCtl_port_instrType_4_port, B1 => n4182, B2 => 
                           n4267, ZN => n4261);
   U5586 : OAI221_X1 port map( B1 => n4183, B2 => n4254, C1 => n4183, C2 => 
                           n4261, A => n6226, ZN => n4199);
   U5587 : INV_X1 port map( A => n4247, ZN => n4524);
   U5588 : NOR4_X1 port map( A1 => n6189, A2 => n6191, A3 => 
                           DecToCtl_port_instrType_5_port, A4 => 
                           DecToCtl_port_instrType_2_port, ZN => n4458);
   U5589 : INV_X1 port map( A => n4458, ZN => n4525);
   U5590 : NAND3_X1 port map( A1 => DecToCtl_port_instrType_5_port, A2 => n6189
                           , A3 => n6191, ZN => n4523);
   U5591 : NAND2_X1 port map( A1 => n4525, A2 => n4523, ZN => n4457);
   U5592 : NAND3_X1 port map( A1 => DecToCtl_port_instrType_2_port, A2 => 
                           DecToCtl_port_instrType_4_port, A3 => n4244, ZN => 
                           n4526);
   U5593 : NOR2_X1 port map( A1 => DecToCtl_port_encType_2_port, A2 => 
                           DecToCtl_port_encType_0_port, ZN => n4224);
   U5594 : INV_X1 port map( A => n4224, ZN => n4230);
   U5595 : NOR2_X1 port map( A1 => n4230, A2 => n6225, ZN => n4543);
   U5596 : OAI221_X1 port map( B1 => n4532, B2 => n4526, C1 => n4184, C2 => 
                           n4460, A => n4543, ZN => n4185);
   U5597 : AOI221_X1 port map( B1 => n4527, B2 => n4524, C1 => n4457, C2 => 
                           n4524, A => n4185, ZN => n4200);
   U5598 : INV_X1 port map( A => n4200, ZN => n4186);
   U5599 : NOR3_X1 port map( A1 => n6191, A2 => n4199, A3 => n4186, ZN => n4462
                           );
   U5600 : NOR2_X1 port map( A1 => IF_CPathxsection_3_port, A2 => n4281, ZN => 
                           n4402);
   U5601 : NAND2_X1 port map( A1 => n4549, A2 => n4402, ZN => n4192);
   U5602 : INV_X1 port map( A => n6185, ZN => n4187);
   U5603 : NOR2_X1 port map( A1 => IF_CPathxsection_2_port, A2 => n4275, ZN => 
                           n4195);
   U5604 : INV_X1 port map( A => n4195, ZN => n6187);
   U5605 : NOR2_X1 port map( A1 => IF_CPathxsection_0_port, A2 => n6187, ZN => 
                           n6186);
   U5606 : AOI22_X1 port map( A1 => n4187, A2 => n4188, B1 => n6186, B2 => 
                           n4546, ZN => n4191);
   U5607 : NAND2_X1 port map( A1 => IF_CPathxsection_0_port, A2 => n4195, ZN =>
                           n6184);
   U5608 : INV_X1 port map( A => n6184, ZN => n4446);
   U5609 : INV_X1 port map( A => n4445, ZN => n4208);
   U5610 : NOR2_X1 port map( A1 => n4188, A2 => n4208, ZN => n4548);
   U5611 : AOI21_X1 port map( B1 => n4446, B2 => IF_CPathxsection_3_port, A => 
                           n4548, ZN => n4198);
   U5612 : NAND4_X1 port map( A1 => n6236, A2 => n6200, A3 => n6192, A4 => 
                           n6190, ZN => n4189);
   U5613 : OAI21_X1 port map( B1 => 
                           IF_CPathxDecToCtl_data_signal_rd_addr_4_port, B2 => 
                           n4189, A => IF_CPathxwb_en_signal, ZN => n4447);
   U5614 : NOR2_X1 port map( A1 => n4198, A2 => n4447, ZN => n4553);
   U5615 : OAI21_X1 port map( B1 => n4413, B2 => n4553, A => n6546, ZN => n4190
                           );
   U5616 : OAI211_X1 port map( C1 => n4462, C2 => n4192, A => n4191, B => n4190
                           , ZN => n4193);
   U5617 : INV_X1 port map( A => n4193, ZN => n4194);
   U5618 : OAI22_X1 port map( A1 => n4521, A2 => n4406, B1 => n6286, B2 => 
                           n4194, ZN => n6685);
   U5619 : INV_X1 port map( A => n4447, ZN => n4451);
   U5620 : NOR2_X1 port map( A1 => n6227, A2 => IF_CPathxsection_0_port, ZN => 
                           n4203);
   U5621 : AOI21_X1 port map( B1 => n4554, B2 => n4203, A => rst, ZN => n4561);
   U5622 : NOR2_X1 port map( A1 => IF_CPathxsection_3_port, A2 => n4195, ZN => 
                           n4558);
   U5623 : NAND2_X1 port map( A1 => IF_CPathxmem_en_signal, A2 => n4548, ZN => 
                           n4556);
   U5624 : INV_X1 port map( A => n4556, ZN => n4196);
   U5625 : AOI221_X1 port map( B1 => n4446, B2 => CtlToMem_port_notify_port, C1
                           => n4558, C2 => CtlToMem_port_notify_port, A => 
                           n4196, ZN => n4197);
   U5626 : OAI211_X1 port map( C1 => n4451, C2 => n4198, A => n4561, B => n4197
                           , ZN => n6684);
   U5627 : NAND2_X1 port map( A1 => n4454, A2 => n4443, ZN => n4440);
   U5628 : INV_X1 port map( A => n4440, ZN => n4201);
   U5629 : AOI21_X1 port map( B1 => DecToCtl_port_encType_2_port, B2 => 
                           DecToCtl_port_encType_1_port, A => 
                           DecToCtl_port_encType_0_port, ZN => n4456);
   U5630 : NAND2_X1 port map( A1 => n4200, A2 => n4199, ZN => n4540);
   U5631 : AND2_X1 port map( A1 => n4456, A2 => n4540, ZN => n4453);
   U5632 : AOI211_X1 port map( C1 => n4201, C2 => IF_CPathxreg_rd_en_signal, A 
                           => n4453, B => n4464, ZN => n4202);
   U5633 : INV_X1 port map( A => n4202, ZN => n4444);
   U5634 : NAND3_X1 port map( A1 => IF_CPathxsection_0_port, A2 => n4279, A3 =>
                           n6227, ZN => n4206);
   U5635 : INV_X1 port map( A => n4203, ZN => n4204);
   U5636 : OAI211_X1 port map( C1 => n6196, C2 => n4204, A => 
                           CtlToALU_port_notify, B => n4547, ZN => n4205);
   U5637 : OAI211_X1 port map( C1 => n4207, C2 => n4444, A => n4206, B => n4205
                           , ZN => n6683);
   U5638 : NOR3_X1 port map( A1 => IF_CPathxmem_en_signal, A2 => n4208, A3 => 
                           n4270, ZN => n4209);
   U5639 : OAI221_X1 port map( B1 => n4209, B2 => n4210, C1 => n4209, C2 => 
                           n4554, A => IF_CPathxsection_0_port, ZN => n4212);
   U5640 : NAND3_X1 port map( A1 => n4549, A2 => n4402, A3 => n4444, ZN => 
                           n4469);
   U5641 : NOR2_X1 port map( A1 => IF_CPathxsection_0_port, A2 => n4275, ZN => 
                           n4555);
   U5642 : NOR2_X1 port map( A1 => n4555, A2 => n6185, ZN => n4448);
   U5643 : OAI221_X1 port map( B1 => n4448, B2 => n4210, C1 => n4448, C2 => 
                           n6196, A => CtlToRegs_port_notify, ZN => n4211);
   U5644 : OAI211_X1 port map( C1 => n4447, C2 => n4212, A => n4469, B => n4211
                           , ZN => n6682);
   U5645 : NOR2_X1 port map( A1 => rst, A2 => n6226, ZN => IF_CPathxN2195);
   U5646 : NOR2_X1 port map( A1 => DecToCtl_port_encType_0_port, A2 => 
                           DecToCtl_port_encType_1_port, ZN => n4213);
   U5647 : OAI221_X1 port map( B1 => n6195, B2 => 
                           DecToCtl_port_instrType_0_port, C1 => n6195, C2 => 
                           n6230, A => n4213, ZN => n4214);
   U5648 : AOI211_X1 port map( C1 => n4214, C2 => n6226, A => 
                           DecToCtl_port_instrType_1_port, B => 
                           DecToCtl_port_instrType_4_port, ZN => n4221);
   U5649 : NAND2_X1 port map( A1 => n4224, A2 => n4254, ZN => n4248);
   U5650 : NOR2_X1 port map( A1 => DecToCtl_port_instrType_2_port, A2 => 
                           DecToCtl_port_instrType_0_port, ZN => n4253);
   U5651 : NAND2_X1 port map( A1 => n4533, A2 => n4253, ZN => n4227);
   U5652 : AOI22_X1 port map( A1 => DecToCtl_port_encType_1_port, A2 => n4248, 
                           B1 => n4227, B2 => n6225, ZN => n4220);
   U5653 : NOR3_X1 port map( A1 => n4225, A2 => DecToCtl_port_encType_1_port, 
                           A3 => DecToCtl_port_instrType_2_port, ZN => n4222);
   U5654 : INV_X1 port map( A => n4222, ZN => n4251);
   U5655 : NAND2_X1 port map( A1 => DecToCtl_port_instrType_4_port, A2 => n4409
                           , ZN => n4461);
   U5656 : NOR2_X1 port map( A1 => n4524, A2 => n6195, ZN => n4215);
   U5657 : OAI211_X1 port map( C1 => DecToCtl_port_instrType_4_port, C2 => 
                           n4532, A => n4215, B => n4543, ZN => n4218);
   U5658 : NOR3_X1 port map( A1 => DecToCtl_port_encType_0_port, A2 => 
                           DecToCtl_port_encType_1_port, A3 => 
                           DecToCtl_port_instrType_2_port, ZN => n4216);
   U5659 : NAND3_X1 port map( A1 => DecToCtl_port_instrType_0_port, A2 => n4216
                           , A3 => n6191, ZN => n4217);
   U5660 : OAI211_X1 port map( C1 => n4251, C2 => n4461, A => n4218, B => n4217
                           , ZN => n4219);
   U5661 : AOI222_X1 port map( A1 => n4221, A2 => n6226, B1 => n4221, B2 => 
                           n4220, C1 => n6226, C2 => n4219, ZN => n4223);
   U5662 : NAND2_X1 port map( A1 => IF_CPathxN2195, A2 => n6191, ZN => n4226);
   U5663 : NAND2_X1 port map( A1 => n4409, A2 => n4222, ZN => n4255);
   U5664 : OAI22_X1 port map( A1 => rst, A2 => n4223, B1 => n4226, B2 => n4255,
                           ZN => n6681);
   U5665 : NOR2_X1 port map( A1 => rst, A2 => n2953, ZN => IF_CPathxN2191);
   U5666 : NOR2_X1 port map( A1 => rst, A2 => n6232, ZN => IF_CPathxN2190);
   U5667 : NAND2_X1 port map( A1 => n4253, A2 => IF_CPathxN2191, ZN => n4240);
   U5668 : NAND3_X1 port map( A1 => n4224, A2 => n4244, A3 => n6191, ZN => 
                           n4538);
   U5669 : NAND4_X1 port map( A1 => n6226, A2 => n6195, A3 => n6189, A4 => 
                           n6191, ZN => n4531);
   U5670 : NOR2_X1 port map( A1 => n4225, A2 => n4531, ZN => n4229);
   U5671 : NAND2_X1 port map( A1 => n6189, A2 => n2953, ZN => n4231);
   U5672 : AOI211_X1 port map( C1 => n4248, C2 => n4227, A => n4226, B => n4231
                           , ZN => n4228);
   U5673 : AOI21_X1 port map( B1 => n4229, B2 => IF_CPathxN2190, A => n4228, ZN
                           => n4239);
   U5674 : AOI211_X1 port map( C1 => n6191, C2 => n2953, A => n6189, B => n4248
                           , ZN => n4237);
   U5675 : NOR2_X1 port map( A1 => DecToCtl_port_instrType_3_port, A2 => n4230,
                           ZN => n4405);
   U5676 : AOI21_X1 port map( B1 => n4267, B2 => n4231, A => 
                           DecToCtl_port_instrType_0_port, ZN => n4232);
   U5677 : AOI22_X1 port map( A1 => n4532, A2 => n4405, B1 => n4533, B2 => 
                           n4232, ZN => n4235);
   U5678 : NAND2_X1 port map( A1 => DecToCtl_port_instrType_2_port, A2 => 
                           DecToCtl_port_instrType_4_port, ZN => n4234);
   U5679 : OAI21_X1 port map( B1 => n4532, B2 => n6197, A => n4242, ZN => n4265
                           );
   U5680 : OAI211_X1 port map( C1 => DecToCtl_port_encType_0_port, C2 => n4528,
                           A => DecToCtl_port_instrType_3_port, B => n6230, ZN 
                           => n4233);
   U5681 : OAI22_X1 port map( A1 => n4235, A2 => n4234, B1 => n4265, B2 => 
                           n4233, ZN => n4236);
   U5682 : OAI211_X1 port map( C1 => n4237, C2 => n4236, A => n4571, B => n6226
                           , ZN => n4238);
   U5683 : OAI211_X1 port map( C1 => n4240, C2 => n4538, A => n4239, B => n4238
                           , ZN => n6680);
   U5684 : NOR2_X1 port map( A1 => DecToCtl_port_instrType_2_port, A2 => n4241,
                           ZN => n4246);
   U5685 : AOI211_X1 port map( C1 => n4242, C2 => n4241, A => rst, B => 
                           DecToCtl_port_encType_0_port, ZN => n4243);
   U5686 : OAI21_X1 port map( B1 => n4244, B2 => n4246, A => n4243, ZN => n4245
                           );
   U5687 : AOI21_X1 port map( B1 => n4246, B2 => n4523, A => n4245, ZN => n6679
                           );
   U5688 : NOR2_X1 port map( A1 => n6226, A2 => n4247, ZN => n4259);
   U5689 : NOR2_X1 port map( A1 => n6225, A2 => n4248, ZN => n4250);
   U5690 : NOR3_X1 port map( A1 => DecToCtl_port_instrType_0_port, A2 => n6195,
                           A3 => n4517, ZN => n4249);
   U5691 : NOR2_X1 port map( A1 => n4250, A2 => n4249, ZN => n4252);
   U5692 : MUX2_X1 port map( A => n4252, B => n4251, S => 
                           DecToCtl_port_instrType_5_port, Z => n4257);
   U5693 : NOR3_X1 port map( A1 => DecToCtl_port_encType_2_port, A2 => 
                           DecToCtl_port_encType_0_port, A3 => 
                           DecToCtl_port_encType_1_port, ZN => n4455);
   U5694 : OAI211_X1 port map( C1 => n4254, C2 => n4253, A => n4455, B => n6226
                           , ZN => n4256);
   U5695 : OAI221_X1 port map( B1 => n2953, B2 => n4257, C1 => 
                           DecToCtl_port_instrType_1_port, C2 => n4256, A => 
                           n4255, ZN => n4258);
   U5696 : AOI21_X1 port map( B1 => n4543, B2 => n4259, A => n4258, ZN => n4260
                           );
   U5697 : NAND2_X1 port map( A1 => n4571, A2 => n6191, ZN => n4411);
   U5698 : NOR2_X1 port map( A1 => n4260, A2 => n4411, ZN => n6678);
   U5699 : NOR2_X1 port map( A1 => rst, A2 => n6195, ZN => IF_CPathxN2192);
   U5700 : AND3_X1 port map( A1 => DecToCtl_port_encType_1_port, A2 => n4261, 
                           A3 => IF_CPathxN2192, ZN => n6677);
   U5701 : NOR2_X1 port map( A1 => rst, A2 => n6189, ZN => IF_CPathxN2193);
   U5702 : OAI221_X1 port map( B1 => DecToCtl_port_encType_0_port, B2 => n4409,
                           C1 => n6197, C2 => DecToCtl_port_encType_1_port, A 
                           => IF_CPathxN2193, ZN => n4264);
   U5703 : OAI211_X1 port map( C1 => n4262, C2 => n6225, A => n4571, B => n6197
                           , ZN => n4263);
   U5704 : OAI21_X1 port map( B1 => n4265, B2 => n4264, A => n4263, ZN => n6676
                           );
   U5705 : AOI211_X1 port map( C1 => n4267, C2 => n4266, A => n6225, B => n4411
                           , ZN => n6675);
   U5706 : OAI22_X1 port map( A1 => n4270, A2 => n6224, B1 => n4268, B2 => 
                           n6329, ZN => n6671);
   U5707 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_0_port, A2 => 
                           n4545, ZN => n4483);
   U5708 : OAI22_X1 port map( A1 => n4275, A2 => n4483, B1 => n6287, B2 => 
                           n4270, ZN => n6641);
   U5709 : INV_X1 port map( A => IF_CPathxN2090, ZN => n4269);
   U5710 : OAI22_X1 port map( A1 => n4275, A2 => n4269, B1 => n6340, B2 => 
                           n4270, ZN => n6640);
   U5711 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_16_port, A2 => 
                           n4671, ZN => n4499);
   U5712 : OAI22_X1 port map( A1 => n4275, A2 => n4499, B1 => n6288, B2 => 
                           n4270, ZN => n6639);
   U5713 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_24_port, A2 => 
                           n4545, ZN => n4507);
   U5714 : OAI22_X1 port map( A1 => n4275, A2 => n4507, B1 => n6289, B2 => 
                           n4270, ZN => n6637);
   U5715 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_28_port, A2 => 
                           n4545, ZN => n4511);
   U5716 : OAI22_X1 port map( A1 => n4275, A2 => n4511, B1 => n6290, B2 => 
                           n4270, ZN => n6635);
   U5717 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_29_port, A2 => 
                           n4671, ZN => n4512);
   U5718 : OAI22_X1 port map( A1 => n4275, A2 => n4512, B1 => n6291, B2 => 
                           n4270, ZN => n6633);
   U5719 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_10_port, A2 => 
                           n4571, ZN => n4493);
   U5720 : OAI22_X1 port map( A1 => n4275, A2 => n4493, B1 => n6292, B2 => 
                           n4270, ZN => n6631);
   U5721 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_26_port, A2 => 
                           n4546, ZN => n4509);
   U5722 : OAI22_X1 port map( A1 => n4275, A2 => n4509, B1 => n6293, B2 => 
                           n4270, ZN => n6629);
   U5723 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_27_port, A2 => 
                           n6178, ZN => n4510);
   U5724 : OAI22_X1 port map( A1 => n4275, A2 => n4510, B1 => n6294, B2 => 
                           n4270, ZN => n6627);
   U5725 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_12_port, A2 => 
                           n6178, ZN => n4495);
   U5726 : OAI22_X1 port map( A1 => n4275, A2 => n4495, B1 => n6295, B2 => 
                           n4270, ZN => n6625);
   U5727 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_20_port, A2 => 
                           n4671, ZN => n4503);
   U5728 : OAI22_X1 port map( A1 => n4275, A2 => n4503, B1 => n6296, B2 => 
                           n4270, ZN => n6623);
   U5729 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_22_port, A2 => 
                           n4545, ZN => n4505);
   U5730 : OAI22_X1 port map( A1 => n4275, A2 => n4505, B1 => n6297, B2 => 
                           n4270, ZN => n6621);
   U5731 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_23_port, A2 => 
                           n6178, ZN => n4506);
   U5732 : OAI22_X1 port map( A1 => n4275, A2 => n4506, B1 => n6298, B2 => 
                           n4270, ZN => n6619);
   U5733 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_8_port, A2 => 
                           n4547, ZN => n4491);
   U5734 : OAI22_X1 port map( A1 => n4275, A2 => n4491, B1 => n6299, B2 => 
                           n4270, ZN => n6617);
   U5735 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_11_port, A2 => 
                           n4545, ZN => n4494);
   U5736 : OAI22_X1 port map( A1 => n4277, A2 => n4494, B1 => n6300, B2 => 
                           n4270, ZN => n6615);
   U5737 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_13_port, A2 => 
                           n4671, ZN => n4496);
   U5738 : OAI22_X1 port map( A1 => n4277, A2 => n4496, B1 => n6301, B2 => 
                           n4276, ZN => n6613);
   U5739 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_15_port, A2 => 
                           n4545, ZN => n4498);
   U5740 : OAI22_X1 port map( A1 => n4275, A2 => n4498, B1 => n6302, B2 => 
                           n4276, ZN => n6611);
   U5741 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_17_port, A2 => 
                           n4546, ZN => n4500);
   U5742 : OAI22_X1 port map( A1 => n4275, A2 => n4500, B1 => n6303, B2 => 
                           n4276, ZN => n6609);
   U5743 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_19_port, A2 => 
                           n4671, ZN => n4502);
   U5744 : OAI22_X1 port map( A1 => n4275, A2 => n4502, B1 => n6304, B2 => 
                           n4276, ZN => n6607);
   U5745 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_21_port, A2 => 
                           n6178, ZN => n4504);
   U5746 : OAI22_X1 port map( A1 => n4275, A2 => n4504, B1 => n6305, B2 => 
                           n4276, ZN => n6605);
   U5747 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_18_port, A2 => 
                           n4546, ZN => n4501);
   U5748 : OAI22_X1 port map( A1 => n4275, A2 => n4501, B1 => n6306, B2 => 
                           n4276, ZN => n6603);
   U5749 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_4_port, A2 => 
                           n4545, ZN => n4487);
   U5750 : OAI22_X1 port map( A1 => n4275, A2 => n4487, B1 => n6307, B2 => 
                           n4276, ZN => n6601);
   U5751 : INV_X1 port map( A => IF_CPathxN2096, ZN => n4271);
   U5752 : OAI22_X1 port map( A1 => n4275, A2 => n4271, B1 => n6341, B2 => 
                           n4276, ZN => n6600);
   U5753 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_14_port, A2 => 
                           n4671, ZN => n4497);
   U5754 : OAI22_X1 port map( A1 => n4275, A2 => n4497, B1 => n6308, B2 => 
                           n4276, ZN => n6599);
   U5755 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_2_port, A2 => 
                           n4546, ZN => n4485);
   U5756 : OAI22_X1 port map( A1 => n4275, A2 => n4485, B1 => n6309, B2 => 
                           n4276, ZN => n6597);
   U5757 : INV_X1 port map( A => IF_CPathxN2094, ZN => n4272);
   U5758 : OAI22_X1 port map( A1 => n4275, A2 => n4272, B1 => n6342, B2 => 
                           n4276, ZN => n6596);
   U5759 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_3_port, A2 => 
                           n4671, ZN => n4486);
   U5760 : OAI22_X1 port map( A1 => n4275, A2 => n4486, B1 => n6310, B2 => 
                           n4276, ZN => n6595);
   U5761 : INV_X1 port map( A => IF_CPathxN2095, ZN => n4273);
   U5762 : OAI22_X1 port map( A1 => n4275, A2 => n4273, B1 => n6343, B2 => 
                           n4276, ZN => n6594);
   U5763 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_1_port, A2 => 
                           n4671, ZN => n4484);
   U5764 : OAI22_X1 port map( A1 => n4275, A2 => n4484, B1 => n6311, B2 => 
                           n4276, ZN => n6593);
   U5765 : INV_X1 port map( A => IF_CPathxN2092, ZN => n4274);
   U5766 : OAI22_X1 port map( A1 => n4275, A2 => n4274, B1 => n6344, B2 => 
                           n4276, ZN => n6592);
   U5767 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_5_port, A2 => 
                           n6178, ZN => n4488);
   U5768 : OAI22_X1 port map( A1 => n4275, A2 => n4488, B1 => n6312, B2 => 
                           n4276, ZN => n6591);
   U5769 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_7_port, A2 => 
                           n6178, ZN => n4490);
   U5770 : OAI22_X1 port map( A1 => n4275, A2 => n4490, B1 => n6313, B2 => 
                           n4276, ZN => n6589);
   U5771 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_25_port, A2 => 
                           n6178, ZN => n4508);
   U5772 : OAI22_X1 port map( A1 => n4275, A2 => n4508, B1 => n6314, B2 => 
                           n4276, ZN => n6587);
   U5773 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_9_port, A2 => 
                           n4671, ZN => n4492);
   U5774 : OAI22_X1 port map( A1 => n4277, A2 => n4492, B1 => n6315, B2 => 
                           n4276, ZN => n6585);
   U5775 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_6_port, A2 => 
                           n4546, ZN => n4489);
   U5776 : OAI22_X1 port map( A1 => n4277, A2 => n4489, B1 => n6316, B2 => 
                           n4276, ZN => n6583);
   U5777 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_30_port, A2 => 
                           n6178, ZN => n4513);
   U5778 : OAI22_X1 port map( A1 => n4277, A2 => n4513, B1 => n6317, B2 => 
                           n4276, ZN => n6581);
   U5779 : NAND2_X1 port map( A1 => RegsToCtl_port_contents2_31_port, A2 => 
                           n4667, ZN => n4514);
   U5780 : OAI22_X1 port map( A1 => n4277, A2 => n4514, B1 => n6318, B2 => 
                           n4276, ZN => n6579);
   U5781 : NOR3_X1 port map( A1 => IF_CPathxwb_sel_signal_1_port, A2 => n4281, 
                           A3 => n6269, ZN => n4362);
   U5782 : INV_X1 port map( A => n4362, ZN => n4383);
   U5783 : INV_X1 port map( A => MemToCtl_port(0), ZN => n4470);
   U5784 : NOR2_X1 port map( A1 => IF_CPathxwb_sel_signal_1_port, A2 => 
                           IF_CPathxwb_sel_signal_0_port, ZN => n4278);
   U5785 : NAND2_X1 port map( A1 => n4279, A2 => n4278, ZN => n4396);
   U5786 : INV_X1 port map( A => n4396, ZN => n4384);
   U5787 : NAND2_X1 port map( A1 => IF_CPathxwb_sel_signal_1_port, A2 => n4671,
                           ZN => n4280);
   U5788 : AOI22_X1 port map( A1 => ALUtoCtl_port_0_port, A2 => n4384, B1 => 
                           n4392, B2 => IF_CPathxpc_reg_signal_0_port, ZN => 
                           n4284);
   U5789 : NOR3_X1 port map( A1 => IF_CPathxwb_sel_signal_1_port, A2 => 
                           IF_CPathxwb_sel_signal_0_port, A3 => n4281, ZN => 
                           n4345);
   U5790 : CLKBUF_X1 port map( A => n4345, Z => n4385);
   U5791 : NOR3_X1 port map( A1 => IF_CPathxwb_sel_signal_1_port, A2 => n4282, 
                           A3 => n6269, ZN => n4369);
   U5792 : CLKBUF_X1 port map( A => n4369, Z => n4391);
   U5793 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_0_port, B1 => n4391, 
                           B2 => IF_CPathxMemToCtl_data_signal_0_port, ZN => 
                           n4283);
   U5794 : OAI211_X1 port map( C1 => n4383, C2 => n4470, A => n4284, B => n4283
                           , ZN => n6578);
   U5795 : AOI22_X1 port map( A1 => n4391, A2 => 
                           IF_CPathxMemToCtl_data_signal_16_port, B1 => n4362, 
                           B2 => MemToCtl_port(16), ZN => n4288);
   U5796 : INV_X1 port map( A => n4285, ZN => n4286);
   U5797 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_16_port, B1 => n4392, 
                           B2 => n4286, ZN => n4287);
   U5798 : OAI211_X1 port map( C1 => n6278, C2 => n4396, A => n4288, B => n4287
                           , ZN => n6577);
   U5799 : INV_X1 port map( A => n4392, ZN => n4388);
   U5800 : CLKBUF_X1 port map( A => n4362, Z => n4390);
   U5801 : AOI22_X1 port map( A1 => ALUtoCtl_port_24_port, A2 => n4384, B1 => 
                           n4390, B2 => MemToCtl_port(24), ZN => n4290);
   U5802 : AOI22_X1 port map( A1 => n4345, A2 => 
                           IF_CPathxALUtoCtl_data_signal_24_port, B1 => n4391, 
                           B2 => IF_CPathxMemToCtl_data_signal_24_port, ZN => 
                           n4289);
   U5803 : OAI211_X1 port map( C1 => n4388, C2 => n4291, A => n4290, B => n4289
                           , ZN => n6576);
   U5804 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_28_port, B1 => n4369, 
                           B2 => IF_CPathxMemToCtl_data_signal_28_port, ZN => 
                           n4295);
   U5805 : INV_X1 port map( A => n4292, ZN => n4293);
   U5806 : AOI22_X1 port map( A1 => n4392, A2 => n4293, B1 => n4390, B2 => 
                           MemToCtl_port(28), ZN => n4294);
   U5807 : OAI211_X1 port map( C1 => n6284, C2 => n4396, A => n4295, B => n4294
                           , ZN => n6575);
   U5808 : AOI22_X1 port map( A1 => n4391, A2 => 
                           IF_CPathxMemToCtl_data_signal_29_port, B1 => n4390, 
                           B2 => MemToCtl_port(29), ZN => n4298);
   U5809 : AOI22_X1 port map( A1 => n4296, A2 => n4392, B1 => n4385, B2 => 
                           IF_CPathxALUtoCtl_data_signal_29_port, ZN => n4297);
   U5810 : OAI211_X1 port map( C1 => n6285, C2 => n4396, A => n4298, B => n4297
                           , ZN => n6574);
   U5811 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_10_port, B1 => n4369, 
                           B2 => IF_CPathxMemToCtl_data_signal_10_port, ZN => 
                           n4302);
   U5812 : INV_X1 port map( A => n4299, ZN => n4300);
   U5813 : AOI22_X1 port map( A1 => n4392, A2 => n4300, B1 => n4390, B2 => 
                           MemToCtl_port(10), ZN => n4301);
   U5814 : OAI211_X1 port map( C1 => n6275, C2 => n4396, A => n4302, B => n4301
                           , ZN => n6573);
   U5815 : AOI22_X1 port map( A1 => ALUtoCtl_port_26_port, A2 => n4384, B1 => 
                           n4390, B2 => MemToCtl_port(26), ZN => n4304);
   U5816 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_26_port, B1 => n4391, 
                           B2 => IF_CPathxMemToCtl_data_signal_26_port, ZN => 
                           n4303);
   U5817 : OAI211_X1 port map( C1 => n4388, C2 => n4305, A => n4304, B => n4303
                           , ZN => n6572);
   U5818 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_27_port, B1 => n4369, 
                           B2 => IF_CPathxMemToCtl_data_signal_27_port, ZN => 
                           n4308);
   U5819 : AOI22_X1 port map( A1 => n4392, A2 => n4306, B1 => n4362, B2 => 
                           MemToCtl_port(27), ZN => n4307);
   U5820 : OAI211_X1 port map( C1 => n6283, C2 => n4396, A => n4308, B => n4307
                           , ZN => n6571);
   U5821 : AOI22_X1 port map( A1 => ALUtoCtl_port_12_port, A2 => n4384, B1 => 
                           n4390, B2 => MemToCtl_port(12), ZN => n4310);
   U5822 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_12_port, B1 => n4369, 
                           B2 => IF_CPathxMemToCtl_data_signal_12_port, ZN => 
                           n4309);
   U5823 : OAI211_X1 port map( C1 => n4388, C2 => n4311, A => n4310, B => n4309
                           , ZN => n6570);
   U5824 : INV_X1 port map( A => MemToCtl_port(20), ZN => n4477);
   U5825 : AOI22_X1 port map( A1 => ALUtoCtl_port_20_port, A2 => n4384, B1 => 
                           n4345, B2 => IF_CPathxALUtoCtl_data_signal_20_port, 
                           ZN => n4315);
   U5826 : INV_X1 port map( A => n4312, ZN => n4313);
   U5827 : AOI22_X1 port map( A1 => n4392, A2 => n4313, B1 => n4369, B2 => 
                           IF_CPathxMemToCtl_data_signal_20_port, ZN => n4314);
   U5828 : OAI211_X1 port map( C1 => n4383, C2 => n4477, A => n4315, B => n4314
                           , ZN => n6569);
   U5829 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_22_port, B1 => n4390, 
                           B2 => MemToCtl_port(22), ZN => n4319);
   U5830 : INV_X1 port map( A => n4316, ZN => n4317);
   U5831 : AOI22_X1 port map( A1 => n4392, A2 => n4317, B1 => n4391, B2 => 
                           IF_CPathxMemToCtl_data_signal_22_port, ZN => n4318);
   U5832 : OAI211_X1 port map( C1 => n6276, C2 => n4396, A => n4319, B => n4318
                           , ZN => n6568);
   U5833 : INV_X1 port map( A => MemToCtl_port(23), ZN => n4479);
   U5834 : AOI22_X1 port map( A1 => ALUtoCtl_port_23_port, A2 => n4384, B1 => 
                           n4345, B2 => IF_CPathxALUtoCtl_data_signal_23_port, 
                           ZN => n4322);
   U5835 : AOI22_X1 port map( A1 => n4392, A2 => n4320, B1 => n4391, B2 => 
                           IF_CPathxMemToCtl_data_signal_23_port, ZN => n4321);
   U5836 : OAI211_X1 port map( C1 => n4383, C2 => n4479, A => n4322, B => n4321
                           , ZN => n6567);
   U5837 : AOI22_X1 port map( A1 => ALUtoCtl_port_8_port, A2 => n4384, B1 => 
                           n4390, B2 => MemToCtl_port(8), ZN => n4324);
   U5838 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_8_port, B1 => n4391, 
                           B2 => IF_CPathxMemToCtl_data_signal_8_port, ZN => 
                           n4323);
   U5839 : OAI211_X1 port map( C1 => n4388, C2 => n4325, A => n4324, B => n4323
                           , ZN => n6566);
   U5840 : INV_X1 port map( A => MemToCtl_port(11), ZN => n4472);
   U5841 : AOI22_X1 port map( A1 => ALUtoCtl_port_11_port, A2 => n4384, B1 => 
                           n4345, B2 => IF_CPathxALUtoCtl_data_signal_11_port, 
                           ZN => n4328);
   U5842 : AOI22_X1 port map( A1 => n4392, A2 => n4326, B1 => n4391, B2 => 
                           IF_CPathxMemToCtl_data_signal_11_port, ZN => n4327);
   U5843 : OAI211_X1 port map( C1 => n4383, C2 => n4472, A => n4328, B => n4327
                           , ZN => n6565);
   U5844 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_13_port, B1 => n4391, 
                           B2 => IF_CPathxMemToCtl_data_signal_13_port, ZN => 
                           n4331);
   U5845 : AOI22_X1 port map( A1 => n4392, A2 => n4329, B1 => n4362, B2 => 
                           MemToCtl_port(13), ZN => n4330);
   U5846 : OAI211_X1 port map( C1 => n6282, C2 => n4396, A => n4331, B => n4330
                           , ZN => n6564);
   U5847 : INV_X1 port map( A => MemToCtl_port(15), ZN => n4474);
   U5848 : AOI22_X1 port map( A1 => ALUtoCtl_port_15_port, A2 => n4384, B1 => 
                           n4345, B2 => IF_CPathxALUtoCtl_data_signal_15_port, 
                           ZN => n4334);
   U5849 : AOI22_X1 port map( A1 => n4392, A2 => n4332, B1 => n4391, B2 => 
                           IF_CPathxMemToCtl_data_signal_15_port, ZN => n4333);
   U5850 : OAI211_X1 port map( C1 => n4383, C2 => n4474, A => n4334, B => n4333
                           , ZN => n6563);
   U5851 : INV_X1 port map( A => MemToCtl_port(17), ZN => n4475);
   U5852 : AOI22_X1 port map( A1 => ALUtoCtl_port_17_port, A2 => n4384, B1 => 
                           n4391, B2 => IF_CPathxMemToCtl_data_signal_17_port, 
                           ZN => n4337);
   U5853 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_17_port, B1 => n4392, 
                           B2 => n4335, ZN => n4336);
   U5854 : OAI211_X1 port map( C1 => n4383, C2 => n4475, A => n4337, B => n4336
                           , ZN => n6562);
   U5855 : INV_X1 port map( A => n4338, ZN => n4341);
   U5856 : AOI22_X1 port map( A1 => ALUtoCtl_port_19_port, A2 => n4384, B1 => 
                           n4390, B2 => MemToCtl_port(19), ZN => n4340);
   U5857 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_19_port, B1 => n4391, 
                           B2 => IF_CPathxMemToCtl_data_signal_19_port, ZN => 
                           n4339);
   U5858 : OAI211_X1 port map( C1 => n4388, C2 => n4341, A => n4340, B => n4339
                           , ZN => n6561);
   U5859 : INV_X1 port map( A => MemToCtl_port(21), ZN => n4478);
   U5860 : AOI22_X1 port map( A1 => ALUtoCtl_port_21_port, A2 => n4384, B1 => 
                           n4345, B2 => IF_CPathxALUtoCtl_data_signal_21_port, 
                           ZN => n4344);
   U5861 : AOI22_X1 port map( A1 => n4392, A2 => n4342, B1 => n4391, B2 => 
                           IF_CPathxMemToCtl_data_signal_21_port, ZN => n4343);
   U5862 : OAI211_X1 port map( C1 => n4383, C2 => n4478, A => n4344, B => n4343
                           , ZN => n6560);
   U5863 : INV_X1 port map( A => MemToCtl_port(18), ZN => n4476);
   U5864 : AOI22_X1 port map( A1 => ALUtoCtl_port_18_port, A2 => n4384, B1 => 
                           n4345, B2 => IF_CPathxALUtoCtl_data_signal_18_port, 
                           ZN => n4349);
   U5865 : INV_X1 port map( A => n4346, ZN => n4347);
   U5866 : AOI22_X1 port map( A1 => n4392, A2 => n4347, B1 => n4391, B2 => 
                           IF_CPathxMemToCtl_data_signal_18_port, ZN => n4348);
   U5867 : OAI211_X1 port map( C1 => n4383, C2 => n4476, A => n4349, B => n4348
                           , ZN => n6559);
   U5868 : AOI22_X1 port map( A1 => ALUtoCtl_port_4_port, A2 => n4384, B1 => 
                           n4390, B2 => MemToCtl_port(4), ZN => n4351);
   U5869 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_4_port, B1 => n4391, 
                           B2 => IF_CPathxMemToCtl_data_signal_4_port, ZN => 
                           n4350);
   U5870 : OAI211_X1 port map( C1 => n4388, C2 => n4352, A => n4351, B => n4350
                           , ZN => n6558);
   U5871 : INV_X1 port map( A => MemToCtl_port(14), ZN => n4473);
   U5872 : AOI22_X1 port map( A1 => ALUtoCtl_port_14_port, A2 => n4384, B1 => 
                           n4391, B2 => IF_CPathxMemToCtl_data_signal_14_port, 
                           ZN => n4356);
   U5873 : INV_X1 port map( A => n4353, ZN => n4354);
   U5874 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_14_port, B1 => n4392, 
                           B2 => n4354, ZN => n4355);
   U5875 : OAI211_X1 port map( C1 => n4383, C2 => n4473, A => n4356, B => n4355
                           , ZN => n6557);
   U5876 : AOI22_X1 port map( A1 => ALUtoCtl_port_2_port, A2 => n4384, B1 => 
                           n4385, B2 => IF_CPathxALUtoCtl_data_signal_2_port, 
                           ZN => n4358);
   U5877 : AOI22_X1 port map( A1 => n4391, A2 => 
                           IF_CPathxMemToCtl_data_signal_2_port, B1 => n4390, 
                           B2 => MemToCtl_port(2), ZN => n4357);
   U5878 : OAI211_X1 port map( C1 => IF_CPathxpc_reg_signal_2_port, C2 => n4388
                           , A => n4358, B => n4357, ZN => n6556);
   U5879 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_3_port, B1 => n4362, 
                           B2 => MemToCtl_port(3), ZN => n4361);
   U5880 : AOI22_X1 port map( A1 => n4392, A2 => n4359, B1 => n4391, B2 => 
                           IF_CPathxMemToCtl_data_signal_3_port, ZN => n4360);
   U5881 : OAI211_X1 port map( C1 => n6277, C2 => n4396, A => n4361, B => n4360
                           , ZN => n6555);
   U5882 : AOI22_X1 port map( A1 => n4391, A2 => 
                           IF_CPathxMemToCtl_data_signal_1_port, B1 => n4362, 
                           B2 => MemToCtl_port(1), ZN => n4364);
   U5883 : AOI22_X1 port map( A1 => ALUtoCtl_port_1_port, A2 => n4384, B1 => 
                           n4385, B2 => IF_CPathxALUtoCtl_data_signal_1_port, 
                           ZN => n4363);
   U5884 : OAI211_X1 port map( C1 => n4388, C2 => n6323, A => n4364, B => n4363
                           , ZN => n6554);
   U5885 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_5_port, B1 => n4391, 
                           B2 => IF_CPathxMemToCtl_data_signal_5_port, ZN => 
                           n4367);
   U5886 : AOI22_X1 port map( A1 => n4392, A2 => n4365, B1 => n4390, B2 => 
                           MemToCtl_port(5), ZN => n4366);
   U5887 : OAI211_X1 port map( C1 => n6280, C2 => n4396, A => n4367, B => n4366
                           , ZN => n6553);
   U5888 : INV_X1 port map( A => n4368, ZN => n4372);
   U5889 : AOI22_X1 port map( A1 => ALUtoCtl_port_7_port, A2 => n4384, B1 => 
                           n4390, B2 => MemToCtl_port(7), ZN => n4371);
   U5890 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_7_port, B1 => n4369, 
                           B2 => IF_CPathxMemToCtl_data_signal_7_port, ZN => 
                           n4370);
   U5891 : OAI211_X1 port map( C1 => n4388, C2 => n4372, A => n4371, B => n4370
                           , ZN => n6552);
   U5892 : INV_X1 port map( A => MemToCtl_port(25), ZN => n4480);
   U5893 : AOI22_X1 port map( A1 => ALUtoCtl_port_25_port, A2 => n4384, B1 => 
                           n4391, B2 => IF_CPathxMemToCtl_data_signal_25_port, 
                           ZN => n4375);
   U5894 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_25_port, B1 => n4392, 
                           B2 => n4373, ZN => n4374);
   U5895 : OAI211_X1 port map( C1 => n4383, C2 => n4480, A => n4375, B => n4374
                           , ZN => n6551);
   U5896 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_9_port, B1 => n4391, 
                           B2 => IF_CPathxMemToCtl_data_signal_9_port, ZN => 
                           n4378);
   U5897 : AOI22_X1 port map( A1 => n4392, A2 => n4376, B1 => n4390, B2 => 
                           MemToCtl_port(9), ZN => n4377);
   U5898 : OAI211_X1 port map( C1 => n6281, C2 => n4396, A => n4378, B => n4377
                           , ZN => n6550);
   U5899 : INV_X1 port map( A => MemToCtl_port(6), ZN => n4471);
   U5900 : AOI22_X1 port map( A1 => ALUtoCtl_port_6_port, A2 => n4384, B1 => 
                           n4391, B2 => IF_CPathxMemToCtl_data_signal_6_port, 
                           ZN => n4382);
   U5901 : INV_X1 port map( A => n4379, ZN => n4380);
   U5902 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_6_port, B1 => n4392, 
                           B2 => n4380, ZN => n4381);
   U5903 : OAI211_X1 port map( C1 => n4383, C2 => n4471, A => n4382, B => n4381
                           , ZN => n6549);
   U5904 : AOI22_X1 port map( A1 => ALUtoCtl_port_30_port, A2 => n4384, B1 => 
                           n4390, B2 => MemToCtl_port(30), ZN => n4387);
   U5905 : AOI22_X1 port map( A1 => n4385, A2 => 
                           IF_CPathxALUtoCtl_data_signal_30_port, B1 => n4391, 
                           B2 => IF_CPathxMemToCtl_data_signal_30_port, ZN => 
                           n4386);
   U5906 : OAI211_X1 port map( C1 => n4389, C2 => n4388, A => n4387, B => n4386
                           , ZN => n6548);
   U5907 : AOI22_X1 port map( A1 => n4391, A2 => 
                           IF_CPathxMemToCtl_data_signal_31_port, B1 => 
                           MemToCtl_port(31), B2 => n4390, ZN => n4395);
   U5908 : AOI22_X1 port map( A1 => n4393, A2 => n4392, B1 => n4385, B2 => 
                           IF_CPathxALUtoCtl_data_signal_31_port, ZN => n4394);
   U5909 : OAI211_X1 port map( C1 => n6279, C2 => n4396, A => n4395, B => n4394
                           , ZN => n6547);
   U5910 : AOI22_X1 port map( A1 => 
                           IF_CPathxDecToCtl_data_signal_rd_addr_0_port, A2 => 
                           n6546, B1 => n4402, B2 => 
                           IF_CPathxCtlToRegs_data_signal_dst_0_port, ZN => 
                           n4397);
   U5911 : INV_X1 port map( A => n4397, ZN => n6545);
   U5912 : AOI22_X1 port map( A1 => 
                           IF_CPathxDecToCtl_data_signal_rd_addr_1_port, A2 => 
                           n6546, B1 => n4402, B2 => 
                           IF_CPathxCtlToRegs_data_signal_dst_1_port, ZN => 
                           n4398);
   U5913 : INV_X1 port map( A => n4398, ZN => n6544);
   U5914 : AOI22_X1 port map( A1 => 
                           IF_CPathxDecToCtl_data_signal_rd_addr_2_port, A2 => 
                           n6546, B1 => n4402, B2 => 
                           IF_CPathxCtlToRegs_data_signal_dst_2_port, ZN => 
                           n4399);
   U5915 : INV_X1 port map( A => n4399, ZN => n6543);
   U5916 : AOI22_X1 port map( A1 => 
                           IF_CPathxDecToCtl_data_signal_rd_addr_3_port, A2 => 
                           n6546, B1 => n4402, B2 => 
                           IF_CPathxCtlToRegs_data_signal_dst_3_port, ZN => 
                           n4400);
   U5917 : INV_X1 port map( A => n4400, ZN => n6542);
   U5918 : AOI22_X1 port map( A1 => 
                           IF_CPathxDecToCtl_data_signal_rd_addr_4_port, A2 => 
                           n6546, B1 => n4402, B2 => 
                           IF_CPathxCtlToRegs_data_signal_dst_4_port, ZN => 
                           n4401);
   U5919 : INV_X1 port map( A => n4401, ZN => n6541);
   U5920 : AND3_X1 port map( A1 => n6195, A2 => DecToCtl_port_instrType_0_port,
                           A3 => n4402, ZN => n6540);
   U5921 : OAI211_X1 port map( C1 => DecToCtl_port_encType_2_port, C2 => 
                           DecToCtl_port_instrType_1_port, A => n4402, B => 
                           DecToCtl_port_instrType_4_port, ZN => n4403);
   U5922 : AOI21_X1 port map( B1 => DecToCtl_port_encType_2_port, B2 => 
                           DecToCtl_port_instrType_1_port, A => n4403, ZN => 
                           n6539);
   U5923 : NAND3_X1 port map( A1 => DecToCtl_port_instrType_2_port, A2 => n6196
                           , A3 => n2953, ZN => n4404);
   U5924 : NAND3_X1 port map( A1 => n4416, A2 => n4571, A3 => n4404, ZN => 
                           n6538);
   U5925 : NOR2_X1 port map( A1 => rst, A2 => n6191, ZN => IF_CPathxN2194);
   U5926 : NAND2_X1 port map( A1 => DecToCtl_port_instrType_2_port, A2 => 
                           DecToCtl_port_instrType_1_port, ZN => n4522);
   U5927 : NAND4_X1 port map( A1 => DecToCtl_port_encType_1_port, A2 => n4405, 
                           A3 => IF_CPathxN2194, A4 => n4522, ZN => n4407);
   U5928 : NAND2_X1 port map( A1 => n4406, A2 => n4407, ZN => n6505);
   U5929 : OAI21_X1 port map( B1 => n4464, B2 => n4455, A => n4667, ZN => n4410
                           );
   U5930 : NAND2_X1 port map( A1 => n4410, A2 => n4407, ZN => n6504);
   U5931 : AOI21_X1 port map( B1 => n4543, B2 => n4409, A => n4408, ZN => n4412
                           );
   U5932 : OAI21_X1 port map( B1 => n4412, B2 => n4411, A => n4410, ZN => n6503
                           );
   U5933 : NOR3_X1 port map( A1 => rst, A2 => DecToCtl_port_encType_2_port, A3 
                           => DecToCtl_port_encType_1_port, ZN => n6502);
   U5934 : AND2_X1 port map( A1 => n4413, A2 => 
                           IF_CPathxmemoryAccess_signal_mask_0_port, ZN => 
                           n6501);
   U5935 : AND2_X1 port map( A1 => n4413, A2 => 
                           IF_CPathxmemoryAccess_signal_mask_1_port, ZN => 
                           n6500);
   U5936 : INV_X1 port map( A => n4415, ZN => n4414);
   U5937 : OR2_X1 port map( A1 => IF_CPathxmemoryAccess_signal_mask_2_port, A2 
                           => n4414, ZN => n6499);
   U5938 : NOR2_X1 port map( A1 => n4414, A2 => n6286, ZN => n6498);
   U5939 : NOR2_X1 port map( A1 => n4414, A2 => n6287, ZN => n6496);
   U5940 : NOR2_X1 port map( A1 => n4414, A2 => n6288, ZN => n6494);
   U5941 : NOR2_X1 port map( A1 => n4414, A2 => n6289, ZN => n6492);
   U5942 : NOR2_X1 port map( A1 => n4414, A2 => n6290, ZN => n6490);
   U5943 : NOR2_X1 port map( A1 => n4414, A2 => n6291, ZN => n6488);
   U5944 : NOR2_X1 port map( A1 => n4414, A2 => n6292, ZN => n6486);
   U5945 : NOR2_X1 port map( A1 => n4414, A2 => n6293, ZN => n6484);
   U5946 : NOR2_X1 port map( A1 => n4414, A2 => n6294, ZN => n6482);
   U5947 : NOR2_X1 port map( A1 => n3251, A2 => n6295, ZN => n6480);
   U5948 : NOR2_X1 port map( A1 => n3251, A2 => n6296, ZN => n6478);
   U5949 : NOR2_X1 port map( A1 => n3251, A2 => n6297, ZN => n6476);
   U5950 : NOR2_X1 port map( A1 => n3251, A2 => n6298, ZN => n6474);
   U5951 : NOR2_X1 port map( A1 => n3251, A2 => n6299, ZN => n6472);
   U5952 : NOR2_X1 port map( A1 => n3251, A2 => n6300, ZN => n6470);
   U5953 : NOR2_X1 port map( A1 => n3251, A2 => n6301, ZN => n6468);
   U5954 : NOR2_X1 port map( A1 => n3251, A2 => n6302, ZN => n6466);
   U5955 : NOR2_X1 port map( A1 => n3251, A2 => n6303, ZN => n6464);
   U5956 : NOR2_X1 port map( A1 => n3251, A2 => n6304, ZN => n6462);
   U5957 : NOR2_X1 port map( A1 => n3251, A2 => n6305, ZN => n6460);
   U5958 : NOR2_X1 port map( A1 => n3251, A2 => n6306, ZN => n6458);
   U5959 : NOR2_X1 port map( A1 => n4414, A2 => n6307, ZN => n6456);
   U5960 : NOR2_X1 port map( A1 => n4414, A2 => n6308, ZN => n6454);
   U5961 : NOR2_X1 port map( A1 => n4414, A2 => n6309, ZN => n6452);
   U5962 : NOR2_X1 port map( A1 => n3251, A2 => n6310, ZN => n6450);
   U5963 : NOR2_X1 port map( A1 => n3251, A2 => n6311, ZN => n6448);
   U5964 : NOR2_X1 port map( A1 => n3251, A2 => n6312, ZN => n6446);
   U5965 : NOR2_X1 port map( A1 => n3251, A2 => n6313, ZN => n6444);
   U5966 : NOR2_X1 port map( A1 => n3251, A2 => n6314, ZN => n6442);
   U5967 : NOR2_X1 port map( A1 => n3251, A2 => n6315, ZN => n6440);
   U5968 : NOR2_X1 port map( A1 => n3251, A2 => n6316, ZN => n6438);
   U5969 : NOR2_X1 port map( A1 => n3251, A2 => n6317, ZN => n6436);
   U5970 : NOR2_X1 port map( A1 => n3251, A2 => n6318, ZN => n6434);
   U5971 : INV_X1 port map( A => n6182, ZN => n4427);
   U5972 : INV_X1 port map( A => n4416, ZN => n4426);
   U5973 : AOI22_X1 port map( A1 => n4427, A2 => DecToCtl_port_rs2_addr_0_port,
                           B1 => IF_CPathxCtlToRegs_data_signal_src2_0_port, B2
                           => n4426, ZN => n4417);
   U5974 : INV_X1 port map( A => n4417, ZN => n6433);
   U5975 : AOI22_X1 port map( A1 => n4427, A2 => DecToCtl_port_rs2_addr_1_port,
                           B1 => IF_CPathxCtlToRegs_data_signal_src2_1_port, B2
                           => n4426, ZN => n4418);
   U5976 : INV_X1 port map( A => n4418, ZN => n6432);
   U5977 : AOI22_X1 port map( A1 => n4427, A2 => DecToCtl_port_rs2_addr_2_port,
                           B1 => IF_CPathxCtlToRegs_data_signal_src2_2_port, B2
                           => n4426, ZN => n4419);
   U5978 : INV_X1 port map( A => n4419, ZN => n6431);
   U5979 : AOI22_X1 port map( A1 => n4427, A2 => DecToCtl_port_rs2_addr_3_port,
                           B1 => IF_CPathxCtlToRegs_data_signal_src2_3_port, B2
                           => n4426, ZN => n4420);
   U5980 : INV_X1 port map( A => n4420, ZN => n6430);
   U5981 : AOI22_X1 port map( A1 => n4427, A2 => DecToCtl_port_rs2_addr_4_port,
                           B1 => IF_CPathxCtlToRegs_data_signal_src2_4_port, B2
                           => n4426, ZN => n4421);
   U5982 : INV_X1 port map( A => n4421, ZN => n6429);
   U5983 : AOI22_X1 port map( A1 => n4427, A2 => DecToCtl_port_rs1_addr_0_port,
                           B1 => IF_CPathxCtlToRegs_data_signal_src1_0_port, B2
                           => n4426, ZN => n4422);
   U5984 : INV_X1 port map( A => n4422, ZN => n6428);
   U5985 : AOI22_X1 port map( A1 => n4427, A2 => DecToCtl_port_rs1_addr_1_port,
                           B1 => IF_CPathxCtlToRegs_data_signal_src1_1_port, B2
                           => n4426, ZN => n4423);
   U5986 : INV_X1 port map( A => n4423, ZN => n6427);
   U5987 : AOI22_X1 port map( A1 => n4427, A2 => DecToCtl_port_rs1_addr_2_port,
                           B1 => IF_CPathxCtlToRegs_data_signal_src1_2_port, B2
                           => n4426, ZN => n4424);
   U5988 : INV_X1 port map( A => n4424, ZN => n6426);
   U5989 : AOI22_X1 port map( A1 => n4427, A2 => DecToCtl_port_rs1_addr_3_port,
                           B1 => IF_CPathxCtlToRegs_data_signal_src1_3_port, B2
                           => n4426, ZN => n4425);
   U5990 : INV_X1 port map( A => n4425, ZN => n6425);
   U5991 : AOI22_X1 port map( A1 => n4427, A2 => DecToCtl_port_rs1_addr_4_port,
                           B1 => IF_CPathxCtlToRegs_data_signal_src1_4_port, B2
                           => n4426, ZN => n4428);
   U5992 : INV_X1 port map( A => n4428, ZN => n6424);
   U5993 : OR2_X1 port map( A1 => rst, A2 => CtlToALU_port_notify, ZN => 
                           IF_ALUxN937);
   U5994 : AOI21_X1 port map( B1 => 
                           IF_CPathxCtlToALU_data_signal_op2_sel_1_port, B2 => 
                           n4430, A => n4429, ZN => n4431);
   U5995 : INV_X1 port map( A => n4431, ZN => IF_CPathxN1668);
   U5996 : INV_X1 port map( A => n4443, ZN => n4452);
   U5997 : AOI211_X1 port map( C1 => n4432, C2 => 
                           IF_CPathxCtlToALU_data_signal_op1_sel_0_port, A => 
                           n4434, B => n4452, ZN => n4433);
   U5998 : AOI22_X1 port map( A1 => n4541, A2 => n4433, B1 => n6345, B2 => 
                           n4521, ZN => IF_CPathxN1664);
   U5999 : NOR2_X1 port map( A1 => n4435, A2 => n4434, ZN => n4518);
   U6000 : OAI21_X1 port map( B1 => n4521, B2 => n4518, A => 
                           IF_CPathxCtlToALU_data_signal_op1_sel_1_port, ZN => 
                           n4436);
   U6001 : OAI21_X1 port map( B1 => n4521, B2 => n4443, A => n4436, ZN => 
                           IF_CPathxN1665);
   U6002 : NAND3_X1 port map( A1 => n4517, A2 => n4438, A3 => n4437, ZN => 
                           n4439);
   U6003 : NAND3_X1 port map( A1 => n4541, A2 => n4440, A3 => n4439, ZN => 
                           n4441);
   U6004 : AND2_X1 port map( A1 => IF_CPathxCtlToALU_data_signal_alu_fun_0_port
                           , A2 => n4441, ZN => IF_CPathxN1628);
   U6005 : AND2_X1 port map( A1 => IF_CPathxCtlToALU_data_signal_alu_fun_2_port
                           , A2 => n4441, ZN => IF_CPathxN1630);
   U6006 : OAI21_X1 port map( B1 => n4521, B2 => n4518, A => 
                           IF_CPathxCtlToALU_data_signal_alu_fun_3_port, ZN => 
                           n4442);
   U6007 : OAI21_X1 port map( B1 => n4521, B2 => n4443, A => n4442, ZN => 
                           IF_CPathxN1631);
   U6008 : NOR2_X1 port map( A1 => n4444, A2 => n4521, ZN => n4550);
   U6009 : AND3_X1 port map( A1 => n6227, A2 => IF_CPathxsection_0_port, A3 => 
                           n4445, ZN => n4468);
   U6010 : NOR2_X1 port map( A1 => n4550, A2 => n4468, ZN => n4515);
   U6011 : NOR2_X1 port map( A1 => rst, A2 => n4515, ZN => IF_CPathxN2396);
   U6012 : NAND2_X1 port map( A1 => n4446, A2 => MemToCtl_port_sync, ZN => 
                           n4559);
   U6013 : NOR2_X1 port map( A1 => n6228, A2 => n4559, ZN => n4467);
   U6014 : AOI21_X1 port map( B1 => n4548, B2 => n6199, A => n4467, ZN => n4450
                           );
   U6015 : NOR2_X1 port map( A1 => n4450, A2 => n4447, ZN => n4481);
   U6016 : INV_X1 port map( A => n4481, ZN => n4482);
   U6017 : OAI21_X1 port map( B1 => rst, B2 => n4482, A => n4469, ZN => 
                           IF_CPathxN2394);
   U6018 : INV_X1 port map( A => n4448, ZN => n4449);
   U6019 : NOR2_X1 port map( A1 => n4559, A2 => n4449, ZN => IF_CPathxN2393);
   U6020 : OAI21_X1 port map( B1 => n4451, B2 => n4450, A => n4561, ZN => 
                           IF_CPathxN2274);
   U6021 : INV_X1 port map( A => IF_CPathxN2274, ZN => n4465);
   U6022 : NAND2_X1 port map( A1 => n4465, A2 => n4556, ZN => IF_CPathxN2316);
   U6023 : NOR2_X1 port map( A1 => n4464, A2 => n4452, ZN => n4519);
   U6024 : AOI21_X1 port map( B1 => n4453, B2 => n4541, A => rst, ZN => n4520);
   U6025 : OAI221_X1 port map( B1 => n4521, B2 => n4519, C1 => n4521, C2 => 
                           n4454, A => n4520, ZN => IF_CPathxN2310);
   U6026 : NOR3_X1 port map( A1 => rst, A2 => n4464, A3 => n4455, ZN => 
                           IF_CPathxN2309);
   U6027 : OAI21_X1 port map( B1 => n4456, B2 => n4464, A => n4667, ZN => n4516
                           );
   U6028 : INV_X1 port map( A => n4516, ZN => IF_CPathxN2308);
   U6029 : OAI211_X1 port map( C1 => DecToCtl_port_instrType_2_port, C2 => 
                           n4458, A => n4528, B => n4457, ZN => n4459);
   U6030 : OAI21_X1 port map( B1 => n4461, B2 => n4460, A => n4459, ZN => n4463
                           );
   U6031 : AOI21_X1 port map( B1 => n4464, B2 => n4463, A => n4462, ZN => n4466
                           );
   U6032 : OAI21_X1 port map( B1 => n4466, B2 => n4521, A => n4465, ZN => 
                           IF_CPathxN2235);
   U6033 : OR2_X1 port map( A1 => rst, A2 => n4467, ZN => IF_CPathxN2201);
   U6034 : AND2_X1 port map( A1 => DecToCtl_port_rd_addr_0_port, A2 => n6180, 
                           ZN => IF_CPathxN2196);
   U6035 : AND2_X1 port map( A1 => DecToCtl_port_rd_addr_1_port, A2 => n6180, 
                           ZN => IF_CPathxN2197);
   U6036 : AND2_X1 port map( A1 => DecToCtl_port_rd_addr_2_port, A2 => n6180, 
                           ZN => IF_CPathxN2198);
   U6037 : AND2_X1 port map( A1 => DecToCtl_port_rd_addr_3_port, A2 => n6180, 
                           ZN => IF_CPathxN2199);
   U6038 : AND2_X1 port map( A1 => DecToCtl_port_rd_addr_4_port, A2 => n6180, 
                           ZN => IF_CPathxN2200);
   U6039 : NAND2_X1 port map( A1 => n4571, A2 => n4521, ZN => IF_CPathxN2157);
   U6040 : OR2_X1 port map( A1 => rst, A2 => n4468, ZN => IF_CPathxN2091);
   U6041 : AND2_X1 port map( A1 => DecToCtl_port_rs2_addr_0_port, A2 => n6180, 
                           ZN => IF_CPathxN2084);
   U6042 : AND2_X1 port map( A1 => DecToCtl_port_rs2_addr_1_port, A2 => n4571, 
                           ZN => IF_CPathxN2085);
   U6043 : AND2_X1 port map( A1 => DecToCtl_port_rs2_addr_2_port, A2 => n4571, 
                           ZN => IF_CPathxN2086);
   U6044 : AND2_X1 port map( A1 => DecToCtl_port_rs2_addr_3_port, A2 => n6180, 
                           ZN => IF_CPathxN2087);
   U6045 : AND2_X1 port map( A1 => DecToCtl_port_rs2_addr_4_port, A2 => n6180, 
                           ZN => IF_CPathxN2088);
   U6046 : AND2_X1 port map( A1 => DecToCtl_port_rs1_addr_0_port, A2 => n4571, 
                           ZN => IF_CPathxN2079);
   U6047 : AND2_X1 port map( A1 => DecToCtl_port_rs1_addr_1_port, A2 => n6180, 
                           ZN => IF_CPathxN2080);
   U6048 : AND2_X1 port map( A1 => DecToCtl_port_rs1_addr_2_port, A2 => n6180, 
                           ZN => IF_CPathxN2081);
   U6049 : AND2_X1 port map( A1 => DecToCtl_port_rs1_addr_3_port, A2 => n4571, 
                           ZN => IF_CPathxN2082);
   U6050 : AND2_X1 port map( A1 => DecToCtl_port_rs1_addr_4_port, A2 => n4571, 
                           ZN => IF_CPathxN2083);
   U6051 : NAND2_X1 port map( A1 => n4571, A2 => n4469, ZN => IF_CPathxN2078);
   U6052 : NOR2_X1 port map( A1 => rst, A2 => n4470, ZN => IF_CPathxN2202);
   U6053 : AND2_X1 port map( A1 => n4667, A2 => MemToCtl_port(1), ZN => 
                           IF_CPathxN2203);
   U6054 : AND2_X1 port map( A1 => n4547, A2 => MemToCtl_port(2), ZN => 
                           IF_CPathxN2204);
   U6055 : AND2_X1 port map( A1 => n4547, A2 => MemToCtl_port(3), ZN => 
                           IF_CPathxN2205);
   U6056 : AND2_X1 port map( A1 => n6178, A2 => MemToCtl_port(4), ZN => 
                           IF_CPathxN2206);
   U6057 : AND2_X1 port map( A1 => n4547, A2 => MemToCtl_port(5), ZN => 
                           IF_CPathxN2207);
   U6058 : NOR2_X1 port map( A1 => rst, A2 => n4471, ZN => IF_CPathxN2208);
   U6059 : AND2_X1 port map( A1 => n4547, A2 => MemToCtl_port(7), ZN => 
                           IF_CPathxN2209);
   U6060 : AND2_X1 port map( A1 => n4546, A2 => MemToCtl_port(8), ZN => 
                           IF_CPathxN2210);
   U6061 : AND2_X1 port map( A1 => n4547, A2 => MemToCtl_port(9), ZN => 
                           IF_CPathxN2211);
   U6062 : AND2_X1 port map( A1 => n4547, A2 => MemToCtl_port(10), ZN => 
                           IF_CPathxN2212);
   U6063 : NOR2_X1 port map( A1 => rst, A2 => n4472, ZN => IF_CPathxN2213);
   U6064 : AND2_X1 port map( A1 => n4545, A2 => MemToCtl_port(12), ZN => 
                           IF_CPathxN2214);
   U6065 : AND2_X1 port map( A1 => n4547, A2 => MemToCtl_port(13), ZN => 
                           IF_CPathxN2215);
   U6066 : NOR2_X1 port map( A1 => rst, A2 => n4473, ZN => IF_CPathxN2216);
   U6067 : NOR2_X1 port map( A1 => rst, A2 => n4474, ZN => IF_CPathxN2217);
   U6068 : AND2_X1 port map( A1 => n4547, A2 => MemToCtl_port(16), ZN => 
                           IF_CPathxN2218);
   U6069 : NOR2_X1 port map( A1 => rst, A2 => n4475, ZN => IF_CPathxN2219);
   U6070 : NOR2_X1 port map( A1 => rst, A2 => n4476, ZN => IF_CPathxN2220);
   U6071 : AND2_X1 port map( A1 => n6180, A2 => MemToCtl_port(19), ZN => 
                           IF_CPathxN2221);
   U6072 : NOR2_X1 port map( A1 => rst, A2 => n4477, ZN => IF_CPathxN2222);
   U6073 : NOR2_X1 port map( A1 => rst, A2 => n4478, ZN => IF_CPathxN2223);
   U6074 : AND2_X1 port map( A1 => n4547, A2 => MemToCtl_port(22), ZN => 
                           IF_CPathxN2224);
   U6075 : NOR2_X1 port map( A1 => rst, A2 => n4479, ZN => IF_CPathxN2225);
   U6076 : AND2_X1 port map( A1 => n4571, A2 => MemToCtl_port(24), ZN => 
                           IF_CPathxN2226);
   U6077 : NOR2_X1 port map( A1 => rst, A2 => n4480, ZN => IF_CPathxN2227);
   U6078 : AND2_X1 port map( A1 => n6178, A2 => MemToCtl_port(26), ZN => 
                           IF_CPathxN2228);
   U6079 : AND2_X1 port map( A1 => n4545, A2 => MemToCtl_port(27), ZN => 
                           IF_CPathxN2229);
   U6080 : AND2_X1 port map( A1 => n4547, A2 => MemToCtl_port(28), ZN => 
                           IF_CPathxN2230);
   U6081 : AND2_X1 port map( A1 => n4671, A2 => MemToCtl_port(29), ZN => 
                           IF_CPathxN2231);
   U6082 : AND2_X1 port map( A1 => n4547, A2 => MemToCtl_port(30), ZN => 
                           IF_CPathxN2232);
   U6083 : AND2_X1 port map( A1 => n4547, A2 => MemToCtl_port(31), ZN => 
                           IF_CPathxN2233);
   U6084 : OAI221_X1 port map( B1 => n4482, B2 => IF_CPathxwb_sel_signal_0_port
                           , C1 => n4482, C2 => IF_CPathxwb_sel_signal_1_port, 
                           A => n4546, ZN => IF_CPathxN2044);
   U6085 : OR2_X1 port map( A1 => n4481, A2 => IF_CPathxN2078, ZN => 
                           IF_CPathxN2038);
   U6086 : NOR2_X1 port map( A1 => rst, A2 => n6236, ZN => IF_CPathxN2033);
   U6087 : NOR2_X1 port map( A1 => rst, A2 => n6200, ZN => IF_CPathxN2034);
   U6088 : NOR2_X1 port map( A1 => rst, A2 => n6192, ZN => IF_CPathxN2035);
   U6089 : NOR2_X1 port map( A1 => rst, A2 => n6190, ZN => IF_CPathxN2036);
   U6090 : AND2_X1 port map( A1 => n4571, A2 => 
                           IF_CPathxDecToCtl_data_signal_rd_addr_4_port, ZN => 
                           IF_CPathxN2037);
   U6091 : NAND2_X1 port map( A1 => n4571, A2 => n4482, ZN => IF_CPathxN2032);
   U6092 : INV_X1 port map( A => n4483, ZN => IF_CPathxN2124);
   U6093 : INV_X1 port map( A => n4484, ZN => IF_CPathxN2125);
   U6094 : INV_X1 port map( A => n4485, ZN => IF_CPathxN2126);
   U6095 : INV_X1 port map( A => n4486, ZN => IF_CPathxN2127);
   U6096 : INV_X1 port map( A => n4487, ZN => IF_CPathxN2128);
   U6097 : INV_X1 port map( A => n4488, ZN => IF_CPathxN2129);
   U6098 : INV_X1 port map( A => n4489, ZN => IF_CPathxN2130);
   U6099 : INV_X1 port map( A => n4490, ZN => IF_CPathxN2131);
   U6100 : INV_X1 port map( A => n4491, ZN => IF_CPathxN2132);
   U6101 : INV_X1 port map( A => n4492, ZN => IF_CPathxN2133);
   U6102 : INV_X1 port map( A => n4493, ZN => IF_CPathxN2134);
   U6103 : INV_X1 port map( A => n4494, ZN => IF_CPathxN2135);
   U6104 : INV_X1 port map( A => n4495, ZN => IF_CPathxN2136);
   U6105 : INV_X1 port map( A => n4496, ZN => IF_CPathxN2137);
   U6106 : INV_X1 port map( A => n4497, ZN => IF_CPathxN2138);
   U6107 : INV_X1 port map( A => n4498, ZN => IF_CPathxN2139);
   U6108 : INV_X1 port map( A => n4499, ZN => IF_CPathxN2140);
   U6109 : INV_X1 port map( A => n4500, ZN => IF_CPathxN2141);
   U6110 : INV_X1 port map( A => n4501, ZN => IF_CPathxN2142);
   U6111 : INV_X1 port map( A => n4502, ZN => IF_CPathxN2143);
   U6112 : INV_X1 port map( A => n4503, ZN => IF_CPathxN2144);
   U6113 : INV_X1 port map( A => n4504, ZN => IF_CPathxN2145);
   U6114 : INV_X1 port map( A => n4505, ZN => IF_CPathxN2146);
   U6115 : INV_X1 port map( A => n4506, ZN => IF_CPathxN2147);
   U6116 : INV_X1 port map( A => n4507, ZN => IF_CPathxN2148);
   U6117 : INV_X1 port map( A => n4508, ZN => IF_CPathxN2149);
   U6118 : INV_X1 port map( A => n4509, ZN => IF_CPathxN2150);
   U6119 : INV_X1 port map( A => n4510, ZN => IF_CPathxN2151);
   U6120 : INV_X1 port map( A => n4511, ZN => IF_CPathxN2152);
   U6121 : INV_X1 port map( A => n4512, ZN => IF_CPathxN2153);
   U6122 : INV_X1 port map( A => n4513, ZN => IF_CPathxN2154);
   U6123 : INV_X1 port map( A => n4514, ZN => IF_CPathxN2155);
   U6124 : NAND2_X1 port map( A1 => n4515, A2 => n4546, ZN => IF_CPathxN1935);
   U6125 : OAI21_X1 port map( B1 => rst, B2 => n4517, A => n4516, ZN => 
                           IF_CPathxN1932);
   U6126 : AND2_X1 port map( A1 => n4519, A2 => n4518, ZN => n4537);
   U6127 : OAI21_X1 port map( B1 => n4537, B2 => n4521, A => n4520, ZN => 
                           IF_CPathxN1930);
   U6128 : INV_X1 port map( A => n4522, ZN => n4539);
   U6129 : NOR3_X1 port map( A1 => DecToCtl_port_instrType_2_port, A2 => n4524,
                           A3 => n4523, ZN => n4535);
   U6130 : OAI21_X1 port map( B1 => DecToCtl_port_instrType_0_port, B2 => n4526
                           , A => n4525, ZN => n4529);
   U6131 : AOI22_X1 port map( A1 => DecToCtl_port_instrType_1_port, A2 => n4529
                           , B1 => n4528, B2 => n4527, ZN => n4530);
   U6132 : OAI21_X1 port map( B1 => n4532, B2 => n4531, A => n4530, ZN => n4534
                           );
   U6133 : OAI211_X1 port map( C1 => n4535, C2 => n4534, A => n4533, B => n6225
                           , ZN => n4536);
   U6134 : OAI211_X1 port map( C1 => n4539, C2 => n4538, A => n4537, B => n4536
                           , ZN => n4542);
   U6135 : OAI211_X1 port map( C1 => n4543, C2 => n4542, A => n4541, B => n4540
                           , ZN => n4544);
   U6136 : NAND2_X1 port map( A1 => n4571, A2 => n4544, ZN => IF_CPathxN1892);
   U6137 : NOR2_X1 port map( A1 => rst, A2 => n6238, ZN => IF_CPathxN1860);
   U6138 : AND2_X1 port map( A1 => n4546, A2 => ALUtoCtl_port_1_port, ZN => 
                           IF_CPathxN1861);
   U6139 : AND2_X1 port map( A1 => n4547, A2 => ALUtoCtl_port_2_port, ZN => 
                           IF_CPathxN1862);
   U6140 : NOR2_X1 port map( A1 => rst, A2 => n6277, ZN => IF_CPathxN1863);
   U6141 : AND2_X1 port map( A1 => n4546, A2 => ALUtoCtl_port_4_port, ZN => 
                           IF_CPathxN1864);
   U6142 : NOR2_X1 port map( A1 => rst, A2 => n6280, ZN => IF_CPathxN1865);
   U6143 : AND2_X1 port map( A1 => n4547, A2 => ALUtoCtl_port_6_port, ZN => 
                           IF_CPathxN1866);
   U6144 : AND2_X1 port map( A1 => n4571, A2 => ALUtoCtl_port_7_port, ZN => 
                           IF_CPathxN1867);
   U6145 : AND2_X1 port map( A1 => n4671, A2 => ALUtoCtl_port_8_port, ZN => 
                           IF_CPathxN1868);
   U6146 : NOR2_X1 port map( A1 => rst, A2 => n6281, ZN => IF_CPathxN1869);
   U6147 : NOR2_X1 port map( A1 => rst, A2 => n6275, ZN => IF_CPathxN1870);
   U6148 : AND2_X1 port map( A1 => n4667, A2 => ALUtoCtl_port_11_port, ZN => 
                           IF_CPathxN1871);
   U6149 : AND2_X1 port map( A1 => n6180, A2 => ALUtoCtl_port_12_port, ZN => 
                           IF_CPathxN1872);
   U6150 : NOR2_X1 port map( A1 => rst, A2 => n6282, ZN => IF_CPathxN1873);
   U6151 : AND2_X1 port map( A1 => n6180, A2 => ALUtoCtl_port_14_port, ZN => 
                           IF_CPathxN1874);
   U6152 : AND2_X1 port map( A1 => n4547, A2 => ALUtoCtl_port_15_port, ZN => 
                           IF_CPathxN1875);
   U6153 : NOR2_X1 port map( A1 => rst, A2 => n6278, ZN => IF_CPathxN1876);
   U6154 : AND2_X1 port map( A1 => n4547, A2 => ALUtoCtl_port_17_port, ZN => 
                           IF_CPathxN1877);
   U6155 : AND2_X1 port map( A1 => n6178, A2 => ALUtoCtl_port_18_port, ZN => 
                           IF_CPathxN1878);
   U6156 : AND2_X1 port map( A1 => n4667, A2 => ALUtoCtl_port_19_port, ZN => 
                           IF_CPathxN1879);
   U6157 : AND2_X1 port map( A1 => n4545, A2 => ALUtoCtl_port_20_port, ZN => 
                           IF_CPathxN1880);
   U6158 : AND2_X1 port map( A1 => n4667, A2 => ALUtoCtl_port_21_port, ZN => 
                           IF_CPathxN1881);
   U6159 : NOR2_X1 port map( A1 => rst, A2 => n6276, ZN => IF_CPathxN1882);
   U6160 : AND2_X1 port map( A1 => n4546, A2 => ALUtoCtl_port_23_port, ZN => 
                           IF_CPathxN1883);
   U6161 : AND2_X1 port map( A1 => n6180, A2 => ALUtoCtl_port_24_port, ZN => 
                           IF_CPathxN1884);
   U6162 : AND2_X1 port map( A1 => n4547, A2 => ALUtoCtl_port_25_port, ZN => 
                           IF_CPathxN1885);
   U6163 : AND2_X1 port map( A1 => n4671, A2 => ALUtoCtl_port_26_port, ZN => 
                           IF_CPathxN1886);
   U6164 : NOR2_X1 port map( A1 => rst, A2 => n6283, ZN => IF_CPathxN1887);
   U6165 : NOR2_X1 port map( A1 => rst, A2 => n6284, ZN => IF_CPathxN1888);
   U6166 : NOR2_X1 port map( A1 => rst, A2 => n6285, ZN => IF_CPathxN1889);
   U6167 : AND2_X1 port map( A1 => n6178, A2 => ALUtoCtl_port_30_port, ZN => 
                           IF_CPathxN1890);
   U6168 : NOR2_X1 port map( A1 => rst, A2 => n6279, ZN => IF_CPathxN1891);
   U6169 : OR2_X1 port map( A1 => rst, A2 => n4548, ZN => IF_CPathxN1859);
   U6170 : NOR2_X1 port map( A1 => n4549, A2 => n4555, ZN => n6179);
   U6171 : AOI21_X1 port map( B1 => n6179, B2 => n6228, A => n4550, ZN => n4552
                           );
   U6172 : OAI21_X1 port map( B1 => n4446, B2 => n6199, A => n4553, ZN => n4551
                           );
   U6173 : AOI21_X1 port map( B1 => n4552, B2 => n4551, A => rst, ZN => 
                           IF_CPathxN1856);
   U6174 : AOI21_X1 port map( B1 => n4555, B2 => n4554, A => n4553, ZN => n4557
                           );
   U6175 : AOI21_X1 port map( B1 => n4557, B2 => n4556, A => rst, ZN => 
                           IF_CPathxN1858);
   U6176 : AOI21_X1 port map( B1 => n6186, B2 => CtlToMem_port_sync, A => n4558
                           , ZN => n4560);
   U6177 : NAND3_X1 port map( A1 => n4561, A2 => n4560, A3 => n4559, ZN => 
                           IF_CPathxN1854);
   U6178 : NOR2_X1 port map( A1 => rst, A2 => CtlToDec_port_notify, ZN => n4643
                           );
   U6179 : INV_X1 port map( A => n4643, ZN => IF_DecoderxN596);
   U6180 : NAND3_X1 port map( A1 => CtlToDec_port_0_port, A2 => 
                           CtlToDec_port_1_port, A3 => n6231, ZN => n4566);
   U6181 : OR2_X1 port map( A1 => CtlToDec_port_6_port, A2 => n4566, ZN => 
                           n4649);
   U6182 : NOR2_X1 port map( A1 => n4649, A2 => n6234, ZN => n4576);
   U6183 : INV_X1 port map( A => n4576, ZN => n4654);
   U6184 : NOR2_X1 port map( A1 => CtlToDec_port_2_port, A2 => n4654, ZN => 
                           n4585);
   U6185 : NAND2_X1 port map( A1 => CtlToDec_port_5_port, A2 => n4585, ZN => 
                           n4608);
   U6186 : NOR2_X1 port map( A1 => n6208, A2 => CtlToDec_port_14_port, ZN => 
                           n4624);
   U6187 : NAND2_X1 port map( A1 => n6259, A2 => n4624, ZN => n4602);
   U6188 : INV_X1 port map( A => n4602, ZN => n4635);
   U6189 : NOR2_X1 port map( A1 => CtlToDec_port_2_port, A2 => n4649, ZN => 
                           n4563);
   U6190 : NAND2_X1 port map( A1 => n4563, A2 => n6234, ZN => n4618);
   U6191 : NOR2_X1 port map( A1 => CtlToDec_port_5_port, A2 => n4618, ZN => 
                           n4574);
   U6192 : OAI21_X1 port map( B1 => n4628, B2 => n4635, A => n4574, ZN => n4616
                           );
   U6193 : OAI21_X1 port map( B1 => CtlToDec_port_12_port, B2 => n4608, A => 
                           n4616, ZN => n4570);
   U6194 : NOR2_X1 port map( A1 => n4654, A2 => n6229, ZN => n4634);
   U6195 : INV_X1 port map( A => n4634, ZN => n4596);
   U6196 : NOR2_X1 port map( A1 => CtlToDec_port_12_port, A2 => n4617, ZN => 
                           n4577);
   U6197 : NAND2_X1 port map( A1 => n4563, A2 => n4562, ZN => n4653);
   U6198 : INV_X1 port map( A => n4653, ZN => n4642);
   U6199 : NAND2_X1 port map( A1 => n4577, A2 => n4642, ZN => n4598);
   U6200 : OAI21_X1 port map( B1 => CtlToDec_port_5_port, B2 => n4596, A => 
                           n4598, ZN => n4569);
   U6201 : NOR2_X1 port map( A1 => n4582, A2 => n6260, ZN => n4592);
   U6202 : NAND2_X1 port map( A1 => n4577, A2 => n4592, ZN => n4629);
   U6203 : INV_X1 port map( A => n4566, ZN => n4564);
   U6204 : NAND2_X1 port map( A1 => n4564, A2 => n4595, ZN => n4645);
   U6205 : NOR3_X1 port map( A1 => CtlToDec_port_2_port, A2 => n4566, A3 => 
                           n4565, ZN => n4587);
   U6206 : OAI211_X1 port map( C1 => CtlToDec_port_14_port, C2 => 
                           CtlToDec_port_12_port, A => n4587, B => n6208, ZN =>
                           n4567);
   U6207 : OAI211_X1 port map( C1 => n4629, C2 => n4608, A => n4645, B => n4567
                           , ZN => n4568);
   U6208 : AOI211_X1 port map( C1 => n4617, C2 => n4570, A => n4569, B => n4568
                           , ZN => n4573);
   U6209 : NOR2_X1 port map( A1 => n4654, A2 => n4648, ZN => n4633);
   U6210 : INV_X1 port map( A => n4633, ZN => n4625);
   U6211 : NAND2_X1 port map( A1 => n4571, A2 => n4625, ZN => n4652);
   U6212 : NOR2_X1 port map( A1 => CtlToDec_port_14_port, A2 => n6259, ZN => 
                           n4623);
   U6213 : AOI221_X1 port map( B1 => n4578, B2 => n6208, C1 => n6259, C2 => 
                           n6208, A => n4623, ZN => n4572);
   U6214 : OAI22_X1 port map( A1 => n4573, A2 => n4652, B1 => n4572, B2 => 
                           n4625, ZN => IF_DecoderxN585);
   U6215 : NOR2_X1 port map( A1 => n6208, A2 => n6261, ZN => n4586);
   U6216 : INV_X1 port map( A => n4574, ZN => n4597);
   U6217 : NOR3_X1 port map( A1 => CtlToDec_port_12_port, A2 => n4586, A3 => 
                           n4597, ZN => n4575);
   U6218 : AOI211_X1 port map( C1 => CtlToDec_port_5_port, C2 => n4576, A => 
                           n4587, B => n4575, ZN => n4581);
   U6219 : OAI21_X1 port map( B1 => n4635, B2 => n4613, A => n4642, ZN => n4580
                           );
   U6220 : NOR2_X1 port map( A1 => n6260, A2 => n4638, ZN => n4622);
   U6221 : NOR3_X1 port map( A1 => n4586, A2 => n4622, A3 => n4608, ZN => n4579
                           );
   U6222 : NAND3_X1 port map( A1 => n4578, A2 => n4577, A3 => n6260, ZN => 
                           n4593);
   U6223 : AOI22_X1 port map( A1 => n4581, A2 => n4580, B1 => n4579, B2 => 
                           n4593, ZN => n4591);
   U6224 : NOR2_X1 port map( A1 => CtlToDec_port_30_port, A2 => n4582, ZN => 
                           n4583);
   U6225 : OAI21_X1 port map( B1 => n4583, B2 => n6259, A => n4628, ZN => n4584
                           );
   U6226 : NAND3_X1 port map( A1 => n4633, A2 => CtlToDec_port_14_port, A3 => 
                           n4584, ZN => n4590);
   U6227 : NOR2_X1 port map( A1 => rst, A2 => n4585, ZN => n4647);
   U6228 : AND2_X1 port map( A1 => n6259, A2 => n4586, ZN => n4621);
   U6229 : INV_X1 port map( A => n4587, ZN => n4611);
   U6230 : NOR2_X1 port map( A1 => n4621, A2 => n4611, ZN => n4601);
   U6231 : NAND2_X1 port map( A1 => n4628, A2 => CtlToDec_port_12_port, ZN => 
                           n4588);
   U6232 : NAND4_X1 port map( A1 => n4647, A2 => n4601, A3 => n4617, A4 => 
                           n4588, ZN => n4589);
   U6233 : OAI211_X1 port map( C1 => n4591, C2 => n4652, A => n4590, B => n4589
                           , ZN => IF_DecoderxN586);
   U6234 : AOI211_X1 port map( C1 => CtlToDec_port_14_port, C2 => n4592, A => 
                           CtlToDec_port_13_port, B => n6259, ZN => n4607);
   U6235 : NOR2_X1 port map( A1 => rst, A2 => n4608, ZN => n4630);
   U6236 : INV_X1 port map( A => n4624, ZN => n4594);
   U6237 : OAI21_X1 port map( B1 => n4594, B2 => n6259, A => n4593, ZN => n4600
                           );
   U6238 : NAND3_X1 port map( A1 => CtlToDec_port_0_port, A2 => 
                           CtlToDec_port_1_port, A3 => n4595, ZN => n4610);
   U6239 : AND2_X1 port map( A1 => n4596, A2 => n4610, ZN => n4651);
   U6240 : NAND3_X1 port map( A1 => n4647, A2 => n4597, A3 => n4611, ZN => 
                           n4641);
   U6241 : AOI21_X1 port map( B1 => n4651, B2 => n4598, A => n4641, ZN => n4599
                           );
   U6242 : AOI21_X1 port map( B1 => n4630, B2 => n4600, A => n4599, ZN => n4606
                           );
   U6243 : INV_X1 port map( A => n4601, ZN => n4604);
   U6244 : OAI21_X1 port map( B1 => n4602, B2 => n4618, A => n4611, ZN => n4603
                           );
   U6245 : OAI211_X1 port map( C1 => n4613, C2 => n4604, A => n4647, B => n4603
                           , ZN => n4605);
   U6246 : OAI211_X1 port map( C1 => n4607, C2 => n4625, A => n4606, B => n4605
                           , ZN => IF_DecoderxN587);
   U6247 : NOR3_X1 port map( A1 => n4624, A2 => n4623, A3 => n4622, ZN => n4615
                           );
   U6248 : NOR2_X1 port map( A1 => n4624, A2 => n4623, ZN => n4609);
   U6249 : NOR2_X1 port map( A1 => n4609, A2 => n4608, ZN => n4620);
   U6250 : OAI21_X1 port map( B1 => n4624, B2 => n4611, A => n4610, ZN => n4612
                           );
   U6251 : AOI211_X1 port map( C1 => n4613, C2 => n4642, A => n4620, B => n4612
                           , ZN => n4614);
   U6252 : OAI22_X1 port map( A1 => n4615, A2 => n4625, B1 => n4614, B2 => 
                           n4652, ZN => IF_DecoderxN588);
   U6253 : OAI21_X1 port map( B1 => n4618, B2 => n4617, A => n4616, ZN => n4619
                           );
   U6254 : AOI211_X1 port map( C1 => n4634, C2 => CtlToDec_port_5_port, A => 
                           n4620, B => n4619, ZN => n4627);
   U6255 : NOR4_X1 port map( A1 => n4624, A2 => n4623, A3 => n4622, A4 => n4621
                           , ZN => n4626);
   U6256 : OAI22_X1 port map( A1 => n4627, A2 => n4652, B1 => n4626, B2 => 
                           n4625, ZN => IF_DecoderxN589);
   U6257 : AOI21_X1 port map( B1 => n4633, B2 => n6260, A => n4630, ZN => n4639
                           );
   U6258 : AND2_X1 port map( A1 => n6259, A2 => n4628, ZN => n4632);
   U6259 : INV_X1 port map( A => n4629, ZN => n4631);
   U6260 : AOI22_X1 port map( A1 => n4633, A2 => n4632, B1 => n4631, B2 => 
                           n4630, ZN => n4637);
   U6261 : NOR2_X1 port map( A1 => n4634, A2 => n4641, ZN => n4646);
   U6262 : NAND3_X1 port map( A1 => n4635, A2 => n4642, A3 => n4646, ZN => 
                           n4636);
   U6263 : OAI211_X1 port map( C1 => n4639, C2 => n4638, A => n4637, B => n4636
                           , ZN => IF_DecoderxN590);
   U6264 : NOR2_X1 port map( A1 => rst, A2 => n6319, ZN => IF_DecoderxN592);
   U6265 : NOR2_X1 port map( A1 => rst, A2 => n6320, ZN => IF_DecoderxN593);
   U6266 : NOR2_X1 port map( A1 => rst, A2 => n6321, ZN => IF_DecoderxN594);
   U6267 : NOR2_X1 port map( A1 => rst, A2 => n6322, ZN => IF_DecoderxN595);
   U6268 : INV_X1 port map( A => n4640, ZN => IF_DecoderxN591);
   U6269 : NOR2_X1 port map( A1 => rst, A2 => n6324, ZN => IF_DecoderxN597);
   U6270 : NOR2_X1 port map( A1 => rst, A2 => n6325, ZN => IF_DecoderxN598);
   U6271 : NOR2_X1 port map( A1 => rst, A2 => n6326, ZN => IF_DecoderxN599);
   U6272 : NOR2_X1 port map( A1 => rst, A2 => n6327, ZN => IF_DecoderxN600);
   U6273 : NOR2_X1 port map( A1 => rst, A2 => n6328, ZN => IF_DecoderxN601);
   U6274 : NOR2_X1 port map( A1 => rst, A2 => n6210, ZN => IF_DecoderxN603);
   U6275 : NOR2_X1 port map( A1 => rst, A2 => n6211, ZN => IF_DecoderxN604);
   U6276 : NOR2_X1 port map( A1 => rst, A2 => n6212, ZN => IF_DecoderxN605);
   U6277 : NOR2_X1 port map( A1 => rst, A2 => n6213, ZN => IF_DecoderxN606);
   U6278 : NOR2_X1 port map( A1 => n4642, A2 => n4641, ZN => n4644);
   U6279 : AOI21_X1 port map( B1 => n4651, B2 => n4644, A => n4643, ZN => 
                           IF_DecoderxN552);
   U6280 : AND2_X1 port map( A1 => n4646, A2 => n4645, ZN => IF_DecoderxN549);
   U6281 : INV_X1 port map( A => n4647, ZN => n4650);
   U6282 : OAI22_X1 port map( A1 => n4651, A2 => n4650, B1 => n4649, B2 => 
                           n4648, ZN => IF_DecoderxN550);
   U6283 : AOI21_X1 port map( B1 => n4654, B2 => n4653, A => n4652, ZN => 
                           IF_DecoderxN551);
   U6284 : NAND3_X1 port map( A1 => CtlToRegs_port_dst_1_port, A2 => 
                           CtlToRegs_port_dst_2_port, A3 => 
                           CtlToRegs_port_dst_0_port, ZN => n4664);
   U6285 : NAND4_X1 port map( A1 => CtlToRegs_port_notify, A2 => 
                           CtlToRegs_port_dst_4_port, A3 => 
                           CtlToRegs_port_dst_3_port, A4 => CtlToRegs_port_req,
                           ZN => n4657);
   U6286 : OAI21_X1 port map( B1 => n4664, B2 => n4657, A => n4667, ZN => 
                           IF_RegsxN659);
   U6287 : NAND3_X1 port map( A1 => CtlToRegs_port_dst_2_port, A2 => 
                           CtlToRegs_port_dst_1_port, A3 => n6233, ZN => n4665)
                           ;
   U6288 : OAI21_X1 port map( B1 => n4657, B2 => n4665, A => n4667, ZN => 
                           IF_RegsxN692);
   U6289 : NAND3_X1 port map( A1 => CtlToRegs_port_dst_2_port, A2 => 
                           CtlToRegs_port_dst_0_port, A3 => n6198, ZN => n4666)
                           ;
   U6290 : OAI21_X1 port map( B1 => n4657, B2 => n4666, A => n4667, ZN => 
                           IF_RegsxN693);
   U6291 : NAND3_X1 port map( A1 => CtlToRegs_port_dst_2_port, A2 => n6198, A3 
                           => n6233, ZN => n4668);
   U6292 : OAI21_X1 port map( B1 => n4657, B2 => n4668, A => n4671, ZN => 
                           IF_RegsxN694);
   U6293 : NOR2_X1 port map( A1 => CtlToRegs_port_dst_2_port, A2 => n6233, ZN 
                           => n4655);
   U6294 : NAND2_X1 port map( A1 => CtlToRegs_port_dst_1_port, A2 => n4655, ZN 
                           => n4669);
   U6295 : OAI21_X1 port map( B1 => n4657, B2 => n4669, A => n4667, ZN => 
                           IF_RegsxN695);
   U6296 : NOR2_X1 port map( A1 => CtlToRegs_port_dst_2_port, A2 => 
                           CtlToRegs_port_dst_0_port, ZN => n4656);
   U6297 : NAND2_X1 port map( A1 => CtlToRegs_port_dst_1_port, A2 => n4656, ZN 
                           => n4670);
   U6298 : OAI21_X1 port map( B1 => n4657, B2 => n4670, A => n6178, ZN => 
                           IF_RegsxN696);
   U6299 : NAND2_X1 port map( A1 => n4655, A2 => n6198, ZN => n4673);
   U6300 : OAI21_X1 port map( B1 => n4657, B2 => n4673, A => n4667, ZN => 
                           IF_RegsxN697);
   U6301 : NAND2_X1 port map( A1 => n4656, A2 => n6198, ZN => n4662);
   U6302 : OAI21_X1 port map( B1 => n4657, B2 => n4662, A => n4671, ZN => 
                           IF_RegsxN698);
   U6303 : NAND2_X1 port map( A1 => CtlToRegs_port_notify, A2 => 
                           CtlToRegs_port_req, ZN => n4659);
   U6304 : NOR2_X1 port map( A1 => CtlToRegs_port_dst_3_port, A2 => n4659, ZN 
                           => n4663);
   U6305 : NAND2_X1 port map( A1 => CtlToRegs_port_dst_4_port, A2 => n4663, ZN 
                           => n4658);
   U6306 : OAI21_X1 port map( B1 => n4664, B2 => n4658, A => n4667, ZN => 
                           IF_RegsxN699);
   U6307 : OAI21_X1 port map( B1 => n4665, B2 => n4658, A => n6178, ZN => 
                           IF_RegsxN700);
   U6308 : OAI21_X1 port map( B1 => n4666, B2 => n4658, A => n4667, ZN => 
                           IF_RegsxN701);
   U6309 : OAI21_X1 port map( B1 => n4668, B2 => n4658, A => n6178, ZN => 
                           IF_RegsxN702);
   U6310 : OAI21_X1 port map( B1 => n4669, B2 => n4658, A => n4667, ZN => 
                           IF_RegsxN703);
   U6311 : OAI21_X1 port map( B1 => n4670, B2 => n4658, A => n4671, ZN => 
                           IF_RegsxN704);
   U6312 : OAI21_X1 port map( B1 => n4673, B2 => n4658, A => n4667, ZN => 
                           IF_RegsxN705);
   U6313 : OAI21_X1 port map( B1 => n4662, B2 => n4658, A => n6178, ZN => 
                           IF_RegsxN706);
   U6314 : INV_X1 port map( A => n4659, ZN => n4660);
   U6315 : NAND3_X1 port map( A1 => CtlToRegs_port_dst_3_port, A2 => n4660, A3 
                           => n6235, ZN => n4661);
   U6316 : OAI21_X1 port map( B1 => n4664, B2 => n4661, A => n4667, ZN => 
                           IF_RegsxN707);
   U6317 : OAI21_X1 port map( B1 => n4665, B2 => n4661, A => n4671, ZN => 
                           IF_RegsxN708);
   U6318 : OAI21_X1 port map( B1 => n4666, B2 => n4661, A => n4667, ZN => 
                           IF_RegsxN709);
   U6319 : OAI21_X1 port map( B1 => n4668, B2 => n4661, A => n6178, ZN => 
                           IF_RegsxN710);
   U6320 : OAI21_X1 port map( B1 => n4669, B2 => n4661, A => n4667, ZN => 
                           IF_RegsxN711);
   U6321 : OAI21_X1 port map( B1 => n4670, B2 => n4661, A => n6178, ZN => 
                           IF_RegsxN712);
   U6322 : OAI21_X1 port map( B1 => n4673, B2 => n4661, A => n4667, ZN => 
                           IF_RegsxN713);
   U6323 : OAI21_X1 port map( B1 => n4662, B2 => n4661, A => n6178, ZN => 
                           IF_RegsxN714);
   U6324 : NAND2_X1 port map( A1 => n4663, A2 => n6235, ZN => n4672);
   U6325 : OAI21_X1 port map( B1 => n4664, B2 => n4672, A => n4667, ZN => 
                           IF_RegsxN715);
   U6326 : OAI21_X1 port map( B1 => n4665, B2 => n4672, A => n6178, ZN => 
                           IF_RegsxN716);
   U6327 : OAI21_X1 port map( B1 => n4666, B2 => n4672, A => n4667, ZN => 
                           IF_RegsxN717);
   U6328 : OAI21_X1 port map( B1 => n4668, B2 => n4672, A => n4667, ZN => 
                           IF_RegsxN718);
   U6329 : OAI21_X1 port map( B1 => n4669, B2 => n4672, A => n6178, ZN => 
                           IF_RegsxN719);
   U6330 : OAI21_X1 port map( B1 => n4670, B2 => n4672, A => n6178, ZN => 
                           IF_RegsxN720);
   U6331 : OAI21_X1 port map( B1 => n4673, B2 => n4672, A => n4671, ZN => 
                           IF_RegsxN721);
   U6332 : NAND2_X1 port map( A1 => CtlToRegs_port_src2_3_port, A2 => 
                           CtlToRegs_port_src2_2_port, ZN => n4674);
   U6333 : OR2_X1 port map( A1 => CtlToRegs_port_src2_4_port, A2 => n4674, ZN 
                           => n4690);
   U6334 : NOR2_X1 port map( A1 => n2952, A2 => n4690, ZN => n5345);
   U6335 : CLKBUF_X1 port map( A => n5345, Z => n5385);
   U6336 : AND2_X1 port map( A1 => CtlToRegs_port_src2_0_port, A2 => n5385, ZN 
                           => n5415);
   U6337 : CLKBUF_X1 port map( A => n6266, Z => n4917);
   U6338 : NAND2_X1 port map( A1 => n2952, A2 => n4917, ZN => n4696);
   U6339 : NOR3_X1 port map( A1 => CtlToRegs_port_src2_3_port, A2 => 
                           CtlToRegs_port_src2_2_port, A3 => n4696, ZN => n4813
                           );
   U6340 : CLKBUF_X1 port map( A => n4813, Z => n5340);
   U6341 : NAND3_X1 port map( A1 => CtlToRegs_port_src2_3_port, A2 => n6206, A3
                           => n6257, ZN => n4687);
   U6342 : NAND2_X1 port map( A1 => CtlToRegs_port_src2_0_port, A2 => n2952, ZN
                           => n4688);
   U6343 : NOR2_X1 port map( A1 => n4687, A2 => n4688, ZN => n5401);
   U6344 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_480_port, B1 
                           => IF_Regsxreg_file_704_port, B2 => n5401, ZN => 
                           n4677);
   U6345 : NAND3_X1 port map( A1 => CtlToRegs_port_src2_2_port, A2 => n6206, A3
                           => n6265, ZN => n4685);
   U6346 : NOR2_X1 port map( A1 => n4685, A2 => n4688, ZN => n5314);
   U6347 : CLKBUF_X1 port map( A => n5314, Z => n5409);
   U6348 : NAND3_X1 port map( A1 => CtlToRegs_port_src2_4_port, A2 => 
                           CtlToRegs_port_src2_3_port, A3 => 
                           CtlToRegs_port_src2_2_port, ZN => n4680);
   U6349 : NOR2_X1 port map( A1 => n4696, A2 => n4680, ZN => n5075);
   U6350 : AOI22_X1 port map( A1 => IF_Regsxreg_file_832_port, A2 => n5409, B1 
                           => IF_Regsxreg_file_96_port, B2 => n5075, ZN => 
                           n4676);
   U6351 : NOR2_X1 port map( A1 => n4680, A2 => n4688, ZN => n5240);
   U6352 : CLKBUF_X1 port map( A => n5240, Z => n5378);
   U6353 : NOR2_X1 port map( A1 => n4690, A2 => n4688, ZN => n5250);
   U6354 : AOI22_X1 port map( A1 => IF_Regsxreg_file_64_port, A2 => n5378, B1 
                           => IF_Regsxreg_file_576_port, B2 => n5250, ZN => 
                           n4675);
   U6355 : NAND3_X1 port map( A1 => n4677, A2 => n4676, A3 => n4675, ZN => 
                           n4678);
   U6356 : AOI21_X1 port map( B1 => IF_Regsxreg_file_512_port, B2 => n5415, A 
                           => n4678, ZN => n4707);
   U6357 : NAND3_X1 port map( A1 => CtlToRegs_port_src2_3_port, A2 => 
                           CtlToRegs_port_src2_4_port, A3 => n6257, ZN => n4689
                           );
   U6358 : NOR2_X1 port map( A1 => n2952, A2 => n4689, ZN => n5294);
   U6359 : CLKBUF_X1 port map( A => n5294, Z => n5387);
   U6360 : NOR2_X1 port map( A1 => n2952, A2 => n4687, ZN => n5391);
   U6361 : CLKBUF_X1 port map( A => n5391, Z => n5320);
   U6362 : AOI22_X1 port map( A1 => IF_Regsxreg_file_160_port, A2 => n5387, B1 
                           => IF_Regsxreg_file_672_port, B2 => n5320, ZN => 
                           n4684);
   U6363 : NOR4_X1 port map( A1 => CtlToRegs_port_src2_4_port, A2 => 
                           CtlToRegs_port_src2_3_port, A3 => 
                           CtlToRegs_port_src2_2_port, A4 => n2952, ZN => n4697
                           );
   U6364 : CLKBUF_X1 port map( A => n4697, Z => n5389);
   U6365 : AOI22_X1 port map( A1 => IF_Regsxreg_file_544_port, A2 => n5385, B1 
                           => IF_Regsxreg_file_928_port, B2 => n5389, ZN => 
                           n4683);
   U6366 : NOR2_X1 port map( A1 => n2952, A2 => n4685, ZN => n5157);
   U6367 : CLKBUF_X1 port map( A => n5157, Z => n5384);
   U6368 : NOR2_X1 port map( A1 => CtlToRegs_port_src2_3_port, A2 => 
                           CtlToRegs_port_src2_2_port, ZN => n4679);
   U6369 : NAND2_X1 port map( A1 => CtlToRegs_port_src2_4_port, A2 => n4679, ZN
                           => n4686);
   U6370 : NOR2_X1 port map( A1 => n2952, A2 => n4686, ZN => n5386);
   U6371 : AOI22_X1 port map( A1 => IF_Regsxreg_file_800_port, A2 => n5384, B1 
                           => IF_Regsxreg_file_416_port, B2 => n5386, ZN => 
                           n4682);
   U6372 : NAND3_X1 port map( A1 => CtlToRegs_port_src2_4_port, A2 => 
                           CtlToRegs_port_src2_2_port, A3 => n6265, ZN => n4695
                           );
   U6373 : NOR2_X1 port map( A1 => n2952, A2 => n4695, ZN => n5390);
   U6374 : CLKBUF_X1 port map( A => n5390, Z => n5346);
   U6375 : NOR2_X1 port map( A1 => n2952, A2 => n4680, ZN => n5388);
   U6376 : CLKBUF_X1 port map( A => n5388, Z => n5319);
   U6377 : AOI22_X1 port map( A1 => IF_Regsxreg_file_288_port, A2 => n5346, B1 
                           => IF_Regsxreg_file_32_port, B2 => n5319, ZN => 
                           n4681);
   U6378 : NAND4_X1 port map( A1 => n4684, A2 => n4683, A3 => n4682, A4 => 
                           n4681, ZN => n4704);
   U6379 : NOR4_X1 port map( A1 => CtlToRegs_port_src2_4_port, A2 => 
                           CtlToRegs_port_src2_3_port, A3 => 
                           CtlToRegs_port_src2_2_port, A4 => n4688, ZN => n5264
                           );
   U6380 : CLKBUF_X1 port map( A => n5264, Z => n5352);
   U6381 : NOR2_X1 port map( A1 => n4695, A2 => n4688, ZN => n5354);
   U6382 : CLKBUF_X1 port map( A => n5354, Z => n5399);
   U6383 : AOI22_X1 port map( A1 => IF_Regsxreg_file_960_port, A2 => n5352, B1 
                           => IF_Regsxreg_file_320_port, B2 => n5399, ZN => 
                           n4694);
   U6384 : NOR2_X1 port map( A1 => n4696, A2 => n4685, ZN => n5396);
   U6385 : CLKBUF_X1 port map( A => n5396, Z => n5300);
   U6386 : NOR2_X1 port map( A1 => n4686, A2 => n4688, ZN => n5373);
   U6387 : CLKBUF_X1 port map( A => n5373, Z => n5325);
   U6388 : AOI22_X1 port map( A1 => IF_Regsxreg_file_864_port, A2 => n5300, B1 
                           => IF_Regsxreg_file_448_port, B2 => n5325, ZN => 
                           n4693);
   U6389 : NOR2_X1 port map( A1 => n4696, A2 => n4689, ZN => n5299);
   U6390 : NOR2_X1 port map( A1 => n4696, A2 => n4687, ZN => n5273);
   U6391 : AOI22_X1 port map( A1 => IF_Regsxreg_file_224_port, A2 => n5299, B1 
                           => IF_Regsxreg_file_736_port, B2 => n5273, ZN => 
                           n4692);
   U6392 : NOR2_X1 port map( A1 => n4689, A2 => n4688, ZN => n5398);
   U6393 : CLKBUF_X1 port map( A => n5398, Z => n5353);
   U6394 : NOR2_X1 port map( A1 => n4696, A2 => n4690, ZN => n5162);
   U6395 : CLKBUF_X1 port map( A => n5162, Z => n5375);
   U6396 : AOI22_X1 port map( A1 => IF_Regsxreg_file_192_port, A2 => n5353, B1 
                           => IF_Regsxreg_file_608_port, B2 => n5375, ZN => 
                           n4691);
   U6397 : NAND4_X1 port map( A1 => n4694, A2 => n4693, A3 => n4692, A4 => 
                           n4691, ZN => n4703);
   U6398 : AND2_X1 port map( A1 => CtlToRegs_port_src2_0_port, A2 => n5384, ZN 
                           => n5411);
   U6399 : CLKBUF_X1 port map( A => n5411, Z => n5279);
   U6400 : NOR2_X1 port map( A1 => n4696, A2 => n4695, ZN => n5400);
   U6401 : CLKBUF_X1 port map( A => n5400, Z => n5351);
   U6402 : AOI22_X1 port map( A1 => IF_Regsxreg_file_768_port, A2 => n5279, B1 
                           => IF_Regsxreg_file_352_port, B2 => n5351, ZN => 
                           n4701);
   U6403 : AND2_X1 port map( A1 => CtlToRegs_port_src2_0_port, A2 => n5346, ZN 
                           => n5363);
   U6404 : AND2_X1 port map( A1 => CtlToRegs_port_src2_0_port, A2 => n5387, ZN 
                           => n5361);
   U6405 : CLKBUF_X1 port map( A => n5361, Z => n5412);
   U6406 : AOI22_X1 port map( A1 => IF_Regsxreg_file_256_port, A2 => n5363, B1 
                           => IF_Regsxreg_file_128_port, B2 => n5412, ZN => 
                           n4700);
   U6407 : CLKBUF_X1 port map( A => n5386, Z => n5293);
   U6408 : AND2_X1 port map( A1 => CtlToRegs_port_src2_0_port, A2 => n5293, ZN 
                           => n5278);
   U6409 : AND2_X1 port map( A1 => CtlToRegs_port_src2_0_port, A2 => n5319, ZN 
                           => n5408);
   U6410 : CLKBUF_X1 port map( A => n5408, Z => n5362);
   U6411 : AOI22_X1 port map( A1 => IF_Regsxreg_file_384_port, A2 => n5278, B1 
                           => IF_Regsxreg_file_0_port, B2 => n5362, ZN => n4699
                           );
   U6412 : CLKBUF_X1 port map( A => n4697, Z => n5245);
   U6413 : AND2_X1 port map( A1 => CtlToRegs_port_src2_0_port, A2 => n5245, ZN 
                           => n5383);
   U6414 : AND2_X1 port map( A1 => CtlToRegs_port_src2_0_port, A2 => n5320, ZN 
                           => n5410);
   U6415 : CLKBUF_X1 port map( A => n5410, Z => n5360);
   U6416 : AOI22_X1 port map( A1 => IF_Regsxreg_file_896_port, A2 => n5383, B1 
                           => IF_Regsxreg_file_640_port, B2 => n5360, ZN => 
                           n4698);
   U6417 : NAND4_X1 port map( A1 => n4701, A2 => n4700, A3 => n4699, A4 => 
                           n4698, ZN => n4702);
   U6418 : AOI211_X1 port map( C1 => n4917, C2 => n4704, A => n4703, B => n4702
                           , ZN => n4706);
   U6419 : AOI21_X1 port map( B1 => n6206, B2 => n5340, A => rst, ZN => n4705);
   U6420 : INV_X1 port map( A => n4705, ZN => n5216);
   U6421 : AOI21_X1 port map( B1 => n4707, B2 => n4706, A => n5216, ZN => 
                           IF_RegsxN627);
   U6422 : AOI22_X1 port map( A1 => n4813, A2 => IF_Regsxreg_file_481_port, B1 
                           => n5373, B2 => IF_Regsxreg_file_449_port, ZN => 
                           n4710);
   U6423 : AOI22_X1 port map( A1 => n5399, A2 => IF_Regsxreg_file_321_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_353_port, ZN => 
                           n4709);
   U6424 : CLKBUF_X1 port map( A => n5299, Z => n5377);
   U6425 : AOI22_X1 port map( A1 => n5075, A2 => IF_Regsxreg_file_97_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_225_port, ZN => 
                           n4708);
   U6426 : NAND3_X1 port map( A1 => n4710, A2 => n4709, A3 => n4708, ZN => 
                           n4711);
   U6427 : AOI21_X1 port map( B1 => n5383, B2 => IF_Regsxreg_file_897_port, A 
                           => n4711, ZN => n4728);
   U6428 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_673_port, B1 
                           => n5385, B2 => IF_Regsxreg_file_545_port, ZN => 
                           n4715);
   U6429 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_161_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_289_port, ZN => 
                           n4714);
   U6430 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_929_port, B1 
                           => n5384, B2 => IF_Regsxreg_file_801_port, ZN => 
                           n4713);
   U6431 : AOI22_X1 port map( A1 => n5293, A2 => IF_Regsxreg_file_417_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_33_port, ZN => 
                           n4712);
   U6432 : NAND4_X1 port map( A1 => n4715, A2 => n4714, A3 => n4713, A4 => 
                           n4712, ZN => n4726);
   U6433 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_833_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_609_port, ZN => 
                           n4719);
   U6434 : CLKBUF_X1 port map( A => n5273, Z => n5402);
   U6435 : AOI22_X1 port map( A1 => n5352, A2 => IF_Regsxreg_file_961_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_737_port, ZN => 
                           n4718);
   U6436 : AOI22_X1 port map( A1 => n5250, A2 => IF_Regsxreg_file_577_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_193_port, ZN => 
                           n4717);
   U6437 : AOI22_X1 port map( A1 => n5401, A2 => IF_Regsxreg_file_705_port, B1 
                           => n5300, B2 => IF_Regsxreg_file_865_port, ZN => 
                           n4716);
   U6438 : NAND4_X1 port map( A1 => n4719, A2 => n4718, A3 => n4717, A4 => 
                           n4716, ZN => n4725);
   U6439 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_65_port, B1 
                           => n5360, B2 => IF_Regsxreg_file_641_port, ZN => 
                           n4723);
   U6440 : AOI22_X1 port map( A1 => n5279, A2 => IF_Regsxreg_file_769_port, B1 
                           => n5412, B2 => IF_Regsxreg_file_129_port, ZN => 
                           n4722);
   U6441 : CLKBUF_X1 port map( A => n5278, Z => n5414);
   U6442 : AOI22_X1 port map( A1 => n5363, A2 => IF_Regsxreg_file_257_port, B1 
                           => n5414, B2 => IF_Regsxreg_file_385_port, ZN => 
                           n4721);
   U6443 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_513_port, B1 
                           => n5362, B2 => IF_Regsxreg_file_1_port, ZN => n4720
                           );
   U6444 : NAND4_X1 port map( A1 => n4723, A2 => n4722, A3 => n4721, A4 => 
                           n4720, ZN => n4724);
   U6445 : AOI211_X1 port map( C1 => n4917, C2 => n4726, A => n4725, B => n4724
                           , ZN => n4727);
   U6446 : AOI21_X1 port map( B1 => n4728, B2 => n4727, A => n5216, ZN => 
                           IF_RegsxN628);
   U6447 : CLKBUF_X1 port map( A => n4813, Z => n5374);
   U6448 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_482_port, B1 
                           => n5314, B2 => IF_Regsxreg_file_834_port, ZN => 
                           n4731);
   U6449 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_66_port, B1 
                           => n5400, B2 => IF_Regsxreg_file_354_port, ZN => 
                           n4730);
   U6450 : CLKBUF_X1 port map( A => n5264, Z => n5376);
   U6451 : AOI22_X1 port map( A1 => n5376, A2 => IF_Regsxreg_file_962_port, B1 
                           => n5399, B2 => IF_Regsxreg_file_322_port, ZN => 
                           n4729);
   U6452 : NAND3_X1 port map( A1 => n4731, A2 => n4730, A3 => n4729, ZN => 
                           n4732);
   U6453 : AOI21_X1 port map( B1 => n5383, B2 => IF_Regsxreg_file_898_port, A 
                           => n4732, ZN => n4749);
   U6454 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_930_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_34_port, ZN => 
                           n4736);
   U6455 : AOI22_X1 port map( A1 => n5385, A2 => IF_Regsxreg_file_546_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_290_port, ZN => 
                           n4735);
   U6456 : AOI22_X1 port map( A1 => n5391, A2 => IF_Regsxreg_file_674_port, B1 
                           => n5384, B2 => IF_Regsxreg_file_802_port, ZN => 
                           n4734);
   U6457 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_162_port, B1 
                           => n5293, B2 => IF_Regsxreg_file_418_port, ZN => 
                           n4733);
   U6458 : NAND4_X1 port map( A1 => n4736, A2 => n4735, A3 => n4734, A4 => 
                           n4733, ZN => n4747);
   U6459 : AOI22_X1 port map( A1 => n5325, A2 => IF_Regsxreg_file_450_port, B1 
                           => n5273, B2 => IF_Regsxreg_file_738_port, ZN => 
                           n4740);
   U6460 : AOI22_X1 port map( A1 => n5300, A2 => IF_Regsxreg_file_866_port, B1 
                           => n5398, B2 => IF_Regsxreg_file_194_port, ZN => 
                           n4739);
   U6461 : CLKBUF_X1 port map( A => n5401, Z => n5330);
   U6462 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_706_port, B1 
                           => n5075, B2 => IF_Regsxreg_file_98_port, ZN => 
                           n4738);
   U6463 : AOI22_X1 port map( A1 => n5250, A2 => IF_Regsxreg_file_578_port, B1 
                           => n5162, B2 => IF_Regsxreg_file_610_port, ZN => 
                           n4737);
   U6464 : NAND4_X1 port map( A1 => n4740, A2 => n4739, A3 => n4738, A4 => 
                           n4737, ZN => n4746);
   U6465 : AOI22_X1 port map( A1 => n5377, A2 => IF_Regsxreg_file_226_port, B1 
                           => n5278, B2 => IF_Regsxreg_file_386_port, ZN => 
                           n4744);
   U6466 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_514_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_2_port, ZN => n4743
                           );
   U6467 : AOI22_X1 port map( A1 => n5411, A2 => IF_Regsxreg_file_770_port, B1 
                           => n5363, B2 => IF_Regsxreg_file_258_port, ZN => 
                           n4742);
   U6468 : AOI22_X1 port map( A1 => n5361, A2 => IF_Regsxreg_file_130_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_642_port, ZN => 
                           n4741);
   U6469 : NAND4_X1 port map( A1 => n4744, A2 => n4743, A3 => n4742, A4 => 
                           n4741, ZN => n4745);
   U6470 : AOI211_X1 port map( C1 => n4917, C2 => n4747, A => n4746, B => n4745
                           , ZN => n4748);
   U6471 : AOI21_X1 port map( B1 => n4749, B2 => n4748, A => n5216, ZN => 
                           IF_RegsxN629);
   U6472 : AOI22_X1 port map( A1 => n4813, A2 => IF_Regsxreg_file_483_port, B1 
                           => n5162, B2 => IF_Regsxreg_file_611_port, ZN => 
                           n4752);
   U6473 : AOI22_X1 port map( A1 => n5314, A2 => IF_Regsxreg_file_835_port, B1 
                           => n5273, B2 => IF_Regsxreg_file_739_port, ZN => 
                           n4751);
   U6474 : CLKBUF_X1 port map( A => n5250, Z => n5397);
   U6475 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_579_port, B1 
                           => n5400, B2 => IF_Regsxreg_file_355_port, ZN => 
                           n4750);
   U6476 : NAND3_X1 port map( A1 => n4752, A2 => n4751, A3 => n4750, ZN => 
                           n4753);
   U6477 : AOI21_X1 port map( B1 => n5383, B2 => IF_Regsxreg_file_899_port, A 
                           => n4753, ZN => n4770);
   U6478 : AOI22_X1 port map( A1 => n5384, A2 => IF_Regsxreg_file_803_port, B1 
                           => n5293, B2 => IF_Regsxreg_file_419_port, ZN => 
                           n4757);
   U6479 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_675_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_291_port, ZN => 
                           n4756);
   U6480 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_931_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_35_port, ZN => 
                           n4755);
   U6481 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_163_port, B1 
                           => n5385, B2 => IF_Regsxreg_file_547_port, ZN => 
                           n4754);
   U6482 : NAND4_X1 port map( A1 => n4757, A2 => n4756, A3 => n4755, A4 => 
                           n4754, ZN => n4768);
   U6483 : AOI22_X1 port map( A1 => n5300, A2 => IF_Regsxreg_file_867_port, B1 
                           => n5373, B2 => IF_Regsxreg_file_451_port, ZN => 
                           n4761);
   U6484 : AOI22_X1 port map( A1 => n5401, A2 => IF_Regsxreg_file_707_port, B1 
                           => n5299, B2 => IF_Regsxreg_file_227_port, ZN => 
                           n4760);
   U6485 : AOI22_X1 port map( A1 => n5376, A2 => IF_Regsxreg_file_963_port, B1 
                           => n5398, B2 => IF_Regsxreg_file_195_port, ZN => 
                           n4759);
   U6486 : AOI22_X1 port map( A1 => n5240, A2 => IF_Regsxreg_file_67_port, B1 
                           => n5354, B2 => IF_Regsxreg_file_323_port, ZN => 
                           n4758);
   U6487 : NAND4_X1 port map( A1 => n4761, A2 => n4760, A3 => n4759, A4 => 
                           n4758, ZN => n4767);
   U6488 : CLKBUF_X1 port map( A => n5075, Z => n5403);
   U6489 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_99_port, B1 
                           => n5363, B2 => IF_Regsxreg_file_259_port, ZN => 
                           n4765);
   U6490 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_515_port, B1 
                           => n5361, B2 => IF_Regsxreg_file_131_port, ZN => 
                           n4764);
   U6491 : AOI22_X1 port map( A1 => n5362, A2 => IF_Regsxreg_file_3_port, B1 =>
                           n5410, B2 => IF_Regsxreg_file_643_port, ZN => n4763)
                           ;
   U6492 : AOI22_X1 port map( A1 => n5411, A2 => IF_Regsxreg_file_771_port, B1 
                           => n5278, B2 => IF_Regsxreg_file_387_port, ZN => 
                           n4762);
   U6493 : NAND4_X1 port map( A1 => n4765, A2 => n4764, A3 => n4763, A4 => 
                           n4762, ZN => n4766);
   U6494 : AOI211_X1 port map( C1 => n4917, C2 => n4768, A => n4767, B => n4766
                           , ZN => n4769);
   U6495 : AOI21_X1 port map( B1 => n4770, B2 => n4769, A => n5216, ZN => 
                           IF_RegsxN630);
   U6496 : AOI22_X1 port map( A1 => n4813, A2 => IF_Regsxreg_file_484_port, B1 
                           => n5400, B2 => IF_Regsxreg_file_356_port, ZN => 
                           n4773);
   U6497 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_580_port, B1 
                           => n5273, B2 => IF_Regsxreg_file_740_port, ZN => 
                           n4772);
   U6498 : AOI22_X1 port map( A1 => n5399, A2 => IF_Regsxreg_file_324_port, B1 
                           => n5299, B2 => IF_Regsxreg_file_228_port, ZN => 
                           n4771);
   U6499 : NAND3_X1 port map( A1 => n4773, A2 => n4772, A3 => n4771, ZN => 
                           n4774);
   U6500 : AOI21_X1 port map( B1 => n5383, B2 => IF_Regsxreg_file_900_port, A 
                           => n4774, ZN => n4791);
   U6501 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_164_port, B1 
                           => n5157, B2 => IF_Regsxreg_file_804_port, ZN => 
                           n4778);
   U6502 : AOI22_X1 port map( A1 => n5293, A2 => IF_Regsxreg_file_420_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_36_port, ZN => 
                           n4777);
   U6503 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_676_port, B1 
                           => n5245, B2 => IF_Regsxreg_file_932_port, ZN => 
                           n4776);
   U6504 : AOI22_X1 port map( A1 => n5345, A2 => IF_Regsxreg_file_548_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_292_port, ZN => 
                           n4775);
   U6505 : NAND4_X1 port map( A1 => n4778, A2 => n4777, A3 => n4776, A4 => 
                           n4775, ZN => n4789);
   U6506 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_836_port, B1 
                           => n5376, B2 => IF_Regsxreg_file_964_port, ZN => 
                           n4782);
   U6507 : AOI22_X1 port map( A1 => n5373, A2 => IF_Regsxreg_file_452_port, B1 
                           => n5162, B2 => IF_Regsxreg_file_612_port, ZN => 
                           n4781);
   U6508 : AOI22_X1 port map( A1 => n5075, A2 => IF_Regsxreg_file_100_port, B1 
                           => n5240, B2 => IF_Regsxreg_file_68_port, ZN => 
                           n4780);
   U6509 : AOI22_X1 port map( A1 => n5396, A2 => IF_Regsxreg_file_868_port, B1 
                           => n5398, B2 => IF_Regsxreg_file_196_port, ZN => 
                           n4779);
   U6510 : NAND4_X1 port map( A1 => n4782, A2 => n4781, A3 => n4780, A4 => 
                           n4779, ZN => n4788);
   U6511 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_708_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_644_port, ZN => 
                           n4786);
   U6512 : CLKBUF_X1 port map( A => n5363, Z => n5413);
   U6513 : AOI22_X1 port map( A1 => n5413, A2 => IF_Regsxreg_file_260_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_4_port, ZN => n4785
                           );
   U6514 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_516_port, B1 
                           => n5278, B2 => IF_Regsxreg_file_388_port, ZN => 
                           n4784);
   U6515 : AOI22_X1 port map( A1 => n5411, A2 => IF_Regsxreg_file_772_port, B1 
                           => n5361, B2 => IF_Regsxreg_file_132_port, ZN => 
                           n4783);
   U6516 : NAND4_X1 port map( A1 => n4786, A2 => n4785, A3 => n4784, A4 => 
                           n4783, ZN => n4787);
   U6517 : AOI211_X1 port map( C1 => n4917, C2 => n4789, A => n4788, B => n4787
                           , ZN => n4790);
   U6518 : AOI21_X1 port map( B1 => n4791, B2 => n4790, A => n5216, ZN => 
                           IF_RegsxN631);
   U6519 : AOI22_X1 port map( A1 => n4813, A2 => IF_Regsxreg_file_485_port, B1 
                           => n5396, B2 => IF_Regsxreg_file_869_port, ZN => 
                           n4794);
   U6520 : AOI22_X1 port map( A1 => n5075, A2 => IF_Regsxreg_file_101_port, B1 
                           => n5273, B2 => IF_Regsxreg_file_741_port, ZN => 
                           n4793);
   U6521 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_709_port, B1 
                           => n5250, B2 => IF_Regsxreg_file_581_port, ZN => 
                           n4792);
   U6522 : NAND3_X1 port map( A1 => n4794, A2 => n4793, A3 => n4792, ZN => 
                           n4795);
   U6523 : AOI21_X1 port map( B1 => n5362, B2 => IF_Regsxreg_file_5_port, A => 
                           n4795, ZN => n4812);
   U6524 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_677_port, B1 
                           => n5157, B2 => IF_Regsxreg_file_805_port, ZN => 
                           n4799);
   U6525 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_933_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_293_port, ZN => 
                           n4798);
   U6526 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_165_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_37_port, ZN => 
                           n4797);
   U6527 : AOI22_X1 port map( A1 => n5345, A2 => IF_Regsxreg_file_549_port, B1 
                           => n5293, B2 => IF_Regsxreg_file_421_port, ZN => 
                           n4796);
   U6528 : NAND4_X1 port map( A1 => n4799, A2 => n4798, A3 => n4797, A4 => 
                           n4796, ZN => n4810);
   U6529 : AOI22_X1 port map( A1 => n5376, A2 => IF_Regsxreg_file_965_port, B1 
                           => n5354, B2 => IF_Regsxreg_file_325_port, ZN => 
                           n4803);
   U6530 : AOI22_X1 port map( A1 => n5325, A2 => IF_Regsxreg_file_453_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_229_port, ZN => 
                           n4802);
   U6531 : AOI22_X1 port map( A1 => n5314, A2 => IF_Regsxreg_file_837_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_613_port, ZN => 
                           n4801);
   U6532 : AOI22_X1 port map( A1 => n5240, A2 => IF_Regsxreg_file_69_port, B1 
                           => n5400, B2 => IF_Regsxreg_file_357_port, ZN => 
                           n4800);
   U6533 : NAND4_X1 port map( A1 => n4803, A2 => n4802, A3 => n4801, A4 => 
                           n4800, ZN => n4809);
   U6534 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_517_port, B1 
                           => n5398, B2 => IF_Regsxreg_file_197_port, ZN => 
                           n4807);
   U6535 : AOI22_X1 port map( A1 => n5411, A2 => IF_Regsxreg_file_773_port, B1 
                           => n5361, B2 => IF_Regsxreg_file_133_port, ZN => 
                           n4806);
   U6536 : AOI22_X1 port map( A1 => n5383, A2 => IF_Regsxreg_file_901_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_645_port, ZN => 
                           n4805);
   U6537 : AOI22_X1 port map( A1 => n5413, A2 => IF_Regsxreg_file_261_port, B1 
                           => n5278, B2 => IF_Regsxreg_file_389_port, ZN => 
                           n4804);
   U6538 : NAND4_X1 port map( A1 => n4807, A2 => n4806, A3 => n4805, A4 => 
                           n4804, ZN => n4808);
   U6539 : AOI211_X1 port map( C1 => n4917, C2 => n4810, A => n4809, B => n4808
                           , ZN => n4811);
   U6540 : AOI21_X1 port map( B1 => n4812, B2 => n4811, A => n5216, ZN => 
                           IF_RegsxN632);
   U6541 : AOI22_X1 port map( A1 => n4813, A2 => IF_Regsxreg_file_486_port, B1 
                           => n5401, B2 => IF_Regsxreg_file_710_port, ZN => 
                           n4816);
   U6542 : AOI22_X1 port map( A1 => n5376, A2 => IF_Regsxreg_file_966_port, B1 
                           => n5273, B2 => IF_Regsxreg_file_742_port, ZN => 
                           n4815);
   U6543 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_102_port, B1 
                           => n5240, B2 => IF_Regsxreg_file_70_port, ZN => 
                           n4814);
   U6544 : NAND3_X1 port map( A1 => n4816, A2 => n4815, A3 => n4814, ZN => 
                           n4817);
   U6545 : AOI21_X1 port map( B1 => n5362, B2 => IF_Regsxreg_file_6_port, A => 
                           n4817, ZN => n4834);
   U6546 : AOI22_X1 port map( A1 => n5384, A2 => IF_Regsxreg_file_806_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_294_port, ZN => 
                           n4821);
   U6547 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_166_port, B1 
                           => n5320, B2 => IF_Regsxreg_file_678_port, ZN => 
                           n4820);
   U6548 : AOI22_X1 port map( A1 => n5293, A2 => IF_Regsxreg_file_422_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_38_port, ZN => 
                           n4819);
   U6549 : AOI22_X1 port map( A1 => n5345, A2 => IF_Regsxreg_file_550_port, B1 
                           => n5245, B2 => IF_Regsxreg_file_934_port, ZN => 
                           n4818);
   U6550 : NAND4_X1 port map( A1 => n4821, A2 => n4820, A3 => n4819, A4 => 
                           n4818, ZN => n4832);
   U6551 : AOI22_X1 port map( A1 => n5325, A2 => IF_Regsxreg_file_454_port, B1 
                           => n5299, B2 => IF_Regsxreg_file_230_port, ZN => 
                           n4825);
   U6552 : AOI22_X1 port map( A1 => n5250, A2 => IF_Regsxreg_file_582_port, B1 
                           => n5300, B2 => IF_Regsxreg_file_870_port, ZN => 
                           n4824);
   U6553 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_838_port, B1 
                           => n5398, B2 => IF_Regsxreg_file_198_port, ZN => 
                           n4823);
   U6554 : AOI22_X1 port map( A1 => n5375, A2 => IF_Regsxreg_file_614_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_358_port, ZN => 
                           n4822);
   U6555 : NAND4_X1 port map( A1 => n4825, A2 => n4824, A3 => n4823, A4 => 
                           n4822, ZN => n4831);
   U6556 : AOI22_X1 port map( A1 => n5399, A2 => IF_Regsxreg_file_326_port, B1 
                           => n5363, B2 => IF_Regsxreg_file_262_port, ZN => 
                           n4829);
   U6557 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_518_port, B1 
                           => n5383, B2 => IF_Regsxreg_file_902_port, ZN => 
                           n4828);
   U6558 : AOI22_X1 port map( A1 => n5411, A2 => IF_Regsxreg_file_774_port, B1 
                           => n5278, B2 => IF_Regsxreg_file_390_port, ZN => 
                           n4827);
   U6559 : AOI22_X1 port map( A1 => n5361, A2 => IF_Regsxreg_file_134_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_646_port, ZN => 
                           n4826);
   U6560 : NAND4_X1 port map( A1 => n4829, A2 => n4828, A3 => n4827, A4 => 
                           n4826, ZN => n4830);
   U6561 : AOI211_X1 port map( C1 => n4917, C2 => n4832, A => n4831, B => n4830
                           , ZN => n4833);
   U6562 : AOI21_X1 port map( B1 => n4834, B2 => n4833, A => n5216, ZN => 
                           IF_RegsxN633);
   U6563 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_487_port, B1 
                           => n5314, B2 => IF_Regsxreg_file_839_port, ZN => 
                           n4837);
   U6564 : AOI22_X1 port map( A1 => n5399, A2 => IF_Regsxreg_file_327_port, B1 
                           => n5398, B2 => IF_Regsxreg_file_199_port, ZN => 
                           n4836);
   U6565 : AOI22_X1 port map( A1 => n5325, A2 => IF_Regsxreg_file_455_port, B1 
                           => n5299, B2 => IF_Regsxreg_file_231_port, ZN => 
                           n4835);
   U6566 : NAND3_X1 port map( A1 => n4837, A2 => n4836, A3 => n4835, ZN => 
                           n4838);
   U6567 : AOI21_X1 port map( B1 => n5411, B2 => IF_Regsxreg_file_775_port, A 
                           => n4838, ZN => n4855);
   U6568 : AOI22_X1 port map( A1 => n5293, A2 => IF_Regsxreg_file_423_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_295_port, ZN => 
                           n4842);
   U6569 : AOI22_X1 port map( A1 => n5385, A2 => IF_Regsxreg_file_551_port, B1 
                           => n5157, B2 => IF_Regsxreg_file_807_port, ZN => 
                           n4841);
   U6570 : AOI22_X1 port map( A1 => n5391, A2 => IF_Regsxreg_file_679_port, B1 
                           => n5245, B2 => IF_Regsxreg_file_935_port, ZN => 
                           n4840);
   U6571 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_167_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_39_port, ZN => 
                           n4839);
   U6572 : NAND4_X1 port map( A1 => n4842, A2 => n4841, A3 => n4840, A4 => 
                           n4839, ZN => n4853);
   U6573 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_583_port, B1 
                           => n5162, B2 => IF_Regsxreg_file_615_port, ZN => 
                           n4846);
   U6574 : AOI22_X1 port map( A1 => n5300, A2 => IF_Regsxreg_file_871_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_743_port, ZN => 
                           n4845);
   U6575 : AOI22_X1 port map( A1 => n5401, A2 => IF_Regsxreg_file_711_port, B1 
                           => n5075, B2 => IF_Regsxreg_file_103_port, ZN => 
                           n4844);
   U6576 : AOI22_X1 port map( A1 => n5376, A2 => IF_Regsxreg_file_967_port, B1 
                           => n5400, B2 => IF_Regsxreg_file_359_port, ZN => 
                           n4843);
   U6577 : NAND4_X1 port map( A1 => n4846, A2 => n4845, A3 => n4844, A4 => 
                           n4843, ZN => n4852);
   U6578 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_71_port, B1 
                           => n5383, B2 => IF_Regsxreg_file_903_port, ZN => 
                           n4850);
   U6579 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_519_port, B1 
                           => n5361, B2 => IF_Regsxreg_file_135_port, ZN => 
                           n4849);
   U6580 : AOI22_X1 port map( A1 => n5278, A2 => IF_Regsxreg_file_391_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_647_port, ZN => 
                           n4848);
   U6581 : AOI22_X1 port map( A1 => n5413, A2 => IF_Regsxreg_file_263_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_7_port, ZN => n4847
                           );
   U6582 : NAND4_X1 port map( A1 => n4850, A2 => n4849, A3 => n4848, A4 => 
                           n4847, ZN => n4851);
   U6583 : AOI211_X1 port map( C1 => n4917, C2 => n4853, A => n4852, B => n4851
                           , ZN => n4854);
   U6584 : AOI21_X1 port map( B1 => n4855, B2 => n4854, A => n5216, ZN => 
                           IF_RegsxN634);
   U6585 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_488_port, B1 
                           => n5325, B2 => IF_Regsxreg_file_456_port, ZN => 
                           n4858);
   U6586 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_584_port, B1 
                           => n5400, B2 => IF_Regsxreg_file_360_port, ZN => 
                           n4857);
   U6587 : AOI22_X1 port map( A1 => n5399, A2 => IF_Regsxreg_file_328_port, B1 
                           => n5299, B2 => IF_Regsxreg_file_232_port, ZN => 
                           n4856);
   U6588 : NAND3_X1 port map( A1 => n4858, A2 => n4857, A3 => n4856, ZN => 
                           n4859);
   U6589 : AOI21_X1 port map( B1 => n5411, B2 => IF_Regsxreg_file_776_port, A 
                           => n4859, ZN => n4876);
   U6590 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_680_port, B1 
                           => n5293, B2 => IF_Regsxreg_file_424_port, ZN => 
                           n4863);
   U6591 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_168_port, B1 
                           => n5157, B2 => IF_Regsxreg_file_808_port, ZN => 
                           n4862);
   U6592 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_936_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_296_port, ZN => 
                           n4861);
   U6593 : AOI22_X1 port map( A1 => n5345, A2 => IF_Regsxreg_file_552_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_40_port, ZN => 
                           n4860);
   U6594 : NAND4_X1 port map( A1 => n4863, A2 => n4862, A3 => n4861, A4 => 
                           n4860, ZN => n4874);
   U6595 : AOI22_X1 port map( A1 => n5376, A2 => IF_Regsxreg_file_968_port, B1 
                           => n5273, B2 => IF_Regsxreg_file_744_port, ZN => 
                           n4867);
   U6596 : AOI22_X1 port map( A1 => n5314, A2 => IF_Regsxreg_file_840_port, B1 
                           => n5162, B2 => IF_Regsxreg_file_616_port, ZN => 
                           n4866);
   U6597 : AOI22_X1 port map( A1 => n5075, A2 => IF_Regsxreg_file_104_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_200_port, ZN => 
                           n4865);
   U6598 : AOI22_X1 port map( A1 => n5401, A2 => IF_Regsxreg_file_712_port, B1 
                           => n5300, B2 => IF_Regsxreg_file_872_port, ZN => 
                           n4864);
   U6599 : NAND4_X1 port map( A1 => n4867, A2 => n4866, A3 => n4865, A4 => 
                           n4864, ZN => n4873);
   U6600 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_72_port, B1 
                           => n5278, B2 => IF_Regsxreg_file_392_port, ZN => 
                           n4871);
   U6601 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_520_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_648_port, ZN => 
                           n4870);
   U6602 : AOI22_X1 port map( A1 => n5361, A2 => IF_Regsxreg_file_136_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_8_port, ZN => n4869
                           );
   U6603 : CLKBUF_X1 port map( A => n5383, Z => n5101);
   U6604 : AOI22_X1 port map( A1 => n5363, A2 => IF_Regsxreg_file_264_port, B1 
                           => n5101, B2 => IF_Regsxreg_file_904_port, ZN => 
                           n4868);
   U6605 : NAND4_X1 port map( A1 => n4871, A2 => n4870, A3 => n4869, A4 => 
                           n4868, ZN => n4872);
   U6606 : AOI211_X1 port map( C1 => n4917, C2 => n4874, A => n4873, B => n4872
                           , ZN => n4875);
   U6607 : AOI21_X1 port map( B1 => n4876, B2 => n4875, A => n5216, ZN => 
                           IF_RegsxN635);
   U6608 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_489_port, B1 
                           => n5325, B2 => IF_Regsxreg_file_457_port, ZN => 
                           n4879);
   U6609 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_585_port, B1 
                           => n5376, B2 => IF_Regsxreg_file_969_port, ZN => 
                           n4878);
   U6610 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_841_port, B1 
                           => n5162, B2 => IF_Regsxreg_file_617_port, ZN => 
                           n4877);
   U6611 : NAND3_X1 port map( A1 => n4879, A2 => n4878, A3 => n4877, ZN => 
                           n4880);
   U6612 : AOI21_X1 port map( B1 => n5415, B2 => IF_Regsxreg_file_521_port, A 
                           => n4880, ZN => n4897);
   U6613 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_937_port, B1 
                           => n5293, B2 => IF_Regsxreg_file_425_port, ZN => 
                           n4884);
   U6614 : AOI22_X1 port map( A1 => n5385, A2 => IF_Regsxreg_file_553_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_297_port, ZN => 
                           n4883);
   U6615 : AOI22_X1 port map( A1 => n5384, A2 => IF_Regsxreg_file_809_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_41_port, ZN => 
                           n4882);
   U6616 : AOI22_X1 port map( A1 => n5294, A2 => IF_Regsxreg_file_169_port, B1 
                           => n5320, B2 => IF_Regsxreg_file_681_port, ZN => 
                           n4881);
   U6617 : NAND4_X1 port map( A1 => n4884, A2 => n4883, A3 => n4882, A4 => 
                           n4881, ZN => n4895);
   U6618 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_105_port, B1 
                           => n5400, B2 => IF_Regsxreg_file_361_port, ZN => 
                           n4888);
   U6619 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_713_port, B1 
                           => n5240, B2 => IF_Regsxreg_file_73_port, ZN => 
                           n4887);
   U6620 : AOI22_X1 port map( A1 => n5399, A2 => IF_Regsxreg_file_329_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_201_port, ZN => 
                           n4886);
   U6621 : AOI22_X1 port map( A1 => n5299, A2 => IF_Regsxreg_file_233_port, B1 
                           => n5273, B2 => IF_Regsxreg_file_745_port, ZN => 
                           n4885);
   U6622 : NAND4_X1 port map( A1 => n4888, A2 => n4887, A3 => n4886, A4 => 
                           n4885, ZN => n4894);
   U6623 : AOI22_X1 port map( A1 => n5300, A2 => IF_Regsxreg_file_873_port, B1 
                           => n5101, B2 => IF_Regsxreg_file_905_port, ZN => 
                           n4892);
   U6624 : AOI22_X1 port map( A1 => n5361, A2 => IF_Regsxreg_file_137_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_649_port, ZN => 
                           n4891);
   U6625 : AOI22_X1 port map( A1 => n5411, A2 => IF_Regsxreg_file_777_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_9_port, ZN => n4890
                           );
   U6626 : AOI22_X1 port map( A1 => n5413, A2 => IF_Regsxreg_file_265_port, B1 
                           => n5278, B2 => IF_Regsxreg_file_393_port, ZN => 
                           n4889);
   U6627 : NAND4_X1 port map( A1 => n4892, A2 => n4891, A3 => n4890, A4 => 
                           n4889, ZN => n4893);
   U6628 : AOI211_X1 port map( C1 => n4917, C2 => n4895, A => n4894, B => n4893
                           , ZN => n4896);
   U6629 : AOI21_X1 port map( B1 => n4897, B2 => n4896, A => n5216, ZN => 
                           IF_RegsxN636);
   U6630 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_490_port, B1 
                           => n5325, B2 => IF_Regsxreg_file_458_port, ZN => 
                           n4900);
   U6631 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_106_port, B1 
                           => n5299, B2 => IF_Regsxreg_file_234_port, ZN => 
                           n4899);
   U6632 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_714_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_362_port, ZN => 
                           n4898);
   U6633 : NAND3_X1 port map( A1 => n4900, A2 => n4899, A3 => n4898, ZN => 
                           n4901);
   U6634 : AOI21_X1 port map( B1 => n5413, B2 => IF_Regsxreg_file_266_port, A 
                           => n4901, ZN => n4919);
   U6635 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_170_port, B1 
                           => n5320, B2 => IF_Regsxreg_file_682_port, ZN => 
                           n4905);
   U6636 : AOI22_X1 port map( A1 => n5385, A2 => IF_Regsxreg_file_554_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_42_port, ZN => 
                           n4904);
   U6637 : AOI22_X1 port map( A1 => n5384, A2 => IF_Regsxreg_file_810_port, B1 
                           => n5390, B2 => IF_Regsxreg_file_298_port, ZN => 
                           n4903);
   U6638 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_938_port, B1 
                           => n5293, B2 => IF_Regsxreg_file_426_port, ZN => 
                           n4902);
   U6639 : NAND4_X1 port map( A1 => n4905, A2 => n4904, A3 => n4903, A4 => 
                           n4902, ZN => n4916);
   U6640 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_586_port, B1 
                           => n5162, B2 => IF_Regsxreg_file_618_port, ZN => 
                           n4909);
   U6641 : AOI22_X1 port map( A1 => n5396, A2 => IF_Regsxreg_file_874_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_202_port, ZN => 
                           n4908);
   U6642 : AOI22_X1 port map( A1 => n5240, A2 => IF_Regsxreg_file_74_port, B1 
                           => n5399, B2 => IF_Regsxreg_file_330_port, ZN => 
                           n4907);
   U6643 : AOI22_X1 port map( A1 => n5314, A2 => IF_Regsxreg_file_842_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_746_port, ZN => 
                           n4906);
   U6644 : NAND4_X1 port map( A1 => n4909, A2 => n4908, A3 => n4907, A4 => 
                           n4906, ZN => n4915);
   U6645 : AOI22_X1 port map( A1 => n5376, A2 => IF_Regsxreg_file_970_port, B1 
                           => n5361, B2 => IF_Regsxreg_file_138_port, ZN => 
                           n4913);
   U6646 : AOI22_X1 port map( A1 => n5278, A2 => IF_Regsxreg_file_394_port, B1 
                           => n5101, B2 => IF_Regsxreg_file_906_port, ZN => 
                           n4912);
   U6647 : AOI22_X1 port map( A1 => n5411, A2 => IF_Regsxreg_file_778_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_650_port, ZN => 
                           n4911);
   U6648 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_522_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_10_port, ZN => 
                           n4910);
   U6649 : NAND4_X1 port map( A1 => n4913, A2 => n4912, A3 => n4911, A4 => 
                           n4910, ZN => n4914);
   U6650 : AOI211_X1 port map( C1 => n4917, C2 => n4916, A => n4915, B => n4914
                           , ZN => n4918);
   U6651 : AOI21_X1 port map( B1 => n4919, B2 => n4918, A => n5216, ZN => 
                           IF_RegsxN637);
   U6652 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_491_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_619_port, ZN => 
                           n4922);
   U6653 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_843_port, B1 
                           => n5264, B2 => IF_Regsxreg_file_971_port, ZN => 
                           n4921);
   U6654 : AOI22_X1 port map( A1 => n5300, A2 => IF_Regsxreg_file_875_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_363_port, ZN => 
                           n4920);
   U6655 : NAND3_X1 port map( A1 => n4922, A2 => n4921, A3 => n4920, ZN => 
                           n4923);
   U6656 : AOI21_X1 port map( B1 => n5278, B2 => IF_Regsxreg_file_395_port, A 
                           => n4923, ZN => n4940);
   U6657 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_683_port, B1 
                           => n5293, B2 => IF_Regsxreg_file_427_port, ZN => 
                           n4927);
   U6658 : AOI22_X1 port map( A1 => n5385, A2 => IF_Regsxreg_file_555_port, B1 
                           => n5157, B2 => IF_Regsxreg_file_811_port, ZN => 
                           n4926);
   U6659 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_939_port, B1 
                           => n5388, B2 => IF_Regsxreg_file_43_port, ZN => 
                           n4925);
   U6660 : AOI22_X1 port map( A1 => n5294, A2 => IF_Regsxreg_file_171_port, B1 
                           => n5390, B2 => IF_Regsxreg_file_299_port, ZN => 
                           n4924);
   U6661 : NAND4_X1 port map( A1 => n4927, A2 => n4926, A3 => n4925, A4 => 
                           n4924, ZN => n4938);
   U6662 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_715_port, B1 
                           => n5354, B2 => IF_Regsxreg_file_331_port, ZN => 
                           n4931);
   U6663 : AOI22_X1 port map( A1 => n5250, A2 => IF_Regsxreg_file_587_port, B1 
                           => n5299, B2 => IF_Regsxreg_file_235_port, ZN => 
                           n4930);
   U6664 : AOI22_X1 port map( A1 => n5075, A2 => IF_Regsxreg_file_107_port, B1 
                           => n5398, B2 => IF_Regsxreg_file_203_port, ZN => 
                           n4929);
   U6665 : AOI22_X1 port map( A1 => n5240, A2 => IF_Regsxreg_file_75_port, B1 
                           => n5325, B2 => IF_Regsxreg_file_459_port, ZN => 
                           n4928);
   U6666 : NAND4_X1 port map( A1 => n4931, A2 => n4930, A3 => n4929, A4 => 
                           n4928, ZN => n4937);
   U6667 : AOI22_X1 port map( A1 => n5402, A2 => IF_Regsxreg_file_747_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_11_port, ZN => 
                           n4935);
   U6668 : AOI22_X1 port map( A1 => n5413, A2 => IF_Regsxreg_file_267_port, B1 
                           => n5101, B2 => IF_Regsxreg_file_907_port, ZN => 
                           n4934);
   U6669 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_523_port, B1 
                           => n5361, B2 => IF_Regsxreg_file_139_port, ZN => 
                           n4933);
   U6670 : AOI22_X1 port map( A1 => n5411, A2 => IF_Regsxreg_file_779_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_651_port, ZN => 
                           n4932);
   U6671 : NAND4_X1 port map( A1 => n4935, A2 => n4934, A3 => n4933, A4 => 
                           n4932, ZN => n4936);
   U6672 : AOI211_X1 port map( C1 => n6266, C2 => n4938, A => n4937, B => n4936
                           , ZN => n4939);
   U6673 : AOI21_X1 port map( B1 => n4940, B2 => n4939, A => n5216, ZN => 
                           IF_RegsxN638);
   U6674 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_492_port, B1 
                           => n5376, B2 => IF_Regsxreg_file_972_port, ZN => 
                           n4943);
   U6675 : AOI22_X1 port map( A1 => n5353, A2 => IF_Regsxreg_file_204_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_620_port, ZN => 
                           n4942);
   U6676 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_76_port, B1 
                           => n5300, B2 => IF_Regsxreg_file_876_port, ZN => 
                           n4941);
   U6677 : NAND3_X1 port map( A1 => n4943, A2 => n4942, A3 => n4941, ZN => 
                           n4944);
   U6678 : AOI21_X1 port map( B1 => n5415, B2 => IF_Regsxreg_file_524_port, A 
                           => n4944, ZN => n4961);
   U6679 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_172_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_44_port, ZN => 
                           n4948);
   U6680 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_940_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_300_port, ZN => 
                           n4947);
   U6681 : AOI22_X1 port map( A1 => n5345, A2 => IF_Regsxreg_file_556_port, B1 
                           => n5293, B2 => IF_Regsxreg_file_428_port, ZN => 
                           n4946);
   U6682 : AOI22_X1 port map( A1 => n5391, A2 => IF_Regsxreg_file_684_port, B1 
                           => n5157, B2 => IF_Regsxreg_file_812_port, ZN => 
                           n4945);
   U6683 : NAND4_X1 port map( A1 => n4948, A2 => n4947, A3 => n4946, A4 => 
                           n4945, ZN => n4959);
   U6684 : AOI22_X1 port map( A1 => n5399, A2 => IF_Regsxreg_file_332_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_748_port, ZN => 
                           n4952);
   U6685 : AOI22_X1 port map( A1 => n5250, A2 => IF_Regsxreg_file_588_port, B1 
                           => n5325, B2 => IF_Regsxreg_file_460_port, ZN => 
                           n4951);
   U6686 : AOI22_X1 port map( A1 => n5314, A2 => IF_Regsxreg_file_844_port, B1 
                           => n5400, B2 => IF_Regsxreg_file_364_port, ZN => 
                           n4950);
   U6687 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_716_port, B1 
                           => n5075, B2 => IF_Regsxreg_file_108_port, ZN => 
                           n4949);
   U6688 : NAND4_X1 port map( A1 => n4952, A2 => n4951, A3 => n4950, A4 => 
                           n4949, ZN => n4958);
   U6689 : AOI22_X1 port map( A1 => n5377, A2 => IF_Regsxreg_file_236_port, B1 
                           => n5278, B2 => IF_Regsxreg_file_396_port, ZN => 
                           n4956);
   U6690 : AOI22_X1 port map( A1 => n5363, A2 => IF_Regsxreg_file_268_port, B1 
                           => n5101, B2 => IF_Regsxreg_file_908_port, ZN => 
                           n4955);
   U6691 : AOI22_X1 port map( A1 => n5279, A2 => IF_Regsxreg_file_780_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_12_port, ZN => 
                           n4954);
   U6692 : AOI22_X1 port map( A1 => n5361, A2 => IF_Regsxreg_file_140_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_652_port, ZN => 
                           n4953);
   U6693 : NAND4_X1 port map( A1 => n4956, A2 => n4955, A3 => n4954, A4 => 
                           n4953, ZN => n4957);
   U6694 : AOI211_X1 port map( C1 => n6266, C2 => n4959, A => n4958, B => n4957
                           , ZN => n4960);
   U6695 : AOI21_X1 port map( B1 => n4961, B2 => n4960, A => n5216, ZN => 
                           IF_RegsxN639);
   U6696 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_493_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_621_port, ZN => 
                           n4964);
   U6697 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_845_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_749_port, ZN => 
                           n4963);
   U6698 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_109_port, B1 
                           => n5354, B2 => IF_Regsxreg_file_333_port, ZN => 
                           n4962);
   U6699 : NAND3_X1 port map( A1 => n4964, A2 => n4963, A3 => n4962, ZN => 
                           n4965);
   U6700 : AOI21_X1 port map( B1 => n5362, B2 => IF_Regsxreg_file_13_port, A =>
                           n4965, ZN => n4982);
   U6701 : AOI22_X1 port map( A1 => n5384, A2 => IF_Regsxreg_file_813_port, B1 
                           => n5386, B2 => IF_Regsxreg_file_429_port, ZN => 
                           n4969);
   U6702 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_941_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_301_port, ZN => 
                           n4968);
   U6703 : AOI22_X1 port map( A1 => n5391, A2 => IF_Regsxreg_file_685_port, B1 
                           => n5385, B2 => IF_Regsxreg_file_557_port, ZN => 
                           n4967);
   U6704 : AOI22_X1 port map( A1 => n5294, A2 => IF_Regsxreg_file_173_port, B1 
                           => n5388, B2 => IF_Regsxreg_file_45_port, ZN => 
                           n4966);
   U6705 : NAND4_X1 port map( A1 => n4969, A2 => n4968, A3 => n4967, A4 => 
                           n4966, ZN => n4980);
   U6706 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_717_port, B1 
                           => n5300, B2 => IF_Regsxreg_file_877_port, ZN => 
                           n4973);
   U6707 : AOI22_X1 port map( A1 => n5250, A2 => IF_Regsxreg_file_589_port, B1 
                           => n5352, B2 => IF_Regsxreg_file_973_port, ZN => 
                           n4972);
   U6708 : AOI22_X1 port map( A1 => n5240, A2 => IF_Regsxreg_file_77_port, B1 
                           => n5398, B2 => IF_Regsxreg_file_205_port, ZN => 
                           n4971);
   U6709 : AOI22_X1 port map( A1 => n5373, A2 => IF_Regsxreg_file_461_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_237_port, ZN => 
                           n4970);
   U6710 : NAND4_X1 port map( A1 => n4973, A2 => n4972, A3 => n4971, A4 => 
                           n4970, ZN => n4979);
   U6711 : AOI22_X1 port map( A1 => n5279, A2 => IF_Regsxreg_file_781_port, B1 
                           => n5400, B2 => IF_Regsxreg_file_365_port, ZN => 
                           n4977);
   U6712 : AOI22_X1 port map( A1 => n5361, A2 => IF_Regsxreg_file_141_port, B1 
                           => n5101, B2 => IF_Regsxreg_file_909_port, ZN => 
                           n4976);
   U6713 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_525_port, B1 
                           => n5363, B2 => IF_Regsxreg_file_269_port, ZN => 
                           n4975);
   U6714 : AOI22_X1 port map( A1 => n5278, A2 => IF_Regsxreg_file_397_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_653_port, ZN => 
                           n4974);
   U6715 : NAND4_X1 port map( A1 => n4977, A2 => n4976, A3 => n4975, A4 => 
                           n4974, ZN => n4978);
   U6716 : AOI211_X1 port map( C1 => n6266, C2 => n4980, A => n4979, B => n4978
                           , ZN => n4981);
   U6717 : AOI21_X1 port map( B1 => n4982, B2 => n4981, A => n5216, ZN => 
                           IF_RegsxN640);
   U6718 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_494_port, B1 
                           => n5401, B2 => IF_Regsxreg_file_718_port, ZN => 
                           n4985);
   U6719 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_846_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_750_port, ZN => 
                           n4984);
   U6720 : AOI22_X1 port map( A1 => n5300, A2 => IF_Regsxreg_file_878_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_366_port, ZN => 
                           n4983);
   U6721 : NAND3_X1 port map( A1 => n4985, A2 => n4984, A3 => n4983, ZN => 
                           n4986);
   U6722 : AOI21_X1 port map( B1 => n5415, B2 => IF_Regsxreg_file_526_port, A 
                           => n4986, ZN => n5003);
   U6723 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_174_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_302_port, ZN => 
                           n4990);
   U6724 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_942_port, B1 
                           => n5157, B2 => IF_Regsxreg_file_814_port, ZN => 
                           n4989);
   U6725 : AOI22_X1 port map( A1 => n5345, A2 => IF_Regsxreg_file_558_port, B1 
                           => n5388, B2 => IF_Regsxreg_file_46_port, ZN => 
                           n4988);
   U6726 : AOI22_X1 port map( A1 => n5391, A2 => IF_Regsxreg_file_686_port, B1 
                           => n5293, B2 => IF_Regsxreg_file_430_port, ZN => 
                           n4987);
   U6727 : NAND4_X1 port map( A1 => n4990, A2 => n4989, A3 => n4988, A4 => 
                           n4987, ZN => n5001);
   U6728 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_110_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_206_port, ZN => 
                           n4994);
   U6729 : AOI22_X1 port map( A1 => n5352, A2 => IF_Regsxreg_file_974_port, B1 
                           => n5325, B2 => IF_Regsxreg_file_462_port, ZN => 
                           n4993);
   U6730 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_78_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_238_port, ZN => 
                           n4992);
   U6731 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_590_port, B1 
                           => n5399, B2 => IF_Regsxreg_file_334_port, ZN => 
                           n4991);
   U6732 : NAND4_X1 port map( A1 => n4994, A2 => n4993, A3 => n4992, A4 => 
                           n4991, ZN => n5000);
   U6733 : AOI22_X1 port map( A1 => n5375, A2 => IF_Regsxreg_file_622_port, B1 
                           => n5411, B2 => IF_Regsxreg_file_782_port, ZN => 
                           n4998);
   U6734 : AOI22_X1 port map( A1 => n5361, A2 => IF_Regsxreg_file_142_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_14_port, ZN => 
                           n4997);
   U6735 : AOI22_X1 port map( A1 => n5278, A2 => IF_Regsxreg_file_398_port, B1 
                           => n5101, B2 => IF_Regsxreg_file_910_port, ZN => 
                           n4996);
   U6736 : AOI22_X1 port map( A1 => n5363, A2 => IF_Regsxreg_file_270_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_654_port, ZN => 
                           n4995);
   U6737 : NAND4_X1 port map( A1 => n4998, A2 => n4997, A3 => n4996, A4 => 
                           n4995, ZN => n4999);
   U6738 : AOI211_X1 port map( C1 => n6266, C2 => n5001, A => n5000, B => n4999
                           , ZN => n5002);
   U6739 : AOI21_X1 port map( B1 => n5003, B2 => n5002, A => n5216, ZN => 
                           IF_RegsxN641);
   U6740 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_495_port, B1 
                           => n5075, B2 => IF_Regsxreg_file_111_port, ZN => 
                           n5006);
   U6741 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_591_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_623_port, ZN => 
                           n5005);
   U6742 : AOI22_X1 port map( A1 => n5300, A2 => IF_Regsxreg_file_879_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_207_port, ZN => 
                           n5004);
   U6743 : NAND3_X1 port map( A1 => n5006, A2 => n5005, A3 => n5004, ZN => 
                           n5007);
   U6744 : AOI21_X1 port map( B1 => n5413, B2 => IF_Regsxreg_file_271_port, A 
                           => n5007, ZN => n5024);
   U6745 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_687_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_47_port, ZN => 
                           n5011);
   U6746 : AOI22_X1 port map( A1 => n5385, A2 => IF_Regsxreg_file_559_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_303_port, ZN => 
                           n5010);
   U6747 : AOI22_X1 port map( A1 => n5294, A2 => IF_Regsxreg_file_175_port, B1 
                           => n5245, B2 => IF_Regsxreg_file_943_port, ZN => 
                           n5009);
   U6748 : AOI22_X1 port map( A1 => n5157, A2 => IF_Regsxreg_file_815_port, B1 
                           => n5386, B2 => IF_Regsxreg_file_431_port, ZN => 
                           n5008);
   U6749 : NAND4_X1 port map( A1 => n5011, A2 => n5010, A3 => n5009, A4 => 
                           n5008, ZN => n5022);
   U6750 : AOI22_X1 port map( A1 => n5352, A2 => IF_Regsxreg_file_975_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_751_port, ZN => 
                           n5015);
   U6751 : AOI22_X1 port map( A1 => n5401, A2 => IF_Regsxreg_file_719_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_239_port, ZN => 
                           n5014);
   U6752 : AOI22_X1 port map( A1 => n5240, A2 => IF_Regsxreg_file_79_port, B1 
                           => n5354, B2 => IF_Regsxreg_file_335_port, ZN => 
                           n5013);
   U6753 : AOI22_X1 port map( A1 => n5373, A2 => IF_Regsxreg_file_463_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_367_port, ZN => 
                           n5012);
   U6754 : NAND4_X1 port map( A1 => n5015, A2 => n5014, A3 => n5013, A4 => 
                           n5012, ZN => n5021);
   U6755 : AOI22_X1 port map( A1 => n5314, A2 => IF_Regsxreg_file_847_port, B1 
                           => n5414, B2 => IF_Regsxreg_file_399_port, ZN => 
                           n5019);
   U6756 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_527_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_655_port, ZN => 
                           n5018);
   U6757 : AOI22_X1 port map( A1 => n5279, A2 => IF_Regsxreg_file_783_port, B1 
                           => n5361, B2 => IF_Regsxreg_file_143_port, ZN => 
                           n5017);
   U6758 : AOI22_X1 port map( A1 => n5362, A2 => IF_Regsxreg_file_15_port, B1 
                           => n5101, B2 => IF_Regsxreg_file_911_port, ZN => 
                           n5016);
   U6759 : NAND4_X1 port map( A1 => n5019, A2 => n5018, A3 => n5017, A4 => 
                           n5016, ZN => n5020);
   U6760 : AOI211_X1 port map( C1 => n6266, C2 => n5022, A => n5021, B => n5020
                           , ZN => n5023);
   U6761 : AOI21_X1 port map( B1 => n5024, B2 => n5023, A => n5216, ZN => 
                           IF_RegsxN642);
   U6762 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_496_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_752_port, ZN => 
                           n5027);
   U6763 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_80_port, B1 
                           => n5300, B2 => IF_Regsxreg_file_880_port, ZN => 
                           n5026);
   U6764 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_720_port, B1 
                           => n5314, B2 => IF_Regsxreg_file_848_port, ZN => 
                           n5025);
   U6765 : NAND3_X1 port map( A1 => n5027, A2 => n5026, A3 => n5025, ZN => 
                           n5028);
   U6766 : AOI21_X1 port map( B1 => n5413, B2 => IF_Regsxreg_file_272_port, A 
                           => n5028, ZN => n5045);
   U6767 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_688_port, B1 
                           => n5385, B2 => IF_Regsxreg_file_560_port, ZN => 
                           n5032);
   U6768 : AOI22_X1 port map( A1 => n5293, A2 => IF_Regsxreg_file_432_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_304_port, ZN => 
                           n5031);
   U6769 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_944_port, B1 
                           => n5388, B2 => IF_Regsxreg_file_48_port, ZN => 
                           n5030);
   U6770 : AOI22_X1 port map( A1 => n5294, A2 => IF_Regsxreg_file_176_port, B1 
                           => n5384, B2 => IF_Regsxreg_file_816_port, ZN => 
                           n5029);
   U6771 : NAND4_X1 port map( A1 => n5032, A2 => n5031, A3 => n5030, A4 => 
                           n5029, ZN => n5043);
   U6772 : AOI22_X1 port map( A1 => n5353, A2 => IF_Regsxreg_file_208_port, B1 
                           => n5162, B2 => IF_Regsxreg_file_624_port, ZN => 
                           n5036);
   U6773 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_112_port, B1 
                           => n5376, B2 => IF_Regsxreg_file_976_port, ZN => 
                           n5035);
   U6774 : AOI22_X1 port map( A1 => n5377, A2 => IF_Regsxreg_file_240_port, B1 
                           => n5400, B2 => IF_Regsxreg_file_368_port, ZN => 
                           n5034);
   U6775 : AOI22_X1 port map( A1 => n5354, A2 => IF_Regsxreg_file_336_port, B1 
                           => n5325, B2 => IF_Regsxreg_file_464_port, ZN => 
                           n5033);
   U6776 : NAND4_X1 port map( A1 => n5036, A2 => n5035, A3 => n5034, A4 => 
                           n5033, ZN => n5042);
   U6777 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_592_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_16_port, ZN => 
                           n5040);
   U6778 : AOI22_X1 port map( A1 => n5279, A2 => IF_Regsxreg_file_784_port, B1 
                           => n5361, B2 => IF_Regsxreg_file_144_port, ZN => 
                           n5039);
   U6779 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_528_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_656_port, ZN => 
                           n5038);
   U6780 : AOI22_X1 port map( A1 => n5278, A2 => IF_Regsxreg_file_400_port, B1 
                           => n5101, B2 => IF_Regsxreg_file_912_port, ZN => 
                           n5037);
   U6781 : NAND4_X1 port map( A1 => n5040, A2 => n5039, A3 => n5038, A4 => 
                           n5037, ZN => n5041);
   U6782 : AOI211_X1 port map( C1 => n6266, C2 => n5043, A => n5042, B => n5041
                           , ZN => n5044);
   U6783 : AOI21_X1 port map( B1 => n5045, B2 => n5044, A => n5216, ZN => 
                           IF_RegsxN643);
   U6784 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_497_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_625_port, ZN => 
                           n5048);
   U6785 : AOI22_X1 port map( A1 => n5352, A2 => IF_Regsxreg_file_977_port, B1 
                           => n5300, B2 => IF_Regsxreg_file_881_port, ZN => 
                           n5047);
   U6786 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_593_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_753_port, ZN => 
                           n5046);
   U6787 : NAND3_X1 port map( A1 => n5048, A2 => n5047, A3 => n5046, ZN => 
                           n5049);
   U6788 : AOI21_X1 port map( B1 => n5362, B2 => IF_Regsxreg_file_17_port, A =>
                           n5049, ZN => n5066);
   U6789 : AOI22_X1 port map( A1 => n5384, A2 => IF_Regsxreg_file_817_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_305_port, ZN => 
                           n5053);
   U6790 : AOI22_X1 port map( A1 => n5294, A2 => IF_Regsxreg_file_177_port, B1 
                           => n5386, B2 => IF_Regsxreg_file_433_port, ZN => 
                           n5052);
   U6791 : AOI22_X1 port map( A1 => n5391, A2 => IF_Regsxreg_file_689_port, B1 
                           => n5385, B2 => IF_Regsxreg_file_561_port, ZN => 
                           n5051);
   U6792 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_945_port, B1 
                           => n5388, B2 => IF_Regsxreg_file_49_port, ZN => 
                           n5050);
   U6793 : NAND4_X1 port map( A1 => n5053, A2 => n5052, A3 => n5051, A4 => 
                           n5050, ZN => n5064);
   U6794 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_721_port, B1 
                           => n5354, B2 => IF_Regsxreg_file_337_port, ZN => 
                           n5057);
   U6795 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_113_port, B1 
                           => n5378, B2 => IF_Regsxreg_file_81_port, ZN => 
                           n5056);
   U6796 : AOI22_X1 port map( A1 => n5377, A2 => IF_Regsxreg_file_241_port, B1 
                           => n5398, B2 => IF_Regsxreg_file_209_port, ZN => 
                           n5055);
   U6797 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_849_port, B1 
                           => n5325, B2 => IF_Regsxreg_file_465_port, ZN => 
                           n5054);
   U6798 : NAND4_X1 port map( A1 => n5057, A2 => n5056, A3 => n5055, A4 => 
                           n5054, ZN => n5063);
   U6799 : AOI22_X1 port map( A1 => n5351, A2 => IF_Regsxreg_file_369_port, B1 
                           => n5101, B2 => IF_Regsxreg_file_913_port, ZN => 
                           n5061);
   U6800 : AOI22_X1 port map( A1 => n5363, A2 => IF_Regsxreg_file_273_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_657_port, ZN => 
                           n5060);
   U6801 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_529_port, B1 
                           => n5411, B2 => IF_Regsxreg_file_785_port, ZN => 
                           n5059);
   U6802 : AOI22_X1 port map( A1 => n5361, A2 => IF_Regsxreg_file_145_port, B1 
                           => n5414, B2 => IF_Regsxreg_file_401_port, ZN => 
                           n5058);
   U6803 : NAND4_X1 port map( A1 => n5061, A2 => n5060, A3 => n5059, A4 => 
                           n5058, ZN => n5062);
   U6804 : AOI211_X1 port map( C1 => n6266, C2 => n5064, A => n5063, B => n5062
                           , ZN => n5065);
   U6805 : AOI21_X1 port map( B1 => n5066, B2 => n5065, A => n5216, ZN => 
                           IF_RegsxN644);
   U6806 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_498_port, B1 
                           => n5325, B2 => IF_Regsxreg_file_466_port, ZN => 
                           n5069);
   U6807 : AOI22_X1 port map( A1 => n5352, A2 => IF_Regsxreg_file_978_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_210_port, ZN => 
                           n5068);
   U6808 : AOI22_X1 port map( A1 => n5377, A2 => IF_Regsxreg_file_242_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_370_port, ZN => 
                           n5067);
   U6809 : NAND3_X1 port map( A1 => n5069, A2 => n5068, A3 => n5067, ZN => 
                           n5070);
   U6810 : AOI21_X1 port map( B1 => n5414, B2 => IF_Regsxreg_file_402_port, A 
                           => n5070, ZN => n5088);
   U6811 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_178_port, B1 
                           => n5157, B2 => IF_Regsxreg_file_818_port, ZN => 
                           n5074);
   U6812 : AOI22_X1 port map( A1 => n5385, A2 => IF_Regsxreg_file_562_port, B1 
                           => n5245, B2 => IF_Regsxreg_file_946_port, ZN => 
                           n5073);
   U6813 : AOI22_X1 port map( A1 => n5293, A2 => IF_Regsxreg_file_434_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_306_port, ZN => 
                           n5072);
   U6814 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_690_port, B1 
                           => n5388, B2 => IF_Regsxreg_file_50_port, ZN => 
                           n5071);
   U6815 : NAND4_X1 port map( A1 => n5074, A2 => n5073, A3 => n5072, A4 => 
                           n5071, ZN => n5086);
   U6816 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_594_port, B1 
                           => n5300, B2 => IF_Regsxreg_file_882_port, ZN => 
                           n5079);
   U6817 : AOI22_X1 port map( A1 => n5240, A2 => IF_Regsxreg_file_82_port, B1 
                           => n5399, B2 => IF_Regsxreg_file_338_port, ZN => 
                           n5078);
   U6818 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_722_port, B1 
                           => n5162, B2 => IF_Regsxreg_file_626_port, ZN => 
                           n5077);
   U6819 : AOI22_X1 port map( A1 => n5075, A2 => IF_Regsxreg_file_114_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_754_port, ZN => 
                           n5076);
   U6820 : NAND4_X1 port map( A1 => n5079, A2 => n5078, A3 => n5077, A4 => 
                           n5076, ZN => n5085);
   U6821 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_850_port, B1 
                           => n5411, B2 => IF_Regsxreg_file_786_port, ZN => 
                           n5083);
   U6822 : AOI22_X1 port map( A1 => n5412, A2 => IF_Regsxreg_file_146_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_658_port, ZN => 
                           n5082);
   U6823 : CLKBUF_X1 port map( A => n5415, Z => n5359);
   U6824 : AOI22_X1 port map( A1 => n5359, A2 => IF_Regsxreg_file_530_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_18_port, ZN => 
                           n5081);
   U6825 : AOI22_X1 port map( A1 => n5363, A2 => IF_Regsxreg_file_274_port, B1 
                           => n5101, B2 => IF_Regsxreg_file_914_port, ZN => 
                           n5080);
   U6826 : NAND4_X1 port map( A1 => n5083, A2 => n5082, A3 => n5081, A4 => 
                           n5080, ZN => n5084);
   U6827 : AOI211_X1 port map( C1 => n6266, C2 => n5086, A => n5085, B => n5084
                           , ZN => n5087);
   U6828 : AOI21_X1 port map( B1 => n5088, B2 => n5087, A => n5216, ZN => 
                           IF_RegsxN645);
   U6829 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_499_port, B1 
                           => n5399, B2 => IF_Regsxreg_file_339_port, ZN => 
                           n5091);
   U6830 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_723_port, B1 
                           => n5314, B2 => IF_Regsxreg_file_851_port, ZN => 
                           n5090);
   U6831 : AOI22_X1 port map( A1 => n5402, A2 => IF_Regsxreg_file_755_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_371_port, ZN => 
                           n5089);
   U6832 : NAND3_X1 port map( A1 => n5091, A2 => n5090, A3 => n5089, ZN => 
                           n5092);
   U6833 : AOI21_X1 port map( B1 => n5412, B2 => IF_Regsxreg_file_147_port, A 
                           => n5092, ZN => n5110);
   U6834 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_179_port, B1 
                           => n5245, B2 => IF_Regsxreg_file_947_port, ZN => 
                           n5096);
   U6835 : AOI22_X1 port map( A1 => n5345, A2 => IF_Regsxreg_file_563_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_307_port, ZN => 
                           n5095);
   U6836 : AOI22_X1 port map( A1 => n5384, A2 => IF_Regsxreg_file_819_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_51_port, ZN => 
                           n5094);
   U6837 : AOI22_X1 port map( A1 => n5391, A2 => IF_Regsxreg_file_691_port, B1 
                           => n5293, B2 => IF_Regsxreg_file_435_port, ZN => 
                           n5093);
   U6838 : NAND4_X1 port map( A1 => n5096, A2 => n5095, A3 => n5094, A4 => 
                           n5093, ZN => n5108);
   U6839 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_83_port, B1 
                           => n5250, B2 => IF_Regsxreg_file_595_port, ZN => 
                           n5100);
   U6840 : AOI22_X1 port map( A1 => n5373, A2 => IF_Regsxreg_file_467_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_243_port, ZN => 
                           n5099);
   U6841 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_115_port, B1 
                           => n5300, B2 => IF_Regsxreg_file_883_port, ZN => 
                           n5098);
   U6842 : AOI22_X1 port map( A1 => n5352, A2 => IF_Regsxreg_file_979_port, B1 
                           => n5162, B2 => IF_Regsxreg_file_627_port, ZN => 
                           n5097);
   U6843 : NAND4_X1 port map( A1 => n5100, A2 => n5099, A3 => n5098, A4 => 
                           n5097, ZN => n5107);
   U6844 : AOI22_X1 port map( A1 => n5353, A2 => IF_Regsxreg_file_211_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_659_port, ZN => 
                           n5105);
   U6845 : AOI22_X1 port map( A1 => n5363, A2 => IF_Regsxreg_file_275_port, B1 
                           => n5414, B2 => IF_Regsxreg_file_403_port, ZN => 
                           n5104);
   U6846 : AOI22_X1 port map( A1 => n5279, A2 => IF_Regsxreg_file_787_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_19_port, ZN => 
                           n5103);
   U6847 : AOI22_X1 port map( A1 => n5359, A2 => IF_Regsxreg_file_531_port, B1 
                           => n5101, B2 => IF_Regsxreg_file_915_port, ZN => 
                           n5102);
   U6848 : NAND4_X1 port map( A1 => n5105, A2 => n5104, A3 => n5103, A4 => 
                           n5102, ZN => n5106);
   U6849 : AOI211_X1 port map( C1 => n6266, C2 => n5108, A => n5107, B => n5106
                           , ZN => n5109);
   U6850 : AOI21_X1 port map( B1 => n5110, B2 => n5109, A => n5216, ZN => 
                           IF_RegsxN646);
   U6851 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_500_port, B1 
                           => n5376, B2 => IF_Regsxreg_file_980_port, ZN => 
                           n5113);
   U6852 : AOI22_X1 port map( A1 => n5300, A2 => IF_Regsxreg_file_884_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_244_port, ZN => 
                           n5112);
   U6853 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_116_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_372_port, ZN => 
                           n5111);
   U6854 : NAND3_X1 port map( A1 => n5113, A2 => n5112, A3 => n5111, ZN => 
                           n5114);
   U6855 : AOI21_X1 port map( B1 => n5415, B2 => IF_Regsxreg_file_532_port, A 
                           => n5114, ZN => n5131);
   U6856 : AOI22_X1 port map( A1 => n5385, A2 => IF_Regsxreg_file_564_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_52_port, ZN => 
                           n5118);
   U6857 : AOI22_X1 port map( A1 => n5294, A2 => IF_Regsxreg_file_180_port, B1 
                           => n5320, B2 => IF_Regsxreg_file_692_port, ZN => 
                           n5117);
   U6858 : AOI22_X1 port map( A1 => n5386, A2 => IF_Regsxreg_file_436_port, B1 
                           => n5390, B2 => IF_Regsxreg_file_308_port, ZN => 
                           n5116);
   U6859 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_948_port, B1 
                           => n5384, B2 => IF_Regsxreg_file_820_port, ZN => 
                           n5115);
   U6860 : NAND4_X1 port map( A1 => n5118, A2 => n5117, A3 => n5116, A4 => 
                           n5115, ZN => n5129);
   U6861 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_84_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_212_port, ZN => 
                           n5122);
   U6862 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_724_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_756_port, ZN => 
                           n5121);
   U6863 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_596_port, B1 
                           => n5325, B2 => IF_Regsxreg_file_468_port, ZN => 
                           n5120);
   U6864 : AOI22_X1 port map( A1 => n5354, A2 => IF_Regsxreg_file_340_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_628_port, ZN => 
                           n5119);
   U6865 : NAND4_X1 port map( A1 => n5122, A2 => n5121, A3 => n5120, A4 => 
                           n5119, ZN => n5128);
   U6866 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_852_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_20_port, ZN => 
                           n5126);
   U6867 : AOI22_X1 port map( A1 => n5279, A2 => IF_Regsxreg_file_788_port, B1 
                           => n5413, B2 => IF_Regsxreg_file_276_port, ZN => 
                           n5125);
   U6868 : AOI22_X1 port map( A1 => n5412, A2 => IF_Regsxreg_file_148_port, B1 
                           => n5414, B2 => IF_Regsxreg_file_404_port, ZN => 
                           n5124);
   U6869 : AOI22_X1 port map( A1 => n5383, A2 => IF_Regsxreg_file_916_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_660_port, ZN => 
                           n5123);
   U6870 : NAND4_X1 port map( A1 => n5126, A2 => n5125, A3 => n5124, A4 => 
                           n5123, ZN => n5127);
   U6871 : AOI211_X1 port map( C1 => n6266, C2 => n5129, A => n5128, B => n5127
                           , ZN => n5130);
   U6872 : AOI21_X1 port map( B1 => n5131, B2 => n5130, A => n5216, ZN => 
                           IF_RegsxN647);
   U6873 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_501_port, B1 
                           => n5399, B2 => IF_Regsxreg_file_341_port, ZN => 
                           n5134);
   U6874 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_117_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_757_port, ZN => 
                           n5133);
   U6875 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_725_port, B1 
                           => n5162, B2 => IF_Regsxreg_file_629_port, ZN => 
                           n5132);
   U6876 : NAND3_X1 port map( A1 => n5134, A2 => n5133, A3 => n5132, ZN => 
                           n5135);
   U6877 : AOI21_X1 port map( B1 => n5411, B2 => IF_Regsxreg_file_789_port, A 
                           => n5135, ZN => n5152);
   U6878 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_693_port, B1 
                           => n5157, B2 => IF_Regsxreg_file_821_port, ZN => 
                           n5139);
   U6879 : AOI22_X1 port map( A1 => n5293, A2 => IF_Regsxreg_file_437_port, B1 
                           => n5390, B2 => IF_Regsxreg_file_309_port, ZN => 
                           n5138);
   U6880 : AOI22_X1 port map( A1 => n5345, A2 => IF_Regsxreg_file_565_port, B1 
                           => n5388, B2 => IF_Regsxreg_file_53_port, ZN => 
                           n5137);
   U6881 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_181_port, B1 
                           => n5245, B2 => IF_Regsxreg_file_949_port, ZN => 
                           n5136);
   U6882 : NAND4_X1 port map( A1 => n5139, A2 => n5138, A3 => n5137, A4 => 
                           n5136, ZN => n5150);
   U6883 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_85_port, B1 
                           => n5373, B2 => IF_Regsxreg_file_469_port, ZN => 
                           n5143);
   U6884 : AOI22_X1 port map( A1 => n5396, A2 => IF_Regsxreg_file_885_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_373_port, ZN => 
                           n5142);
   U6885 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_853_port, B1 
                           => n5376, B2 => IF_Regsxreg_file_981_port, ZN => 
                           n5141);
   U6886 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_597_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_245_port, ZN => 
                           n5140);
   U6887 : NAND4_X1 port map( A1 => n5143, A2 => n5142, A3 => n5141, A4 => 
                           n5140, ZN => n5149);
   U6888 : AOI22_X1 port map( A1 => n5353, A2 => IF_Regsxreg_file_213_port, B1 
                           => n5412, B2 => IF_Regsxreg_file_149_port, ZN => 
                           n5147);
   U6889 : AOI22_X1 port map( A1 => n5359, A2 => IF_Regsxreg_file_533_port, B1 
                           => n5363, B2 => IF_Regsxreg_file_277_port, ZN => 
                           n5146);
   U6890 : AOI22_X1 port map( A1 => n5383, A2 => IF_Regsxreg_file_917_port, B1 
                           => n5360, B2 => IF_Regsxreg_file_661_port, ZN => 
                           n5145);
   U6891 : AOI22_X1 port map( A1 => n5278, A2 => IF_Regsxreg_file_405_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_21_port, ZN => 
                           n5144);
   U6892 : NAND4_X1 port map( A1 => n5147, A2 => n5146, A3 => n5145, A4 => 
                           n5144, ZN => n5148);
   U6893 : AOI211_X1 port map( C1 => n6266, C2 => n5150, A => n5149, B => n5148
                           , ZN => n5151);
   U6894 : AOI21_X1 port map( B1 => n5152, B2 => n5151, A => n5216, ZN => 
                           IF_RegsxN648);
   U6895 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_502_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_758_port, ZN => 
                           n5155);
   U6896 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_118_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_246_port, ZN => 
                           n5154);
   U6897 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_854_port, B1 
                           => n5396, B2 => IF_Regsxreg_file_886_port, ZN => 
                           n5153);
   U6898 : NAND3_X1 port map( A1 => n5155, A2 => n5154, A3 => n5153, ZN => 
                           n5156);
   U6899 : AOI21_X1 port map( B1 => n5413, B2 => IF_Regsxreg_file_278_port, A 
                           => n5156, ZN => n5175);
   U6900 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_182_port, B1 
                           => n5157, B2 => IF_Regsxreg_file_822_port, ZN => 
                           n5161);
   U6901 : AOI22_X1 port map( A1 => n5345, A2 => IF_Regsxreg_file_566_port, B1 
                           => n5389, B2 => IF_Regsxreg_file_950_port, ZN => 
                           n5160);
   U6902 : AOI22_X1 port map( A1 => n5293, A2 => IF_Regsxreg_file_438_port, B1 
                           => n5390, B2 => IF_Regsxreg_file_310_port, ZN => 
                           n5159);
   U6903 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_694_port, B1 
                           => n5388, B2 => IF_Regsxreg_file_54_port, ZN => 
                           n5158);
   U6904 : NAND4_X1 port map( A1 => n5161, A2 => n5160, A3 => n5159, A4 => 
                           n5158, ZN => n5173);
   U6905 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_86_port, B1 
                           => n5352, B2 => IF_Regsxreg_file_982_port, ZN => 
                           n5166);
   U6906 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_726_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_374_port, ZN => 
                           n5165);
   U6907 : AOI22_X1 port map( A1 => n5399, A2 => IF_Regsxreg_file_342_port, B1 
                           => n5398, B2 => IF_Regsxreg_file_214_port, ZN => 
                           n5164);
   U6908 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_598_port, B1 
                           => n5162, B2 => IF_Regsxreg_file_630_port, ZN => 
                           n5163);
   U6909 : NAND4_X1 port map( A1 => n5166, A2 => n5165, A3 => n5164, A4 => 
                           n5163, ZN => n5172);
   U6910 : AOI22_X1 port map( A1 => n5325, A2 => IF_Regsxreg_file_470_port, B1 
                           => n5383, B2 => IF_Regsxreg_file_918_port, ZN => 
                           n5170);
   U6911 : AOI22_X1 port map( A1 => n5359, A2 => IF_Regsxreg_file_534_port, B1 
                           => n5411, B2 => IF_Regsxreg_file_790_port, ZN => 
                           n5169);
   U6912 : AOI22_X1 port map( A1 => n5278, A2 => IF_Regsxreg_file_406_port, B1 
                           => n5360, B2 => IF_Regsxreg_file_662_port, ZN => 
                           n5168);
   U6913 : AOI22_X1 port map( A1 => n5412, A2 => IF_Regsxreg_file_150_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_22_port, ZN => 
                           n5167);
   U6914 : NAND4_X1 port map( A1 => n5170, A2 => n5169, A3 => n5168, A4 => 
                           n5167, ZN => n5171);
   U6915 : AOI211_X1 port map( C1 => n6266, C2 => n5173, A => n5172, B => n5171
                           , ZN => n5174);
   U6916 : AOI21_X1 port map( B1 => n5175, B2 => n5174, A => n5216, ZN => 
                           IF_RegsxN649);
   U6917 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_503_port, B1 
                           => n5399, B2 => IF_Regsxreg_file_343_port, ZN => 
                           n5178);
   U6918 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_855_port, B1 
                           => n5250, B2 => IF_Regsxreg_file_599_port, ZN => 
                           n5177);
   U6919 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_87_port, B1 
                           => n5273, B2 => IF_Regsxreg_file_759_port, ZN => 
                           n5176);
   U6920 : NAND3_X1 port map( A1 => n5178, A2 => n5177, A3 => n5176, ZN => 
                           n5179);
   U6921 : AOI21_X1 port map( B1 => n5383, B2 => IF_Regsxreg_file_919_port, A 
                           => n5179, ZN => n5196);
   U6922 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_951_port, B1 
                           => n5384, B2 => IF_Regsxreg_file_823_port, ZN => 
                           n5183);
   U6923 : AOI22_X1 port map( A1 => n5294, A2 => IF_Regsxreg_file_183_port, B1 
                           => n5390, B2 => IF_Regsxreg_file_311_port, ZN => 
                           n5182);
   U6924 : AOI22_X1 port map( A1 => n5391, A2 => IF_Regsxreg_file_695_port, B1 
                           => n5386, B2 => IF_Regsxreg_file_439_port, ZN => 
                           n5181);
   U6925 : AOI22_X1 port map( A1 => n5385, A2 => IF_Regsxreg_file_567_port, B1 
                           => n5388, B2 => IF_Regsxreg_file_55_port, ZN => 
                           n5180);
   U6926 : NAND4_X1 port map( A1 => n5183, A2 => n5182, A3 => n5181, A4 => 
                           n5180, ZN => n5194);
   U6927 : AOI22_X1 port map( A1 => n5325, A2 => IF_Regsxreg_file_471_port, B1 
                           => n5400, B2 => IF_Regsxreg_file_375_port, ZN => 
                           n5187);
   U6928 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_119_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_247_port, ZN => 
                           n5186);
   U6929 : AOI22_X1 port map( A1 => n5396, A2 => IF_Regsxreg_file_887_port, B1 
                           => n5398, B2 => IF_Regsxreg_file_215_port, ZN => 
                           n5185);
   U6930 : AOI22_X1 port map( A1 => n5352, A2 => IF_Regsxreg_file_983_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_631_port, ZN => 
                           n5184);
   U6931 : NAND4_X1 port map( A1 => n5187, A2 => n5186, A3 => n5185, A4 => 
                           n5184, ZN => n5193);
   U6932 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_727_port, B1 
                           => n5360, B2 => IF_Regsxreg_file_663_port, ZN => 
                           n5191);
   U6933 : AOI22_X1 port map( A1 => n5279, A2 => IF_Regsxreg_file_791_port, B1 
                           => n5414, B2 => IF_Regsxreg_file_407_port, ZN => 
                           n5190);
   U6934 : AOI22_X1 port map( A1 => n5359, A2 => IF_Regsxreg_file_535_port, B1 
                           => n5363, B2 => IF_Regsxreg_file_279_port, ZN => 
                           n5189);
   U6935 : AOI22_X1 port map( A1 => n5412, A2 => IF_Regsxreg_file_151_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_23_port, ZN => 
                           n5188);
   U6936 : NAND4_X1 port map( A1 => n5191, A2 => n5190, A3 => n5189, A4 => 
                           n5188, ZN => n5192);
   U6937 : AOI211_X1 port map( C1 => n6266, C2 => n5194, A => n5193, B => n5192
                           , ZN => n5195);
   U6938 : AOI21_X1 port map( B1 => n5196, B2 => n5195, A => n5216, ZN => 
                           IF_RegsxN650);
   U6939 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_504_port, B1 
                           => n5399, B2 => IF_Regsxreg_file_344_port, ZN => 
                           n5199);
   U6940 : AOI22_X1 port map( A1 => n5352, A2 => IF_Regsxreg_file_984_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_248_port, ZN => 
                           n5198);
   U6941 : AOI22_X1 port map( A1 => n5325, A2 => IF_Regsxreg_file_472_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_216_port, ZN => 
                           n5197);
   U6942 : NAND3_X1 port map( A1 => n5199, A2 => n5198, A3 => n5197, ZN => 
                           n5200);
   U6943 : AOI21_X1 port map( B1 => n5362, B2 => IF_Regsxreg_file_24_port, A =>
                           n5200, ZN => n5218);
   U6944 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_696_port, B1 
                           => n5384, B2 => IF_Regsxreg_file_824_port, ZN => 
                           n5204);
   U6945 : AOI22_X1 port map( A1 => n5294, A2 => IF_Regsxreg_file_184_port, B1 
                           => n5390, B2 => IF_Regsxreg_file_312_port, ZN => 
                           n5203);
   U6946 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_952_port, B1 
                           => n5386, B2 => IF_Regsxreg_file_440_port, ZN => 
                           n5202);
   U6947 : AOI22_X1 port map( A1 => n5345, A2 => IF_Regsxreg_file_568_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_56_port, ZN => 
                           n5201);
   U6948 : NAND4_X1 port map( A1 => n5204, A2 => n5203, A3 => n5202, A4 => 
                           n5201, ZN => n5215);
   U6949 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_728_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_376_port, ZN => 
                           n5208);
   U6950 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_120_port, B1 
                           => n5378, B2 => IF_Regsxreg_file_88_port, ZN => 
                           n5207);
   U6951 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_856_port, B1 
                           => n5397, B2 => IF_Regsxreg_file_600_port, ZN => 
                           n5206);
   U6952 : AOI22_X1 port map( A1 => n5273, A2 => IF_Regsxreg_file_760_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_632_port, ZN => 
                           n5205);
   U6953 : NAND4_X1 port map( A1 => n5208, A2 => n5207, A3 => n5206, A4 => 
                           n5205, ZN => n5214);
   U6954 : AOI22_X1 port map( A1 => n5300, A2 => IF_Regsxreg_file_888_port, B1 
                           => n5363, B2 => IF_Regsxreg_file_280_port, ZN => 
                           n5212);
   U6955 : AOI22_X1 port map( A1 => n5359, A2 => IF_Regsxreg_file_536_port, B1 
                           => n5411, B2 => IF_Regsxreg_file_792_port, ZN => 
                           n5211);
   U6956 : AOI22_X1 port map( A1 => n5278, A2 => IF_Regsxreg_file_408_port, B1 
                           => n5360, B2 => IF_Regsxreg_file_664_port, ZN => 
                           n5210);
   U6957 : AOI22_X1 port map( A1 => n5361, A2 => IF_Regsxreg_file_152_port, B1 
                           => n5383, B2 => IF_Regsxreg_file_920_port, ZN => 
                           n5209);
   U6958 : NAND4_X1 port map( A1 => n5212, A2 => n5211, A3 => n5210, A4 => 
                           n5209, ZN => n5213);
   U6959 : AOI211_X1 port map( C1 => n6266, C2 => n5215, A => n5214, B => n5213
                           , ZN => n5217);
   U6960 : CLKBUF_X1 port map( A => n5216, Z => n5423);
   U6961 : AOI21_X1 port map( B1 => n5218, B2 => n5217, A => n5423, ZN => 
                           IF_RegsxN651);
   U6962 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_505_port, B1 
                           => n5396, B2 => IF_Regsxreg_file_889_port, ZN => 
                           n5221);
   U6963 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_601_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_217_port, ZN => 
                           n5220);
   U6964 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_729_port, B1 
                           => n5399, B2 => IF_Regsxreg_file_345_port, ZN => 
                           n5219);
   U6965 : NAND3_X1 port map( A1 => n5221, A2 => n5220, A3 => n5219, ZN => 
                           n5222);
   U6966 : AOI21_X1 port map( B1 => n5360, B2 => IF_Regsxreg_file_665_port, A 
                           => n5222, ZN => n5239);
   U6967 : AOI22_X1 port map( A1 => n5385, A2 => IF_Regsxreg_file_569_port, B1 
                           => n5386, B2 => IF_Regsxreg_file_441_port, ZN => 
                           n5226);
   U6968 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_185_port, B1 
                           => n5388, B2 => IF_Regsxreg_file_57_port, ZN => 
                           n5225);
   U6969 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_953_port, B1 
                           => n5384, B2 => IF_Regsxreg_file_825_port, ZN => 
                           n5224);
   U6970 : AOI22_X1 port map( A1 => n5391, A2 => IF_Regsxreg_file_697_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_313_port, ZN => 
                           n5223);
   U6971 : NAND4_X1 port map( A1 => n5226, A2 => n5225, A3 => n5224, A4 => 
                           n5223, ZN => n5237);
   U6972 : AOI22_X1 port map( A1 => n5352, A2 => IF_Regsxreg_file_985_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_633_port, ZN => 
                           n5230);
   U6973 : AOI22_X1 port map( A1 => n5299, A2 => IF_Regsxreg_file_249_port, B1 
                           => n5273, B2 => IF_Regsxreg_file_761_port, ZN => 
                           n5229);
   U6974 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_857_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_377_port, ZN => 
                           n5228);
   U6975 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_89_port, B1 
                           => n5325, B2 => IF_Regsxreg_file_473_port, ZN => 
                           n5227);
   U6976 : NAND4_X1 port map( A1 => n5230, A2 => n5229, A3 => n5228, A4 => 
                           n5227, ZN => n5236);
   U6977 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_121_port, B1 
                           => n5412, B2 => IF_Regsxreg_file_153_port, ZN => 
                           n5234);
   U6978 : AOI22_X1 port map( A1 => n5279, A2 => IF_Regsxreg_file_793_port, B1 
                           => n5383, B2 => IF_Regsxreg_file_921_port, ZN => 
                           n5233);
   U6979 : AOI22_X1 port map( A1 => n5359, A2 => IF_Regsxreg_file_537_port, B1 
                           => n5414, B2 => IF_Regsxreg_file_409_port, ZN => 
                           n5232);
   U6980 : AOI22_X1 port map( A1 => n5363, A2 => IF_Regsxreg_file_281_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_25_port, ZN => 
                           n5231);
   U6981 : NAND4_X1 port map( A1 => n5234, A2 => n5233, A3 => n5232, A4 => 
                           n5231, ZN => n5235);
   U6982 : AOI211_X1 port map( C1 => n6266, C2 => n5237, A => n5236, B => n5235
                           , ZN => n5238);
   U6983 : AOI21_X1 port map( B1 => n5239, B2 => n5238, A => n5423, ZN => 
                           IF_RegsxN652);
   U6984 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_506_port, B1 
                           => n5240, B2 => IF_Regsxreg_file_90_port, ZN => 
                           n5243);
   U6985 : AOI22_X1 port map( A1 => n5402, A2 => IF_Regsxreg_file_762_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_378_port, ZN => 
                           n5242);
   U6986 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_858_port, B1 
                           => n5373, B2 => IF_Regsxreg_file_474_port, ZN => 
                           n5241);
   U6987 : NAND3_X1 port map( A1 => n5243, A2 => n5242, A3 => n5241, ZN => 
                           n5244);
   U6988 : AOI21_X1 port map( B1 => n5278, B2 => IF_Regsxreg_file_410_port, A 
                           => n5244, ZN => n5263);
   U6989 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_698_port, B1 
                           => n5385, B2 => IF_Regsxreg_file_570_port, ZN => 
                           n5249);
   U6990 : AOI22_X1 port map( A1 => n5293, A2 => IF_Regsxreg_file_442_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_58_port, ZN => 
                           n5248);
   U6991 : AOI22_X1 port map( A1 => n5384, A2 => IF_Regsxreg_file_826_port, B1 
                           => n5390, B2 => IF_Regsxreg_file_314_port, ZN => 
                           n5247);
   U6992 : AOI22_X1 port map( A1 => n5294, A2 => IF_Regsxreg_file_186_port, B1 
                           => n5245, B2 => IF_Regsxreg_file_954_port, ZN => 
                           n5246);
   U6993 : NAND4_X1 port map( A1 => n5249, A2 => n5248, A3 => n5247, A4 => 
                           n5246, ZN => n5261);
   U6994 : AOI22_X1 port map( A1 => n5352, A2 => IF_Regsxreg_file_986_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_218_port, ZN => 
                           n5254);
   U6995 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_730_port, B1 
                           => n5250, B2 => IF_Regsxreg_file_602_port, ZN => 
                           n5253);
   U6996 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_122_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_250_port, ZN => 
                           n5252);
   U6997 : AOI22_X1 port map( A1 => n5354, A2 => IF_Regsxreg_file_346_port, B1 
                           => n5300, B2 => IF_Regsxreg_file_890_port, ZN => 
                           n5251);
   U6998 : NAND4_X1 port map( A1 => n5254, A2 => n5253, A3 => n5252, A4 => 
                           n5251, ZN => n5260);
   U6999 : AOI22_X1 port map( A1 => n5375, A2 => IF_Regsxreg_file_634_port, B1 
                           => n5383, B2 => IF_Regsxreg_file_922_port, ZN => 
                           n5258);
   U7000 : AOI22_X1 port map( A1 => n5359, A2 => IF_Regsxreg_file_538_port, B1 
                           => n5363, B2 => IF_Regsxreg_file_282_port, ZN => 
                           n5257);
   U7001 : AOI22_X1 port map( A1 => n5362, A2 => IF_Regsxreg_file_26_port, B1 
                           => n5360, B2 => IF_Regsxreg_file_666_port, ZN => 
                           n5256);
   U7002 : AOI22_X1 port map( A1 => n5279, A2 => IF_Regsxreg_file_794_port, B1 
                           => n5412, B2 => IF_Regsxreg_file_154_port, ZN => 
                           n5255);
   U7003 : NAND4_X1 port map( A1 => n5258, A2 => n5257, A3 => n5256, A4 => 
                           n5255, ZN => n5259);
   U7004 : AOI211_X1 port map( C1 => n6266, C2 => n5261, A => n5260, B => n5259
                           , ZN => n5262);
   U7005 : AOI21_X1 port map( B1 => n5263, B2 => n5262, A => n5423, ZN => 
                           IF_RegsxN653);
   U7006 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_507_port, B1 
                           => n5399, B2 => IF_Regsxreg_file_347_port, ZN => 
                           n5267);
   U7007 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_859_port, B1 
                           => n5396, B2 => IF_Regsxreg_file_891_port, ZN => 
                           n5266);
   U7008 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_123_port, B1 
                           => n5264, B2 => IF_Regsxreg_file_987_port, ZN => 
                           n5265);
   U7009 : NAND3_X1 port map( A1 => n5267, A2 => n5266, A3 => n5265, ZN => 
                           n5268);
   U7010 : AOI21_X1 port map( B1 => n5413, B2 => IF_Regsxreg_file_283_port, A 
                           => n5268, ZN => n5288);
   U7011 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_699_port, B1 
                           => n5386, B2 => IF_Regsxreg_file_443_port, ZN => 
                           n5272);
   U7012 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_187_port, B1 
                           => n5385, B2 => IF_Regsxreg_file_571_port, ZN => 
                           n5271);
   U7013 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_955_port, B1 
                           => n5390, B2 => IF_Regsxreg_file_315_port, ZN => 
                           n5270);
   U7014 : AOI22_X1 port map( A1 => n5384, A2 => IF_Regsxreg_file_827_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_59_port, ZN => 
                           n5269);
   U7015 : NAND4_X1 port map( A1 => n5272, A2 => n5271, A3 => n5270, A4 => 
                           n5269, ZN => n5286);
   U7016 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_731_port, B1 
                           => n5273, B2 => IF_Regsxreg_file_763_port, ZN => 
                           n5277);
   U7017 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_603_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_251_port, ZN => 
                           n5276);
   U7018 : AOI22_X1 port map( A1 => n5373, A2 => IF_Regsxreg_file_475_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_635_port, ZN => 
                           n5275);
   U7019 : AOI22_X1 port map( A1 => n5353, A2 => IF_Regsxreg_file_219_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_379_port, ZN => 
                           n5274);
   U7020 : NAND4_X1 port map( A1 => n5277, A2 => n5276, A3 => n5275, A4 => 
                           n5274, ZN => n5285);
   U7021 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_91_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_27_port, ZN => 
                           n5283);
   U7022 : AOI22_X1 port map( A1 => n5278, A2 => IF_Regsxreg_file_411_port, B1 
                           => n5360, B2 => IF_Regsxreg_file_667_port, ZN => 
                           n5282);
   U7023 : AOI22_X1 port map( A1 => n5279, A2 => IF_Regsxreg_file_795_port, B1 
                           => n5412, B2 => IF_Regsxreg_file_155_port, ZN => 
                           n5281);
   U7024 : AOI22_X1 port map( A1 => n5359, A2 => IF_Regsxreg_file_539_port, B1 
                           => n5383, B2 => IF_Regsxreg_file_923_port, ZN => 
                           n5280);
   U7025 : NAND4_X1 port map( A1 => n5283, A2 => n5282, A3 => n5281, A4 => 
                           n5280, ZN => n5284);
   U7026 : AOI211_X1 port map( C1 => n6266, C2 => n5286, A => n5285, B => n5284
                           , ZN => n5287);
   U7027 : AOI21_X1 port map( B1 => n5288, B2 => n5287, A => n5423, ZN => 
                           IF_RegsxN654);
   U7028 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_508_port, B1 
                           => n5401, B2 => IF_Regsxreg_file_732_port, ZN => 
                           n5291);
   U7029 : AOI22_X1 port map( A1 => n5352, A2 => IF_Regsxreg_file_988_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_764_port, ZN => 
                           n5290);
   U7030 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_92_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_380_port, ZN => 
                           n5289);
   U7031 : NAND3_X1 port map( A1 => n5291, A2 => n5290, A3 => n5289, ZN => 
                           n5292);
   U7032 : AOI21_X1 port map( B1 => n5383, B2 => IF_Regsxreg_file_924_port, A 
                           => n5292, ZN => n5313);
   U7033 : AOI22_X1 port map( A1 => n5293, A2 => IF_Regsxreg_file_444_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_60_port, ZN => 
                           n5298);
   U7034 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_700_port, B1 
                           => n5385, B2 => IF_Regsxreg_file_572_port, ZN => 
                           n5297);
   U7035 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_956_port, B1 
                           => n5390, B2 => IF_Regsxreg_file_316_port, ZN => 
                           n5296);
   U7036 : AOI22_X1 port map( A1 => n5294, A2 => IF_Regsxreg_file_188_port, B1 
                           => n5384, B2 => IF_Regsxreg_file_828_port, ZN => 
                           n5295);
   U7037 : NAND4_X1 port map( A1 => n5298, A2 => n5297, A3 => n5296, A4 => 
                           n5295, ZN => n5311);
   U7038 : AOI22_X1 port map( A1 => n5325, A2 => IF_Regsxreg_file_476_port, B1 
                           => n5299, B2 => IF_Regsxreg_file_252_port, ZN => 
                           n5304);
   U7039 : AOI22_X1 port map( A1 => n5300, A2 => IF_Regsxreg_file_892_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_636_port, ZN => 
                           n5303);
   U7040 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_860_port, B1 
                           => n5397, B2 => IF_Regsxreg_file_604_port, ZN => 
                           n5302);
   U7041 : AOI22_X1 port map( A1 => n5354, A2 => IF_Regsxreg_file_348_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_220_port, ZN => 
                           n5301);
   U7042 : NAND4_X1 port map( A1 => n5304, A2 => n5303, A3 => n5302, A4 => 
                           n5301, ZN => n5310);
   U7043 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_124_port, B1 
                           => n5411, B2 => IF_Regsxreg_file_796_port, ZN => 
                           n5308);
   U7044 : AOI22_X1 port map( A1 => n5359, A2 => IF_Regsxreg_file_540_port, B1 
                           => n5360, B2 => IF_Regsxreg_file_668_port, ZN => 
                           n5307);
   U7045 : AOI22_X1 port map( A1 => n5361, A2 => IF_Regsxreg_file_156_port, B1 
                           => n5414, B2 => IF_Regsxreg_file_412_port, ZN => 
                           n5306);
   U7046 : AOI22_X1 port map( A1 => n5363, A2 => IF_Regsxreg_file_284_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_28_port, ZN => 
                           n5305);
   U7047 : NAND4_X1 port map( A1 => n5308, A2 => n5307, A3 => n5306, A4 => 
                           n5305, ZN => n5309);
   U7048 : AOI211_X1 port map( C1 => n6266, C2 => n5311, A => n5310, B => n5309
                           , ZN => n5312);
   U7049 : AOI21_X1 port map( B1 => n5313, B2 => n5312, A => n5423, ZN => 
                           IF_RegsxN655);
   U7050 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_509_port, B1 
                           => n5314, B2 => IF_Regsxreg_file_861_port, ZN => 
                           n5317);
   U7051 : AOI22_X1 port map( A1 => n5377, A2 => IF_Regsxreg_file_253_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_221_port, ZN => 
                           n5316);
   U7052 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_93_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_765_port, ZN => 
                           n5315);
   U7053 : NAND3_X1 port map( A1 => n5317, A2 => n5316, A3 => n5315, ZN => 
                           n5318);
   U7054 : AOI21_X1 port map( B1 => n5411, B2 => IF_Regsxreg_file_797_port, A 
                           => n5318, ZN => n5339);
   U7055 : AOI22_X1 port map( A1 => n5384, A2 => IF_Regsxreg_file_829_port, B1 
                           => n5319, B2 => IF_Regsxreg_file_61_port, ZN => 
                           n5324);
   U7056 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_957_port, B1 
                           => n5386, B2 => IF_Regsxreg_file_445_port, ZN => 
                           n5323);
   U7057 : AOI22_X1 port map( A1 => n5320, A2 => IF_Regsxreg_file_701_port, B1 
                           => n5385, B2 => IF_Regsxreg_file_573_port, ZN => 
                           n5322);
   U7058 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_189_port, B1 
                           => n5390, B2 => IF_Regsxreg_file_317_port, ZN => 
                           n5321);
   U7059 : NAND4_X1 port map( A1 => n5324, A2 => n5323, A3 => n5322, A4 => 
                           n5321, ZN => n5337);
   U7060 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_605_port, B1 
                           => n5399, B2 => IF_Regsxreg_file_349_port, ZN => 
                           n5329);
   U7061 : AOI22_X1 port map( A1 => n5375, A2 => IF_Regsxreg_file_637_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_381_port, ZN => 
                           n5328);
   U7062 : AOI22_X1 port map( A1 => n5396, A2 => IF_Regsxreg_file_893_port, B1 
                           => n5325, B2 => IF_Regsxreg_file_477_port, ZN => 
                           n5327);
   U7063 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_125_port, B1 
                           => n5376, B2 => IF_Regsxreg_file_989_port, ZN => 
                           n5326);
   U7064 : NAND4_X1 port map( A1 => n5329, A2 => n5328, A3 => n5327, A4 => 
                           n5326, ZN => n5336);
   U7065 : AOI22_X1 port map( A1 => n5330, A2 => IF_Regsxreg_file_733_port, B1 
                           => n5362, B2 => IF_Regsxreg_file_29_port, ZN => 
                           n5334);
   U7066 : AOI22_X1 port map( A1 => n5359, A2 => IF_Regsxreg_file_541_port, B1 
                           => n5414, B2 => IF_Regsxreg_file_413_port, ZN => 
                           n5333);
   U7067 : AOI22_X1 port map( A1 => n5361, A2 => IF_Regsxreg_file_157_port, B1 
                           => n5383, B2 => IF_Regsxreg_file_925_port, ZN => 
                           n5332);
   U7068 : AOI22_X1 port map( A1 => n5363, A2 => IF_Regsxreg_file_285_port, B1 
                           => n5360, B2 => IF_Regsxreg_file_669_port, ZN => 
                           n5331);
   U7069 : NAND4_X1 port map( A1 => n5334, A2 => n5333, A3 => n5332, A4 => 
                           n5331, ZN => n5335);
   U7070 : AOI211_X1 port map( C1 => n6266, C2 => n5337, A => n5336, B => n5335
                           , ZN => n5338);
   U7071 : AOI21_X1 port map( B1 => n5339, B2 => n5338, A => n5423, ZN => 
                           IF_RegsxN656);
   U7072 : AOI22_X1 port map( A1 => n5340, A2 => IF_Regsxreg_file_510_port, B1 
                           => n5401, B2 => IF_Regsxreg_file_734_port, ZN => 
                           n5343);
   U7073 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_862_port, B1 
                           => n5396, B2 => IF_Regsxreg_file_894_port, ZN => 
                           n5342);
   U7074 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_126_port, B1 
                           => n5373, B2 => IF_Regsxreg_file_478_port, ZN => 
                           n5341);
   U7075 : NAND3_X1 port map( A1 => n5343, A2 => n5342, A3 => n5341, ZN => 
                           n5344);
   U7076 : AOI21_X1 port map( B1 => n5383, B2 => IF_Regsxreg_file_926_port, A 
                           => n5344, ZN => n5372);
   U7077 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_958_port, B1 
                           => n5384, B2 => IF_Regsxreg_file_830_port, ZN => 
                           n5350);
   U7078 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_190_port, B1 
                           => n5388, B2 => IF_Regsxreg_file_62_port, ZN => 
                           n5349);
   U7079 : AOI22_X1 port map( A1 => n5345, A2 => IF_Regsxreg_file_574_port, B1 
                           => n5386, B2 => IF_Regsxreg_file_446_port, ZN => 
                           n5348);
   U7080 : AOI22_X1 port map( A1 => n5391, A2 => IF_Regsxreg_file_702_port, B1 
                           => n5346, B2 => IF_Regsxreg_file_318_port, ZN => 
                           n5347);
   U7081 : NAND4_X1 port map( A1 => n5350, A2 => n5349, A3 => n5348, A4 => 
                           n5347, ZN => n5370);
   U7082 : AOI22_X1 port map( A1 => n5402, A2 => IF_Regsxreg_file_766_port, B1 
                           => n5351, B2 => IF_Regsxreg_file_382_port, ZN => 
                           n5358);
   U7083 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_94_port, B1 
                           => n5352, B2 => IF_Regsxreg_file_990_port, ZN => 
                           n5357);
   U7084 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_606_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_638_port, ZN => 
                           n5356);
   U7085 : AOI22_X1 port map( A1 => n5354, A2 => IF_Regsxreg_file_350_port, B1 
                           => n5353, B2 => IF_Regsxreg_file_222_port, ZN => 
                           n5355);
   U7086 : NAND4_X1 port map( A1 => n5358, A2 => n5357, A3 => n5356, A4 => 
                           n5355, ZN => n5369);
   U7087 : AOI22_X1 port map( A1 => n5377, A2 => IF_Regsxreg_file_254_port, B1 
                           => n5414, B2 => IF_Regsxreg_file_414_port, ZN => 
                           n5367);
   U7088 : AOI22_X1 port map( A1 => n5359, A2 => IF_Regsxreg_file_542_port, B1 
                           => n5411, B2 => IF_Regsxreg_file_798_port, ZN => 
                           n5366);
   U7089 : AOI22_X1 port map( A1 => n5361, A2 => IF_Regsxreg_file_158_port, B1 
                           => n5360, B2 => IF_Regsxreg_file_670_port, ZN => 
                           n5365);
   U7090 : AOI22_X1 port map( A1 => n5363, A2 => IF_Regsxreg_file_286_port, B1 
                           => n5362, B2 => IF_Regsxreg_file_30_port, ZN => 
                           n5364);
   U7091 : NAND4_X1 port map( A1 => n5367, A2 => n5366, A3 => n5365, A4 => 
                           n5364, ZN => n5368);
   U7092 : AOI211_X1 port map( C1 => n6266, C2 => n5370, A => n5369, B => n5368
                           , ZN => n5371);
   U7093 : AOI21_X1 port map( B1 => n5372, B2 => n5371, A => n5423, ZN => 
                           IF_RegsxN657);
   U7094 : AOI22_X1 port map( A1 => n5374, A2 => IF_Regsxreg_file_511_port, B1 
                           => n5373, B2 => IF_Regsxreg_file_479_port, ZN => 
                           n5381);
   U7095 : AOI22_X1 port map( A1 => n5376, A2 => IF_Regsxreg_file_991_port, B1 
                           => n5375, B2 => IF_Regsxreg_file_639_port, ZN => 
                           n5380);
   U7096 : AOI22_X1 port map( A1 => n5378, A2 => IF_Regsxreg_file_95_port, B1 
                           => n5377, B2 => IF_Regsxreg_file_255_port, ZN => 
                           n5379);
   U7097 : NAND3_X1 port map( A1 => n5381, A2 => n5380, A3 => n5379, ZN => 
                           n5382);
   U7098 : AOI21_X1 port map( B1 => n5383, B2 => IF_Regsxreg_file_927_port, A 
                           => n5382, ZN => n5425);
   U7099 : AOI22_X1 port map( A1 => n5385, A2 => IF_Regsxreg_file_575_port, B1 
                           => n5384, B2 => IF_Regsxreg_file_831_port, ZN => 
                           n5395);
   U7100 : AOI22_X1 port map( A1 => n5387, A2 => IF_Regsxreg_file_191_port, B1 
                           => n5386, B2 => IF_Regsxreg_file_447_port, ZN => 
                           n5394);
   U7101 : AOI22_X1 port map( A1 => n5389, A2 => IF_Regsxreg_file_959_port, B1 
                           => n5388, B2 => IF_Regsxreg_file_63_port, ZN => 
                           n5393);
   U7102 : AOI22_X1 port map( A1 => n5391, A2 => IF_Regsxreg_file_703_port, B1 
                           => n5390, B2 => IF_Regsxreg_file_319_port, ZN => 
                           n5392);
   U7103 : NAND4_X1 port map( A1 => n5395, A2 => n5394, A3 => n5393, A4 => 
                           n5392, ZN => n5422);
   U7104 : AOI22_X1 port map( A1 => n5397, A2 => IF_Regsxreg_file_607_port, B1 
                           => n5396, B2 => IF_Regsxreg_file_895_port, ZN => 
                           n5407);
   U7105 : AOI22_X1 port map( A1 => n5399, A2 => IF_Regsxreg_file_351_port, B1 
                           => n5398, B2 => IF_Regsxreg_file_223_port, ZN => 
                           n5406);
   U7106 : AOI22_X1 port map( A1 => n5401, A2 => IF_Regsxreg_file_735_port, B1 
                           => n5400, B2 => IF_Regsxreg_file_383_port, ZN => 
                           n5405);
   U7107 : AOI22_X1 port map( A1 => n5403, A2 => IF_Regsxreg_file_127_port, B1 
                           => n5402, B2 => IF_Regsxreg_file_767_port, ZN => 
                           n5404);
   U7108 : NAND4_X1 port map( A1 => n5407, A2 => n5406, A3 => n5405, A4 => 
                           n5404, ZN => n5421);
   U7109 : AOI22_X1 port map( A1 => n5409, A2 => IF_Regsxreg_file_863_port, B1 
                           => n5408, B2 => IF_Regsxreg_file_31_port, ZN => 
                           n5419);
   U7110 : AOI22_X1 port map( A1 => n5411, A2 => IF_Regsxreg_file_799_port, B1 
                           => n5410, B2 => IF_Regsxreg_file_671_port, ZN => 
                           n5418);
   U7111 : AOI22_X1 port map( A1 => n5413, A2 => IF_Regsxreg_file_287_port, B1 
                           => n5412, B2 => IF_Regsxreg_file_159_port, ZN => 
                           n5417);
   U7112 : AOI22_X1 port map( A1 => n5415, A2 => IF_Regsxreg_file_543_port, B1 
                           => n5414, B2 => IF_Regsxreg_file_415_port, ZN => 
                           n5416);
   U7113 : NAND4_X1 port map( A1 => n5419, A2 => n5418, A3 => n5417, A4 => 
                           n5416, ZN => n5420);
   U7114 : AOI211_X1 port map( C1 => n6266, C2 => n5422, A => n5421, B => n5420
                           , ZN => n5424);
   U7115 : AOI21_X1 port map( B1 => n5425, B2 => n5424, A => n5423, ZN => 
                           IF_RegsxN658);
   U7116 : CLKBUF_X1 port map( A => n6267, Z => n5626);
   U7117 : NOR2_X1 port map( A1 => CtlToRegs_port_src1_3_port, A2 => 
                           CtlToRegs_port_src1_2_port, ZN => n5436);
   U7118 : NAND3_X1 port map( A1 => CtlToRegs_port_src1_4_port, A2 => 
                           CtlToRegs_port_src1_1_port, A3 => n5436, ZN => n5431
                           );
   U7119 : NOR2_X1 port map( A1 => n5626, A2 => n5431, ZN => n6079);
   U7120 : CLKBUF_X1 port map( A => n6079, Z => n6163);
   U7121 : NAND2_X1 port map( A1 => n5626, A2 => n6194, ZN => n5442);
   U7122 : NOR3_X1 port map( A1 => CtlToRegs_port_src1_3_port, A2 => 
                           CtlToRegs_port_src1_2_port, A3 => n5442, ZN => n6015
                           );
   U7123 : CLKBUF_X1 port map( A => n6015, Z => n6126);
   U7124 : NAND3_X1 port map( A1 => CtlToRegs_port_src1_2_port, A2 => n6205, A3
                           => n6256, ZN => n5430);
   U7125 : NAND2_X1 port map( A1 => CtlToRegs_port_src1_0_port, A2 => n6194, ZN
                           => n5447);
   U7126 : NOR2_X1 port map( A1 => n5430, A2 => n5447, ZN => n6148);
   U7127 : AOI22_X1 port map( A1 => IF_Regsxreg_file_480_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_832_port, B2 => n6148, ZN => 
                           n5428);
   U7128 : NAND3_X1 port map( A1 => CtlToRegs_port_src1_3_port, A2 => n6205, A3
                           => n6258, ZN => n5439);
   U7129 : NOR2_X1 port map( A1 => n5439, A2 => n5447, ZN => n6109);
   U7130 : CLKBUF_X1 port map( A => n6109, Z => n6127);
   U7131 : NOR2_X1 port map( A1 => n5442, A2 => n5430, ZN => n6107);
   U7132 : AOI22_X1 port map( A1 => IF_Regsxreg_file_704_port, A2 => n6127, B1 
                           => IF_Regsxreg_file_864_port, B2 => n6107, ZN => 
                           n5427);
   U7133 : NOR4_X1 port map( A1 => CtlToRegs_port_src1_4_port, A2 => 
                           CtlToRegs_port_src1_3_port, A3 => 
                           CtlToRegs_port_src1_2_port, A4 => n5447, ZN => n6090
                           );
   U7134 : CLKBUF_X1 port map( A => n6090, Z => n6154);
   U7135 : NAND3_X1 port map( A1 => CtlToRegs_port_src1_3_port, A2 => 
                           CtlToRegs_port_src1_4_port, A3 => n6258, ZN => n5440
                           );
   U7136 : NOR2_X1 port map( A1 => n5442, A2 => n5440, ZN => n6046);
   U7137 : CLKBUF_X1 port map( A => n6046, Z => n6152);
   U7138 : AOI22_X1 port map( A1 => IF_Regsxreg_file_960_port, A2 => n6154, B1 
                           => IF_Regsxreg_file_224_port, B2 => n6152, ZN => 
                           n5426);
   U7139 : NAND3_X1 port map( A1 => n5428, A2 => n5427, A3 => n5426, ZN => 
                           n5429);
   U7140 : AOI21_X1 port map( B1 => IF_Regsxreg_file_384_port, B2 => n6163, A 
                           => n5429, ZN => n5459);
   U7141 : NOR2_X1 port map( A1 => n6194, A2 => n5430, ZN => n6067);
   U7142 : CLKBUF_X1 port map( A => n6067, Z => n6137);
   U7143 : INV_X1 port map( A => n5431, ZN => n6136);
   U7144 : AOI22_X1 port map( A1 => IF_Regsxreg_file_800_port, A2 => n6137, B1 
                           => IF_Regsxreg_file_416_port, B2 => n6136, ZN => 
                           n5435);
   U7145 : NOR2_X1 port map( A1 => n6194, A2 => n5439, ZN => n6041);
   U7146 : CLKBUF_X1 port map( A => n6041, Z => n6140);
   U7147 : NAND3_X1 port map( A1 => CtlToRegs_port_src1_3_port, A2 => 
                           CtlToRegs_port_src1_2_port, A3 => n6205, ZN => n5438
                           );
   U7148 : NOR2_X1 port map( A1 => n6194, A2 => n5438, ZN => n6096);
   U7149 : AOI22_X1 port map( A1 => IF_Regsxreg_file_672_port, A2 => n6140, B1 
                           => IF_Regsxreg_file_544_port, B2 => n6096, ZN => 
                           n5434);
   U7150 : NAND3_X1 port map( A1 => CtlToRegs_port_src1_4_port, A2 => 
                           CtlToRegs_port_src1_2_port, A3 => n6256, ZN => n5441
                           );
   U7151 : NOR2_X1 port map( A1 => n6194, A2 => n5441, ZN => n6141);
   U7152 : NAND3_X1 port map( A1 => CtlToRegs_port_src1_4_port, A2 => 
                           CtlToRegs_port_src1_3_port, A3 => 
                           CtlToRegs_port_src1_2_port, ZN => n5448);
   U7153 : NOR2_X1 port map( A1 => n6194, A2 => n5448, ZN => n6142);
   U7154 : AOI22_X1 port map( A1 => IF_Regsxreg_file_288_port, A2 => n6141, B1 
                           => IF_Regsxreg_file_32_port, B2 => n6142, ZN => 
                           n5433);
   U7155 : NOR2_X1 port map( A1 => n6194, A2 => n5440, ZN => n6097);
   U7156 : NOR4_X1 port map( A1 => CtlToRegs_port_src1_4_port, A2 => 
                           CtlToRegs_port_src1_3_port, A3 => 
                           CtlToRegs_port_src1_2_port, A4 => n6194, ZN => n5449
                           );
   U7157 : CLKBUF_X1 port map( A => n5449, Z => n6138);
   U7158 : AOI22_X1 port map( A1 => IF_Regsxreg_file_160_port, A2 => n6097, B1 
                           => IF_Regsxreg_file_928_port, B2 => n6138, ZN => 
                           n5432);
   U7159 : NAND4_X1 port map( A1 => n5435, A2 => n5434, A3 => n5433, A4 => 
                           n5432, ZN => n5456);
   U7160 : NAND2_X1 port map( A1 => CtlToRegs_port_src1_4_port, A2 => n5436, ZN
                           => n5437);
   U7161 : NOR2_X1 port map( A1 => n5437, A2 => n5447, ZN => n6155);
   U7162 : CLKBUF_X1 port map( A => n6155, Z => n6106);
   U7163 : NOR2_X1 port map( A1 => n5442, A2 => n5438, ZN => n6005);
   U7164 : CLKBUF_X1 port map( A => n6005, Z => n6153);
   U7165 : AOI22_X1 port map( A1 => IF_Regsxreg_file_448_port, A2 => n6106, B1 
                           => IF_Regsxreg_file_608_port, B2 => n6153, ZN => 
                           n5446);
   U7166 : NOR2_X1 port map( A1 => n5442, A2 => n5448, ZN => n6114);
   U7167 : CLKBUF_X1 port map( A => n6114, Z => n6129);
   U7168 : NOR2_X1 port map( A1 => n5441, A2 => n5447, ZN => n6104);
   U7169 : AOI22_X1 port map( A1 => IF_Regsxreg_file_96_port, A2 => n6129, B1 
                           => IF_Regsxreg_file_320_port, B2 => n6104, ZN => 
                           n5445);
   U7170 : NOR2_X1 port map( A1 => n5438, A2 => n5447, ZN => n6074);
   U7171 : CLKBUF_X1 port map( A => n6074, Z => n6151);
   U7172 : NOR2_X1 port map( A1 => n5442, A2 => n5439, ZN => n6150);
   U7173 : CLKBUF_X1 port map( A => n6150, Z => n6091);
   U7174 : AOI22_X1 port map( A1 => IF_Regsxreg_file_576_port, A2 => n6151, B1 
                           => IF_Regsxreg_file_736_port, B2 => n6091, ZN => 
                           n5444);
   U7175 : NOR2_X1 port map( A1 => n5440, A2 => n5447, ZN => n5826);
   U7176 : NOR2_X1 port map( A1 => n5442, A2 => n5441, ZN => n6108);
   U7177 : CLKBUF_X1 port map( A => n6108, Z => n6130);
   U7178 : AOI22_X1 port map( A1 => IF_Regsxreg_file_192_port, A2 => n5826, B1 
                           => IF_Regsxreg_file_352_port, B2 => n6130, ZN => 
                           n5443);
   U7179 : NAND4_X1 port map( A1 => n5446, A2 => n5445, A3 => n5444, A4 => 
                           n5443, ZN => n5455);
   U7180 : NOR2_X1 port map( A1 => n5448, A2 => n5447, ZN => n6062);
   U7181 : CLKBUF_X1 port map( A => n6062, Z => n6149);
   U7182 : CLKBUF_X1 port map( A => n6141, Z => n6098);
   U7183 : AND2_X1 port map( A1 => CtlToRegs_port_src1_0_port, A2 => n6098, ZN 
                           => n6160);
   U7184 : AOI22_X1 port map( A1 => IF_Regsxreg_file_64_port, A2 => n6149, B1 
                           => IF_Regsxreg_file_256_port, B2 => n6160, ZN => 
                           n5453);
   U7185 : CLKBUF_X1 port map( A => n6142, Z => n6068);
   U7186 : AND2_X1 port map( A1 => CtlToRegs_port_src1_0_port, A2 => n6068, ZN 
                           => n6165);
   U7187 : AND2_X1 port map( A1 => CtlToRegs_port_src1_0_port, A2 => n6140, ZN 
                           => n6166);
   U7188 : AOI22_X1 port map( A1 => IF_Regsxreg_file_0_port, A2 => n6165, B1 =>
                           IF_Regsxreg_file_640_port, B2 => n6166, ZN => n5452)
                           ;
   U7189 : CLKBUF_X1 port map( A => n6097, Z => n6139);
   U7190 : AND2_X1 port map( A1 => CtlToRegs_port_src1_0_port, A2 => n6139, ZN 
                           => n6115);
   U7191 : CLKBUF_X1 port map( A => n5449, Z => n5886);
   U7192 : AND2_X1 port map( A1 => CtlToRegs_port_src1_0_port, A2 => n5886, ZN 
                           => n6167);
   U7193 : AOI22_X1 port map( A1 => IF_Regsxreg_file_128_port, A2 => n6115, B1 
                           => IF_Regsxreg_file_896_port, B2 => n6167, ZN => 
                           n5451);
   U7194 : CLKBUF_X1 port map( A => n6096, Z => n6143);
   U7195 : AND2_X1 port map( A1 => CtlToRegs_port_src1_0_port, A2 => n6143, ZN 
                           => n6080);
   U7196 : AND2_X1 port map( A1 => CtlToRegs_port_src1_0_port, A2 => n6137, ZN 
                           => n6135);
   U7197 : CLKBUF_X1 port map( A => n6135, Z => n6051);
   U7198 : AOI22_X1 port map( A1 => IF_Regsxreg_file_512_port, A2 => n6080, B1 
                           => IF_Regsxreg_file_768_port, B2 => n6051, ZN => 
                           n5450);
   U7199 : NAND4_X1 port map( A1 => n5453, A2 => n5452, A3 => n5451, A4 => 
                           n5450, ZN => n5454);
   U7200 : AOI211_X1 port map( C1 => n5626, C2 => n5456, A => n5455, B => n5454
                           , ZN => n5458);
   U7201 : CLKBUF_X1 port map( A => n6015, Z => n5926);
   U7202 : AOI21_X1 port map( B1 => n6205, B2 => n5926, A => rst, ZN => n5457);
   U7203 : INV_X1 port map( A => n5457, ZN => n5968);
   U7204 : AOI21_X1 port map( B1 => n5459, B2 => n5458, A => n5968, ZN => 
                           IF_RegsxN595);
   U7205 : CLKBUF_X1 port map( A => n6165, Z => n6052);
   U7206 : AOI22_X1 port map( A1 => IF_Regsxreg_file_481_port, A2 => n5926, B1 
                           => IF_Regsxreg_file_865_port, B2 => n6107, ZN => 
                           n5462);
   U7207 : CLKBUF_X1 port map( A => n5826, Z => n6125);
   U7208 : AOI22_X1 port map( A1 => IF_Regsxreg_file_737_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_193_port, B2 => n6125, ZN => 
                           n5461);
   U7209 : CLKBUF_X1 port map( A => n6104, Z => n6161);
   U7210 : AOI22_X1 port map( A1 => IF_Regsxreg_file_321_port, A2 => n6161, B1 
                           => IF_Regsxreg_file_65_port, B2 => n6062, ZN => 
                           n5460);
   U7211 : NAND3_X1 port map( A1 => n5462, A2 => n5461, A3 => n5460, ZN => 
                           n5463);
   U7212 : AOI21_X1 port map( B1 => IF_Regsxreg_file_1_port, B2 => n6052, A => 
                           n5463, ZN => n5480);
   U7213 : AOI22_X1 port map( A1 => IF_Regsxreg_file_673_port, A2 => n6140, B1 
                           => IF_Regsxreg_file_545_port, B2 => n6143, ZN => 
                           n5467);
   U7214 : AOI22_X1 port map( A1 => IF_Regsxreg_file_289_port, A2 => n6098, B1 
                           => IF_Regsxreg_file_801_port, B2 => n6137, ZN => 
                           n5466);
   U7215 : AOI22_X1 port map( A1 => IF_Regsxreg_file_929_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_417_port, B2 => n6136, ZN => 
                           n5465);
   U7216 : AOI22_X1 port map( A1 => IF_Regsxreg_file_161_port, A2 => n6139, B1 
                           => IF_Regsxreg_file_33_port, B2 => n6068, ZN => 
                           n5464);
   U7217 : NAND4_X1 port map( A1 => n5467, A2 => n5466, A3 => n5465, A4 => 
                           n5464, ZN => n5478);
   U7218 : AOI22_X1 port map( A1 => IF_Regsxreg_file_577_port, A2 => n6151, B1 
                           => IF_Regsxreg_file_705_port, B2 => n6127, ZN => 
                           n5471);
   U7219 : AOI22_X1 port map( A1 => IF_Regsxreg_file_225_port, A2 => n6152, B1 
                           => IF_Regsxreg_file_961_port, B2 => n6154, ZN => 
                           n5470);
   U7220 : AOI22_X1 port map( A1 => IF_Regsxreg_file_353_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_97_port, B2 => n6129, ZN => 
                           n5469);
   U7221 : AOI22_X1 port map( A1 => IF_Regsxreg_file_449_port, A2 => n6155, B1 
                           => IF_Regsxreg_file_609_port, B2 => n6005, ZN => 
                           n5468);
   U7222 : NAND4_X1 port map( A1 => n5471, A2 => n5470, A3 => n5469, A4 => 
                           n5468, ZN => n5477);
   U7223 : CLKBUF_X1 port map( A => n6148, Z => n6105);
   U7224 : AOI22_X1 port map( A1 => IF_Regsxreg_file_833_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_769_port, B2 => n6051, ZN => 
                           n5475);
   U7225 : CLKBUF_X1 port map( A => n6115, Z => n6164);
   U7226 : AOI22_X1 port map( A1 => IF_Regsxreg_file_641_port, A2 => n6166, B1 
                           => IF_Regsxreg_file_129_port, B2 => n6164, ZN => 
                           n5474);
   U7227 : AOI22_X1 port map( A1 => IF_Regsxreg_file_897_port, A2 => n6167, B1 
                           => IF_Regsxreg_file_257_port, B2 => n6160, ZN => 
                           n5473);
   U7228 : CLKBUF_X1 port map( A => n6080, Z => n6162);
   U7229 : AOI22_X1 port map( A1 => IF_Regsxreg_file_385_port, A2 => n6079, B1 
                           => IF_Regsxreg_file_513_port, B2 => n6162, ZN => 
                           n5472);
   U7230 : NAND4_X1 port map( A1 => n5475, A2 => n5474, A3 => n5473, A4 => 
                           n5472, ZN => n5476);
   U7231 : AOI211_X1 port map( C1 => n5626, C2 => n5478, A => n5477, B => n5476
                           , ZN => n5479);
   U7232 : AOI21_X1 port map( B1 => n5480, B2 => n5479, A => n5968, ZN => 
                           IF_RegsxN596);
   U7233 : CLKBUF_X1 port map( A => n6160, Z => n5952);
   U7234 : AOI22_X1 port map( A1 => IF_Regsxreg_file_482_port, A2 => n5926, B1 
                           => IF_Regsxreg_file_578_port, B2 => n6074, ZN => 
                           n5483);
   U7235 : AOI22_X1 port map( A1 => IF_Regsxreg_file_354_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_98_port, B2 => n6114, ZN => 
                           n5482);
   U7236 : AOI22_X1 port map( A1 => IF_Regsxreg_file_962_port, A2 => n6154, B1 
                           => IF_Regsxreg_file_706_port, B2 => n6109, ZN => 
                           n5481);
   U7237 : NAND3_X1 port map( A1 => n5483, A2 => n5482, A3 => n5481, ZN => 
                           n5484);
   U7238 : AOI21_X1 port map( B1 => IF_Regsxreg_file_258_port, B2 => n5952, A 
                           => n5484, ZN => n5501);
   U7239 : AOI22_X1 port map( A1 => IF_Regsxreg_file_34_port, A2 => n6068, B1 
                           => IF_Regsxreg_file_802_port, B2 => n6137, ZN => 
                           n5488);
   U7240 : AOI22_X1 port map( A1 => IF_Regsxreg_file_674_port, A2 => n6140, B1 
                           => IF_Regsxreg_file_162_port, B2 => n6139, ZN => 
                           n5487);
   U7241 : AOI22_X1 port map( A1 => IF_Regsxreg_file_930_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_290_port, B2 => n6098, ZN => 
                           n5486);
   U7242 : AOI22_X1 port map( A1 => IF_Regsxreg_file_546_port, A2 => n6143, B1 
                           => IF_Regsxreg_file_418_port, B2 => n6136, ZN => 
                           n5485);
   U7243 : NAND4_X1 port map( A1 => n5488, A2 => n5487, A3 => n5486, A4 => 
                           n5485, ZN => n5499);
   U7244 : AOI22_X1 port map( A1 => IF_Regsxreg_file_322_port, A2 => n6161, B1 
                           => IF_Regsxreg_file_866_port, B2 => n6107, ZN => 
                           n5492);
   U7245 : AOI22_X1 port map( A1 => IF_Regsxreg_file_450_port, A2 => n6106, B1 
                           => IF_Regsxreg_file_738_port, B2 => n6150, ZN => 
                           n5491);
   U7246 : AOI22_X1 port map( A1 => IF_Regsxreg_file_66_port, A2 => n6149, B1 
                           => IF_Regsxreg_file_194_port, B2 => n6125, ZN => 
                           n5490);
   U7247 : AOI22_X1 port map( A1 => IF_Regsxreg_file_834_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_226_port, B2 => n6152, ZN => 
                           n5489);
   U7248 : NAND4_X1 port map( A1 => n5492, A2 => n5491, A3 => n5490, A4 => 
                           n5489, ZN => n5498);
   U7249 : AOI22_X1 port map( A1 => IF_Regsxreg_file_610_port, A2 => n6153, B1 
                           => IF_Regsxreg_file_130_port, B2 => n6115, ZN => 
                           n5496);
   U7250 : AOI22_X1 port map( A1 => IF_Regsxreg_file_2_port, A2 => n6165, B1 =>
                           IF_Regsxreg_file_514_port, B2 => n6080, ZN => n5495)
                           ;
   U7251 : AOI22_X1 port map( A1 => IF_Regsxreg_file_386_port, A2 => n6163, B1 
                           => IF_Regsxreg_file_770_port, B2 => n6135, ZN => 
                           n5494);
   U7252 : AOI22_X1 port map( A1 => IF_Regsxreg_file_898_port, A2 => n6167, B1 
                           => IF_Regsxreg_file_642_port, B2 => n6166, ZN => 
                           n5493);
   U7253 : NAND4_X1 port map( A1 => n5496, A2 => n5495, A3 => n5494, A4 => 
                           n5493, ZN => n5497);
   U7254 : AOI211_X1 port map( C1 => n5626, C2 => n5499, A => n5498, B => n5497
                           , ZN => n5500);
   U7255 : AOI21_X1 port map( B1 => n5501, B2 => n5500, A => n5968, ZN => 
                           IF_RegsxN597);
   U7256 : AOI22_X1 port map( A1 => IF_Regsxreg_file_483_port, A2 => n6015, B1 
                           => IF_Regsxreg_file_867_port, B2 => n6107, ZN => 
                           n5504);
   U7257 : AOI22_X1 port map( A1 => IF_Regsxreg_file_835_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_195_port, B2 => n5826, ZN => 
                           n5503);
   U7258 : AOI22_X1 port map( A1 => IF_Regsxreg_file_323_port, A2 => n6161, B1 
                           => IF_Regsxreg_file_67_port, B2 => n6062, ZN => 
                           n5502);
   U7259 : NAND3_X1 port map( A1 => n5504, A2 => n5503, A3 => n5502, ZN => 
                           n5505);
   U7260 : AOI21_X1 port map( B1 => IF_Regsxreg_file_515_port, B2 => n6162, A 
                           => n5505, ZN => n5522);
   U7261 : AOI22_X1 port map( A1 => IF_Regsxreg_file_803_port, A2 => n6137, B1 
                           => IF_Regsxreg_file_163_port, B2 => n6139, ZN => 
                           n5509);
   U7262 : AOI22_X1 port map( A1 => IF_Regsxreg_file_675_port, A2 => n6140, B1 
                           => IF_Regsxreg_file_931_port, B2 => n5886, ZN => 
                           n5508);
   U7263 : CLKBUF_X1 port map( A => n6136, Z => n6099);
   U7264 : AOI22_X1 port map( A1 => IF_Regsxreg_file_419_port, A2 => n6099, B1 
                           => IF_Regsxreg_file_547_port, B2 => n6143, ZN => 
                           n5507);
   U7265 : AOI22_X1 port map( A1 => IF_Regsxreg_file_291_port, A2 => n6098, B1 
                           => IF_Regsxreg_file_35_port, B2 => n6068, ZN => 
                           n5506);
   U7266 : NAND4_X1 port map( A1 => n5509, A2 => n5508, A3 => n5507, A4 => 
                           n5506, ZN => n5520);
   U7267 : AOI22_X1 port map( A1 => IF_Regsxreg_file_611_port, A2 => n6153, B1 
                           => IF_Regsxreg_file_963_port, B2 => n6154, ZN => 
                           n5513);
   U7268 : AOI22_X1 port map( A1 => IF_Regsxreg_file_451_port, A2 => n6106, B1 
                           => IF_Regsxreg_file_707_port, B2 => n6109, ZN => 
                           n5512);
   U7269 : AOI22_X1 port map( A1 => IF_Regsxreg_file_739_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_355_port, B2 => n6108, ZN => 
                           n5511);
   U7270 : AOI22_X1 port map( A1 => IF_Regsxreg_file_579_port, A2 => n6151, B1 
                           => IF_Regsxreg_file_227_port, B2 => n6152, ZN => 
                           n5510);
   U7271 : NAND4_X1 port map( A1 => n5513, A2 => n5512, A3 => n5511, A4 => 
                           n5510, ZN => n5519);
   U7272 : AOI22_X1 port map( A1 => IF_Regsxreg_file_99_port, A2 => n6129, B1 
                           => IF_Regsxreg_file_643_port, B2 => n6166, ZN => 
                           n5517);
   U7273 : AOI22_X1 port map( A1 => IF_Regsxreg_file_259_port, A2 => n6160, B1 
                           => IF_Regsxreg_file_3_port, B2 => n6052, ZN => n5516
                           );
   U7274 : AOI22_X1 port map( A1 => IF_Regsxreg_file_387_port, A2 => n6163, B1 
                           => IF_Regsxreg_file_771_port, B2 => n6135, ZN => 
                           n5515);
   U7275 : AOI22_X1 port map( A1 => IF_Regsxreg_file_899_port, A2 => n6167, B1 
                           => IF_Regsxreg_file_131_port, B2 => n6115, ZN => 
                           n5514);
   U7276 : NAND4_X1 port map( A1 => n5517, A2 => n5516, A3 => n5515, A4 => 
                           n5514, ZN => n5518);
   U7277 : AOI211_X1 port map( C1 => n5626, C2 => n5520, A => n5519, B => n5518
                           , ZN => n5521);
   U7278 : AOI21_X1 port map( B1 => n5522, B2 => n5521, A => n5968, ZN => 
                           IF_RegsxN598);
   U7279 : AOI22_X1 port map( A1 => IF_Regsxreg_file_484_port, A2 => n5926, B1 
                           => IF_Regsxreg_file_196_port, B2 => n5826, ZN => 
                           n5525);
   U7280 : AOI22_X1 port map( A1 => IF_Regsxreg_file_580_port, A2 => n6151, B1 
                           => IF_Regsxreg_file_324_port, B2 => n6104, ZN => 
                           n5524);
   U7281 : AOI22_X1 port map( A1 => IF_Regsxreg_file_68_port, A2 => n6149, B1 
                           => IF_Regsxreg_file_708_port, B2 => n6109, ZN => 
                           n5523);
   U7282 : NAND3_X1 port map( A1 => n5525, A2 => n5524, A3 => n5523, ZN => 
                           n5526);
   U7283 : AOI21_X1 port map( B1 => IF_Regsxreg_file_388_port, B2 => n6163, A 
                           => n5526, ZN => n5543);
   U7284 : AOI22_X1 port map( A1 => IF_Regsxreg_file_164_port, A2 => n6139, B1 
                           => IF_Regsxreg_file_420_port, B2 => n6136, ZN => 
                           n5530);
   U7285 : AOI22_X1 port map( A1 => IF_Regsxreg_file_36_port, A2 => n6068, B1 
                           => IF_Regsxreg_file_292_port, B2 => n6141, ZN => 
                           n5529);
   U7286 : AOI22_X1 port map( A1 => IF_Regsxreg_file_804_port, A2 => n6137, B1 
                           => IF_Regsxreg_file_676_port, B2 => n6140, ZN => 
                           n5528);
   U7287 : AOI22_X1 port map( A1 => IF_Regsxreg_file_932_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_548_port, B2 => n6143, ZN => 
                           n5527);
   U7288 : NAND4_X1 port map( A1 => n5530, A2 => n5529, A3 => n5528, A4 => 
                           n5527, ZN => n5541);
   U7289 : AOI22_X1 port map( A1 => IF_Regsxreg_file_356_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_740_port, B2 => n6150, ZN => 
                           n5534);
   U7290 : AOI22_X1 port map( A1 => IF_Regsxreg_file_964_port, A2 => n6154, B1 
                           => IF_Regsxreg_file_100_port, B2 => n6129, ZN => 
                           n5533);
   U7291 : AOI22_X1 port map( A1 => IF_Regsxreg_file_228_port, A2 => n6152, B1 
                           => IF_Regsxreg_file_612_port, B2 => n6005, ZN => 
                           n5532);
   U7292 : AOI22_X1 port map( A1 => IF_Regsxreg_file_452_port, A2 => n6155, B1 
                           => IF_Regsxreg_file_868_port, B2 => n6107, ZN => 
                           n5531);
   U7293 : NAND4_X1 port map( A1 => n5534, A2 => n5533, A3 => n5532, A4 => 
                           n5531, ZN => n5540);
   U7294 : AOI22_X1 port map( A1 => IF_Regsxreg_file_836_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_132_port, B2 => n6115, ZN => 
                           n5538);
   U7295 : AOI22_X1 port map( A1 => IF_Regsxreg_file_260_port, A2 => n6160, B1 
                           => IF_Regsxreg_file_516_port, B2 => n6080, ZN => 
                           n5537);
   U7296 : AOI22_X1 port map( A1 => IF_Regsxreg_file_900_port, A2 => n6167, B1 
                           => IF_Regsxreg_file_772_port, B2 => n6135, ZN => 
                           n5536);
   U7297 : AOI22_X1 port map( A1 => IF_Regsxreg_file_644_port, A2 => n6166, B1 
                           => IF_Regsxreg_file_4_port, B2 => n6165, ZN => n5535
                           );
   U7298 : NAND4_X1 port map( A1 => n5538, A2 => n5537, A3 => n5536, A4 => 
                           n5535, ZN => n5539);
   U7299 : AOI211_X1 port map( C1 => n5626, C2 => n5541, A => n5540, B => n5539
                           , ZN => n5542);
   U7300 : AOI21_X1 port map( B1 => n5543, B2 => n5542, A => n5968, ZN => 
                           IF_RegsxN599);
   U7301 : AOI22_X1 port map( A1 => IF_Regsxreg_file_485_port, A2 => n5926, B1 
                           => IF_Regsxreg_file_101_port, B2 => n6129, ZN => 
                           n5546);
   U7302 : AOI22_X1 port map( A1 => IF_Regsxreg_file_69_port, A2 => n6149, B1 
                           => IF_Regsxreg_file_197_port, B2 => n5826, ZN => 
                           n5545);
   U7303 : AOI22_X1 port map( A1 => IF_Regsxreg_file_581_port, A2 => n6151, B1 
                           => IF_Regsxreg_file_453_port, B2 => n6106, ZN => 
                           n5544);
   U7304 : NAND3_X1 port map( A1 => n5546, A2 => n5545, A3 => n5544, ZN => 
                           n5547);
   U7305 : AOI21_X1 port map( B1 => IF_Regsxreg_file_133_port, B2 => n6164, A 
                           => n5547, ZN => n5564);
   U7306 : AOI22_X1 port map( A1 => IF_Regsxreg_file_933_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_165_port, B2 => n6139, ZN => 
                           n5551);
   U7307 : AOI22_X1 port map( A1 => IF_Regsxreg_file_293_port, A2 => n6098, B1 
                           => IF_Regsxreg_file_549_port, B2 => n6143, ZN => 
                           n5550);
   U7308 : AOI22_X1 port map( A1 => IF_Regsxreg_file_37_port, A2 => n6068, B1 
                           => IF_Regsxreg_file_421_port, B2 => n6136, ZN => 
                           n5549);
   U7309 : AOI22_X1 port map( A1 => IF_Regsxreg_file_677_port, A2 => n6041, B1 
                           => IF_Regsxreg_file_805_port, B2 => n6137, ZN => 
                           n5548);
   U7310 : NAND4_X1 port map( A1 => n5551, A2 => n5550, A3 => n5549, A4 => 
                           n5548, ZN => n5562);
   U7311 : AOI22_X1 port map( A1 => IF_Regsxreg_file_325_port, A2 => n6161, B1 
                           => IF_Regsxreg_file_229_port, B2 => n6046, ZN => 
                           n5555);
   U7312 : AOI22_X1 port map( A1 => IF_Regsxreg_file_741_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_357_port, B2 => n6108, ZN => 
                           n5554);
   U7313 : CLKBUF_X1 port map( A => n6107, Z => n6128);
   U7314 : AOI22_X1 port map( A1 => IF_Regsxreg_file_869_port, A2 => n6128, B1 
                           => IF_Regsxreg_file_709_port, B2 => n6127, ZN => 
                           n5553);
   U7315 : AOI22_X1 port map( A1 => IF_Regsxreg_file_965_port, A2 => n6154, B1 
                           => IF_Regsxreg_file_613_port, B2 => n6005, ZN => 
                           n5552);
   U7316 : NAND4_X1 port map( A1 => n5555, A2 => n5554, A3 => n5553, A4 => 
                           n5552, ZN => n5561);
   U7317 : AOI22_X1 port map( A1 => IF_Regsxreg_file_837_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_773_port, B2 => n6135, ZN => 
                           n5559);
   U7318 : AOI22_X1 port map( A1 => IF_Regsxreg_file_261_port, A2 => n6160, B1 
                           => IF_Regsxreg_file_389_port, B2 => n6079, ZN => 
                           n5558);
   U7319 : CLKBUF_X1 port map( A => n6166, Z => n5895);
   U7320 : AOI22_X1 port map( A1 => IF_Regsxreg_file_5_port, A2 => n6165, B1 =>
                           IF_Regsxreg_file_645_port, B2 => n5895, ZN => n5557)
                           ;
   U7321 : AOI22_X1 port map( A1 => IF_Regsxreg_file_517_port, A2 => n6080, B1 
                           => IF_Regsxreg_file_901_port, B2 => n6167, ZN => 
                           n5556);
   U7322 : NAND4_X1 port map( A1 => n5559, A2 => n5558, A3 => n5557, A4 => 
                           n5556, ZN => n5560);
   U7323 : AOI211_X1 port map( C1 => n5626, C2 => n5562, A => n5561, B => n5560
                           , ZN => n5563);
   U7324 : AOI21_X1 port map( B1 => n5564, B2 => n5563, A => n5968, ZN => 
                           IF_RegsxN600);
   U7325 : AOI22_X1 port map( A1 => IF_Regsxreg_file_486_port, A2 => n5926, B1 
                           => IF_Regsxreg_file_358_port, B2 => n6108, ZN => 
                           n5567);
   U7326 : AOI22_X1 port map( A1 => IF_Regsxreg_file_710_port, A2 => n6127, B1 
                           => IF_Regsxreg_file_966_port, B2 => n6154, ZN => 
                           n5566);
   U7327 : AOI22_X1 port map( A1 => IF_Regsxreg_file_742_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_454_port, B2 => n6155, ZN => 
                           n5565);
   U7328 : NAND3_X1 port map( A1 => n5567, A2 => n5566, A3 => n5565, ZN => 
                           n5568);
   U7329 : AOI21_X1 port map( B1 => IF_Regsxreg_file_134_port, B2 => n6164, A 
                           => n5568, ZN => n5585);
   U7330 : AOI22_X1 port map( A1 => IF_Regsxreg_file_806_port, A2 => n6137, B1 
                           => IF_Regsxreg_file_678_port, B2 => n6140, ZN => 
                           n5572);
   U7331 : AOI22_X1 port map( A1 => IF_Regsxreg_file_38_port, A2 => n6068, B1 
                           => IF_Regsxreg_file_934_port, B2 => n5886, ZN => 
                           n5571);
   U7332 : AOI22_X1 port map( A1 => IF_Regsxreg_file_294_port, A2 => n6098, B1 
                           => IF_Regsxreg_file_550_port, B2 => n6143, ZN => 
                           n5570);
   U7333 : AOI22_X1 port map( A1 => IF_Regsxreg_file_166_port, A2 => n6139, B1 
                           => IF_Regsxreg_file_422_port, B2 => n6136, ZN => 
                           n5569);
   U7334 : NAND4_X1 port map( A1 => n5572, A2 => n5571, A3 => n5570, A4 => 
                           n5569, ZN => n5583);
   U7335 : AOI22_X1 port map( A1 => IF_Regsxreg_file_870_port, A2 => n6128, B1 
                           => IF_Regsxreg_file_582_port, B2 => n6151, ZN => 
                           n5576);
   U7336 : AOI22_X1 port map( A1 => IF_Regsxreg_file_70_port, A2 => n6149, B1 
                           => IF_Regsxreg_file_198_port, B2 => n5826, ZN => 
                           n5575);
   U7337 : AOI22_X1 port map( A1 => IF_Regsxreg_file_230_port, A2 => n6046, B1 
                           => IF_Regsxreg_file_326_port, B2 => n6161, ZN => 
                           n5574);
   U7338 : AOI22_X1 port map( A1 => IF_Regsxreg_file_102_port, A2 => n6129, B1 
                           => IF_Regsxreg_file_614_port, B2 => n6005, ZN => 
                           n5573);
   U7339 : NAND4_X1 port map( A1 => n5576, A2 => n5575, A3 => n5574, A4 => 
                           n5573, ZN => n5582);
   U7340 : AOI22_X1 port map( A1 => IF_Regsxreg_file_838_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_518_port, B2 => n6080, ZN => 
                           n5580);
   U7341 : AOI22_X1 port map( A1 => IF_Regsxreg_file_902_port, A2 => n6167, B1 
                           => IF_Regsxreg_file_390_port, B2 => n6079, ZN => 
                           n5579);
   U7342 : AOI22_X1 port map( A1 => IF_Regsxreg_file_262_port, A2 => n6160, B1 
                           => IF_Regsxreg_file_774_port, B2 => n6135, ZN => 
                           n5578);
   U7343 : AOI22_X1 port map( A1 => IF_Regsxreg_file_6_port, A2 => n6165, B1 =>
                           IF_Regsxreg_file_646_port, B2 => n5895, ZN => n5577)
                           ;
   U7344 : NAND4_X1 port map( A1 => n5580, A2 => n5579, A3 => n5578, A4 => 
                           n5577, ZN => n5581);
   U7345 : AOI211_X1 port map( C1 => n5626, C2 => n5583, A => n5582, B => n5581
                           , ZN => n5584);
   U7346 : AOI21_X1 port map( B1 => n5585, B2 => n5584, A => n5968, ZN => 
                           IF_RegsxN601);
   U7347 : AOI22_X1 port map( A1 => IF_Regsxreg_file_487_port, A2 => n6015, B1 
                           => IF_Regsxreg_file_711_port, B2 => n6109, ZN => 
                           n5588);
   U7348 : AOI22_X1 port map( A1 => IF_Regsxreg_file_359_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_71_port, B2 => n6149, ZN => 
                           n5587);
   U7349 : AOI22_X1 port map( A1 => IF_Regsxreg_file_327_port, A2 => n6161, B1 
                           => IF_Regsxreg_file_871_port, B2 => n6128, ZN => 
                           n5586);
   U7350 : NAND3_X1 port map( A1 => n5588, A2 => n5587, A3 => n5586, ZN => 
                           n5589);
   U7351 : AOI21_X1 port map( B1 => IF_Regsxreg_file_391_port, B2 => n6163, A 
                           => n5589, ZN => n5606);
   U7352 : AOI22_X1 port map( A1 => IF_Regsxreg_file_39_port, A2 => n6068, B1 
                           => IF_Regsxreg_file_167_port, B2 => n6139, ZN => 
                           n5593);
   U7353 : AOI22_X1 port map( A1 => IF_Regsxreg_file_551_port, A2 => n6143, B1 
                           => IF_Regsxreg_file_679_port, B2 => n6140, ZN => 
                           n5592);
   U7354 : AOI22_X1 port map( A1 => IF_Regsxreg_file_295_port, A2 => n6098, B1 
                           => IF_Regsxreg_file_423_port, B2 => n6136, ZN => 
                           n5591);
   U7355 : AOI22_X1 port map( A1 => IF_Regsxreg_file_807_port, A2 => n6137, B1 
                           => IF_Regsxreg_file_935_port, B2 => n5886, ZN => 
                           n5590);
   U7356 : NAND4_X1 port map( A1 => n5593, A2 => n5592, A3 => n5591, A4 => 
                           n5590, ZN => n5604);
   U7357 : AOI22_X1 port map( A1 => IF_Regsxreg_file_615_port, A2 => n6153, B1 
                           => IF_Regsxreg_file_743_port, B2 => n6150, ZN => 
                           n5597);
   U7358 : AOI22_X1 port map( A1 => IF_Regsxreg_file_231_port, A2 => n6152, B1 
                           => IF_Regsxreg_file_967_port, B2 => n6154, ZN => 
                           n5596);
   U7359 : AOI22_X1 port map( A1 => IF_Regsxreg_file_455_port, A2 => n6155, B1 
                           => IF_Regsxreg_file_583_port, B2 => n6151, ZN => 
                           n5595);
   U7360 : AOI22_X1 port map( A1 => IF_Regsxreg_file_199_port, A2 => n5826, B1 
                           => IF_Regsxreg_file_103_port, B2 => n6129, ZN => 
                           n5594);
   U7361 : NAND4_X1 port map( A1 => n5597, A2 => n5596, A3 => n5595, A4 => 
                           n5594, ZN => n5603);
   U7362 : AOI22_X1 port map( A1 => IF_Regsxreg_file_775_port, A2 => n6135, B1 
                           => IF_Regsxreg_file_839_port, B2 => n6148, ZN => 
                           n5601);
   U7363 : AOI22_X1 port map( A1 => IF_Regsxreg_file_519_port, A2 => n6080, B1 
                           => IF_Regsxreg_file_263_port, B2 => n6160, ZN => 
                           n5600);
   U7364 : AOI22_X1 port map( A1 => IF_Regsxreg_file_135_port, A2 => n6115, B1 
                           => IF_Regsxreg_file_7_port, B2 => n6165, ZN => n5599
                           );
   U7365 : AOI22_X1 port map( A1 => IF_Regsxreg_file_903_port, A2 => n6167, B1 
                           => IF_Regsxreg_file_647_port, B2 => n5895, ZN => 
                           n5598);
   U7366 : NAND4_X1 port map( A1 => n5601, A2 => n5600, A3 => n5599, A4 => 
                           n5598, ZN => n5602);
   U7367 : AOI211_X1 port map( C1 => n5626, C2 => n5604, A => n5603, B => n5602
                           , ZN => n5605);
   U7368 : AOI21_X1 port map( B1 => n5606, B2 => n5605, A => n5968, ZN => 
                           IF_RegsxN602);
   U7369 : CLKBUF_X1 port map( A => n6167, Z => n5996);
   U7370 : AOI22_X1 port map( A1 => IF_Regsxreg_file_488_port, A2 => n6015, B1 
                           => IF_Regsxreg_file_712_port, B2 => n6109, ZN => 
                           n5609);
   U7371 : AOI22_X1 port map( A1 => IF_Regsxreg_file_616_port, A2 => n6153, B1 
                           => IF_Regsxreg_file_200_port, B2 => n5826, ZN => 
                           n5608);
   U7372 : AOI22_X1 port map( A1 => IF_Regsxreg_file_968_port, A2 => n6154, B1 
                           => IF_Regsxreg_file_104_port, B2 => n6129, ZN => 
                           n5607);
   U7373 : NAND3_X1 port map( A1 => n5609, A2 => n5608, A3 => n5607, ZN => 
                           n5610);
   U7374 : AOI21_X1 port map( B1 => IF_Regsxreg_file_904_port, B2 => n5996, A 
                           => n5610, ZN => n5628);
   U7375 : AOI22_X1 port map( A1 => IF_Regsxreg_file_680_port, A2 => n6140, B1 
                           => IF_Regsxreg_file_40_port, B2 => n6068, ZN => 
                           n5614);
   U7376 : AOI22_X1 port map( A1 => IF_Regsxreg_file_808_port, A2 => n6137, B1 
                           => IF_Regsxreg_file_296_port, B2 => n6141, ZN => 
                           n5613);
   U7377 : AOI22_X1 port map( A1 => IF_Regsxreg_file_424_port, A2 => n6099, B1 
                           => IF_Regsxreg_file_168_port, B2 => n6139, ZN => 
                           n5612);
   U7378 : AOI22_X1 port map( A1 => IF_Regsxreg_file_936_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_552_port, B2 => n6143, ZN => 
                           n5611);
   U7379 : NAND4_X1 port map( A1 => n5614, A2 => n5613, A3 => n5612, A4 => 
                           n5611, ZN => n5625);
   U7380 : AOI22_X1 port map( A1 => IF_Regsxreg_file_360_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_840_port, B2 => n6148, ZN => 
                           n5618);
   U7381 : AOI22_X1 port map( A1 => IF_Regsxreg_file_456_port, A2 => n6106, B1 
                           => IF_Regsxreg_file_872_port, B2 => n6128, ZN => 
                           n5617);
   U7382 : AOI22_X1 port map( A1 => IF_Regsxreg_file_584_port, A2 => n6151, B1 
                           => IF_Regsxreg_file_328_port, B2 => n6161, ZN => 
                           n5616);
   U7383 : AOI22_X1 port map( A1 => IF_Regsxreg_file_744_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_72_port, B2 => n6149, ZN => 
                           n5615);
   U7384 : NAND4_X1 port map( A1 => n5618, A2 => n5617, A3 => n5616, A4 => 
                           n5615, ZN => n5624);
   U7385 : AOI22_X1 port map( A1 => IF_Regsxreg_file_776_port, A2 => n6135, B1 
                           => IF_Regsxreg_file_232_port, B2 => n6046, ZN => 
                           n5622);
   U7386 : AOI22_X1 port map( A1 => IF_Regsxreg_file_136_port, A2 => n6115, B1 
                           => IF_Regsxreg_file_264_port, B2 => n6160, ZN => 
                           n5621);
   U7387 : AOI22_X1 port map( A1 => IF_Regsxreg_file_392_port, A2 => n6079, B1 
                           => IF_Regsxreg_file_8_port, B2 => n6052, ZN => n5620
                           );
   U7388 : AOI22_X1 port map( A1 => IF_Regsxreg_file_648_port, A2 => n6166, B1 
                           => IF_Regsxreg_file_520_port, B2 => n6080, ZN => 
                           n5619);
   U7389 : NAND4_X1 port map( A1 => n5622, A2 => n5621, A3 => n5620, A4 => 
                           n5619, ZN => n5623);
   U7390 : AOI211_X1 port map( C1 => n5626, C2 => n5625, A => n5624, B => n5623
                           , ZN => n5627);
   U7391 : AOI21_X1 port map( B1 => n5628, B2 => n5627, A => n5968, ZN => 
                           IF_RegsxN603);
   U7392 : AOI22_X1 port map( A1 => IF_Regsxreg_file_489_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_73_port, B2 => n6149, ZN => 
                           n5631);
   U7393 : AOI22_X1 port map( A1 => IF_Regsxreg_file_201_port, A2 => n6125, B1 
                           => IF_Regsxreg_file_233_port, B2 => n6046, ZN => 
                           n5630);
   U7394 : AOI22_X1 port map( A1 => IF_Regsxreg_file_585_port, A2 => n6151, B1 
                           => IF_Regsxreg_file_361_port, B2 => n6108, ZN => 
                           n5629);
   U7395 : NAND3_X1 port map( A1 => n5631, A2 => n5630, A3 => n5629, ZN => 
                           n5632);
   U7396 : AOI21_X1 port map( B1 => IF_Regsxreg_file_9_port, B2 => n6052, A => 
                           n5632, ZN => n5649);
   U7397 : AOI22_X1 port map( A1 => IF_Regsxreg_file_425_port, A2 => n6099, B1 
                           => IF_Regsxreg_file_681_port, B2 => n6041, ZN => 
                           n5636);
   U7398 : AOI22_X1 port map( A1 => IF_Regsxreg_file_937_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_169_port, B2 => n6139, ZN => 
                           n5635);
   U7399 : AOI22_X1 port map( A1 => IF_Regsxreg_file_297_port, A2 => n6098, B1 
                           => IF_Regsxreg_file_41_port, B2 => n6068, ZN => 
                           n5634);
   U7400 : AOI22_X1 port map( A1 => IF_Regsxreg_file_553_port, A2 => n6096, B1 
                           => IF_Regsxreg_file_809_port, B2 => n6137, ZN => 
                           n5633);
   U7401 : NAND4_X1 port map( A1 => n5636, A2 => n5635, A3 => n5634, A4 => 
                           n5633, ZN => n5647);
   U7402 : AOI22_X1 port map( A1 => IF_Regsxreg_file_969_port, A2 => n6154, B1 
                           => IF_Regsxreg_file_873_port, B2 => n6128, ZN => 
                           n5640);
   U7403 : AOI22_X1 port map( A1 => IF_Regsxreg_file_457_port, A2 => n6106, B1 
                           => IF_Regsxreg_file_105_port, B2 => n6129, ZN => 
                           n5639);
   U7404 : AOI22_X1 port map( A1 => IF_Regsxreg_file_841_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_713_port, B2 => n6127, ZN => 
                           n5638);
   U7405 : AOI22_X1 port map( A1 => IF_Regsxreg_file_617_port, A2 => n6005, B1 
                           => IF_Regsxreg_file_329_port, B2 => n6161, ZN => 
                           n5637);
   U7406 : NAND4_X1 port map( A1 => n5640, A2 => n5639, A3 => n5638, A4 => 
                           n5637, ZN => n5646);
   U7407 : AOI22_X1 port map( A1 => IF_Regsxreg_file_745_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_777_port, B2 => n6135, ZN => 
                           n5644);
   U7408 : AOI22_X1 port map( A1 => IF_Regsxreg_file_521_port, A2 => n6080, B1 
                           => IF_Regsxreg_file_265_port, B2 => n5952, ZN => 
                           n5643);
   U7409 : AOI22_X1 port map( A1 => IF_Regsxreg_file_905_port, A2 => n6167, B1 
                           => IF_Regsxreg_file_137_port, B2 => n6115, ZN => 
                           n5642);
   U7410 : AOI22_X1 port map( A1 => IF_Regsxreg_file_649_port, A2 => n6166, B1 
                           => IF_Regsxreg_file_393_port, B2 => n6163, ZN => 
                           n5641);
   U7411 : NAND4_X1 port map( A1 => n5644, A2 => n5643, A3 => n5642, A4 => 
                           n5641, ZN => n5645);
   U7412 : AOI211_X1 port map( C1 => n6267, C2 => n5647, A => n5646, B => n5645
                           , ZN => n5648);
   U7413 : AOI21_X1 port map( B1 => n5649, B2 => n5648, A => n5968, ZN => 
                           IF_RegsxN604);
   U7414 : AOI22_X1 port map( A1 => IF_Regsxreg_file_458_port, A2 => n6106, B1 
                           => IF_Regsxreg_file_490_port, B2 => n5926, ZN => 
                           n5652);
   U7415 : AOI22_X1 port map( A1 => IF_Regsxreg_file_746_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_970_port, B2 => n6154, ZN => 
                           n5651);
   U7416 : AOI22_X1 port map( A1 => IF_Regsxreg_file_106_port, A2 => n6129, B1 
                           => IF_Regsxreg_file_714_port, B2 => n6109, ZN => 
                           n5650);
   U7417 : NAND3_X1 port map( A1 => n5652, A2 => n5651, A3 => n5650, ZN => 
                           n5653);
   U7418 : AOI21_X1 port map( B1 => IF_Regsxreg_file_778_port, B2 => n6135, A 
                           => n5653, ZN => n5670);
   U7419 : AOI22_X1 port map( A1 => IF_Regsxreg_file_682_port, A2 => n6140, B1 
                           => IF_Regsxreg_file_554_port, B2 => n6143, ZN => 
                           n5657);
   U7420 : AOI22_X1 port map( A1 => IF_Regsxreg_file_42_port, A2 => n6068, B1 
                           => IF_Regsxreg_file_938_port, B2 => n5886, ZN => 
                           n5656);
   U7421 : AOI22_X1 port map( A1 => IF_Regsxreg_file_170_port, A2 => n6097, B1 
                           => IF_Regsxreg_file_810_port, B2 => n6067, ZN => 
                           n5655);
   U7422 : AOI22_X1 port map( A1 => IF_Regsxreg_file_298_port, A2 => n6141, B1 
                           => IF_Regsxreg_file_426_port, B2 => n6136, ZN => 
                           n5654);
   U7423 : NAND4_X1 port map( A1 => n5657, A2 => n5656, A3 => n5655, A4 => 
                           n5654, ZN => n5668);
   U7424 : AOI22_X1 port map( A1 => IF_Regsxreg_file_202_port, A2 => n6125, B1 
                           => IF_Regsxreg_file_74_port, B2 => n6149, ZN => 
                           n5661);
   U7425 : AOI22_X1 port map( A1 => IF_Regsxreg_file_234_port, A2 => n6152, B1 
                           => IF_Regsxreg_file_874_port, B2 => n6128, ZN => 
                           n5660);
   U7426 : AOI22_X1 port map( A1 => IF_Regsxreg_file_362_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_618_port, B2 => n6153, ZN => 
                           n5659);
   U7427 : AOI22_X1 port map( A1 => IF_Regsxreg_file_586_port, A2 => n6074, B1 
                           => IF_Regsxreg_file_330_port, B2 => n6161, ZN => 
                           n5658);
   U7428 : NAND4_X1 port map( A1 => n5661, A2 => n5660, A3 => n5659, A4 => 
                           n5658, ZN => n5667);
   U7429 : AOI22_X1 port map( A1 => IF_Regsxreg_file_842_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_138_port, B2 => n6115, ZN => 
                           n5665);
   U7430 : AOI22_X1 port map( A1 => IF_Regsxreg_file_394_port, A2 => n6163, B1 
                           => IF_Regsxreg_file_650_port, B2 => n5895, ZN => 
                           n5664);
   U7431 : AOI22_X1 port map( A1 => IF_Regsxreg_file_266_port, A2 => n6160, B1 
                           => IF_Regsxreg_file_906_port, B2 => n6167, ZN => 
                           n5663);
   U7432 : AOI22_X1 port map( A1 => IF_Regsxreg_file_10_port, A2 => n6165, B1 
                           => IF_Regsxreg_file_522_port, B2 => n6080, ZN => 
                           n5662);
   U7433 : NAND4_X1 port map( A1 => n5665, A2 => n5664, A3 => n5663, A4 => 
                           n5662, ZN => n5666);
   U7434 : AOI211_X1 port map( C1 => n6267, C2 => n5668, A => n5667, B => n5666
                           , ZN => n5669);
   U7435 : AOI21_X1 port map( B1 => n5670, B2 => n5669, A => n5968, ZN => 
                           IF_RegsxN605);
   U7436 : AOI22_X1 port map( A1 => IF_Regsxreg_file_491_port, A2 => n5926, B1 
                           => IF_Regsxreg_file_971_port, B2 => n6154, ZN => 
                           n5673);
   U7437 : AOI22_X1 port map( A1 => IF_Regsxreg_file_843_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_715_port, B2 => n6127, ZN => 
                           n5672);
   U7438 : AOI22_X1 port map( A1 => IF_Regsxreg_file_107_port, A2 => n6129, B1 
                           => IF_Regsxreg_file_459_port, B2 => n6155, ZN => 
                           n5671);
   U7439 : NAND3_X1 port map( A1 => n5673, A2 => n5672, A3 => n5671, ZN => 
                           n5674);
   U7440 : AOI21_X1 port map( B1 => IF_Regsxreg_file_907_port, B2 => n5996, A 
                           => n5674, ZN => n5691);
   U7441 : AOI22_X1 port map( A1 => IF_Regsxreg_file_939_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_299_port, B2 => n6141, ZN => 
                           n5678);
   U7442 : AOI22_X1 port map( A1 => IF_Regsxreg_file_427_port, A2 => n6099, B1 
                           => IF_Regsxreg_file_555_port, B2 => n6143, ZN => 
                           n5677);
   U7443 : AOI22_X1 port map( A1 => IF_Regsxreg_file_683_port, A2 => n6041, B1 
                           => IF_Regsxreg_file_811_port, B2 => n6137, ZN => 
                           n5676);
   U7444 : AOI22_X1 port map( A1 => IF_Regsxreg_file_43_port, A2 => n6142, B1 
                           => IF_Regsxreg_file_171_port, B2 => n6139, ZN => 
                           n5675);
   U7445 : NAND4_X1 port map( A1 => n5678, A2 => n5677, A3 => n5676, A4 => 
                           n5675, ZN => n5689);
   U7446 : AOI22_X1 port map( A1 => IF_Regsxreg_file_363_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_75_port, B2 => n6149, ZN => 
                           n5682);
   U7447 : AOI22_X1 port map( A1 => IF_Regsxreg_file_331_port, A2 => n6104, B1 
                           => IF_Regsxreg_file_587_port, B2 => n6151, ZN => 
                           n5681);
   U7448 : AOI22_X1 port map( A1 => IF_Regsxreg_file_235_port, A2 => n6046, B1 
                           => IF_Regsxreg_file_747_port, B2 => n6091, ZN => 
                           n5680);
   U7449 : AOI22_X1 port map( A1 => IF_Regsxreg_file_619_port, A2 => n6005, B1 
                           => IF_Regsxreg_file_203_port, B2 => n6125, ZN => 
                           n5679);
   U7450 : NAND4_X1 port map( A1 => n5682, A2 => n5681, A3 => n5680, A4 => 
                           n5679, ZN => n5688);
   U7451 : AOI22_X1 port map( A1 => IF_Regsxreg_file_875_port, A2 => n6128, B1 
                           => IF_Regsxreg_file_139_port, B2 => n6115, ZN => 
                           n5686);
   U7452 : AOI22_X1 port map( A1 => IF_Regsxreg_file_523_port, A2 => n6080, B1 
                           => IF_Regsxreg_file_651_port, B2 => n5895, ZN => 
                           n5685);
   U7453 : AOI22_X1 port map( A1 => IF_Regsxreg_file_395_port, A2 => n6079, B1 
                           => IF_Regsxreg_file_11_port, B2 => n6165, ZN => 
                           n5684);
   U7454 : AOI22_X1 port map( A1 => IF_Regsxreg_file_267_port, A2 => n6160, B1 
                           => IF_Regsxreg_file_779_port, B2 => n6135, ZN => 
                           n5683);
   U7455 : NAND4_X1 port map( A1 => n5686, A2 => n5685, A3 => n5684, A4 => 
                           n5683, ZN => n5687);
   U7456 : AOI211_X1 port map( C1 => n6267, C2 => n5689, A => n5688, B => n5687
                           , ZN => n5690);
   U7457 : AOI21_X1 port map( B1 => n5691, B2 => n5690, A => n5968, ZN => 
                           IF_RegsxN606);
   U7458 : CLKBUF_X1 port map( A => n6090, Z => n6073);
   U7459 : AOI22_X1 port map( A1 => IF_Regsxreg_file_972_port, A2 => n6073, B1 
                           => IF_Regsxreg_file_492_port, B2 => n5926, ZN => 
                           n5694);
   U7460 : AOI22_X1 port map( A1 => IF_Regsxreg_file_460_port, A2 => n6106, B1 
                           => IF_Regsxreg_file_108_port, B2 => n6129, ZN => 
                           n5693);
   U7461 : AOI22_X1 port map( A1 => IF_Regsxreg_file_620_port, A2 => n6153, B1 
                           => IF_Regsxreg_file_588_port, B2 => n6151, ZN => 
                           n5692);
   U7462 : NAND3_X1 port map( A1 => n5694, A2 => n5693, A3 => n5692, ZN => 
                           n5695);
   U7463 : AOI21_X1 port map( B1 => IF_Regsxreg_file_268_port, B2 => n5952, A 
                           => n5695, ZN => n5712);
   U7464 : AOI22_X1 port map( A1 => IF_Regsxreg_file_556_port, A2 => n6143, B1 
                           => IF_Regsxreg_file_684_port, B2 => n6041, ZN => 
                           n5699);
   U7465 : AOI22_X1 port map( A1 => IF_Regsxreg_file_940_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_812_port, B2 => n6067, ZN => 
                           n5698);
   U7466 : AOI22_X1 port map( A1 => IF_Regsxreg_file_172_port, A2 => n6097, B1 
                           => IF_Regsxreg_file_300_port, B2 => n6098, ZN => 
                           n5697);
   U7467 : AOI22_X1 port map( A1 => IF_Regsxreg_file_44_port, A2 => n6142, B1 
                           => IF_Regsxreg_file_428_port, B2 => n6136, ZN => 
                           n5696);
   U7468 : NAND4_X1 port map( A1 => n5699, A2 => n5698, A3 => n5697, A4 => 
                           n5696, ZN => n5710);
   U7469 : AOI22_X1 port map( A1 => IF_Regsxreg_file_204_port, A2 => n6125, B1 
                           => IF_Regsxreg_file_844_port, B2 => n6148, ZN => 
                           n5703);
   U7470 : AOI22_X1 port map( A1 => IF_Regsxreg_file_876_port, A2 => n6128, B1 
                           => IF_Regsxreg_file_236_port, B2 => n6046, ZN => 
                           n5702);
   U7471 : AOI22_X1 port map( A1 => IF_Regsxreg_file_364_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_716_port, B2 => n6127, ZN => 
                           n5701);
   U7472 : AOI22_X1 port map( A1 => IF_Regsxreg_file_76_port, A2 => n6062, B1 
                           => IF_Regsxreg_file_748_port, B2 => n6091, ZN => 
                           n5700);
   U7473 : NAND4_X1 port map( A1 => n5703, A2 => n5702, A3 => n5701, A4 => 
                           n5700, ZN => n5709);
   U7474 : AOI22_X1 port map( A1 => IF_Regsxreg_file_332_port, A2 => n6161, B1 
                           => IF_Regsxreg_file_780_port, B2 => n6135, ZN => 
                           n5707);
   U7475 : AOI22_X1 port map( A1 => IF_Regsxreg_file_396_port, A2 => n6163, B1 
                           => IF_Regsxreg_file_12_port, B2 => n6165, ZN => 
                           n5706);
   U7476 : AOI22_X1 port map( A1 => IF_Regsxreg_file_524_port, A2 => n6080, B1 
                           => IF_Regsxreg_file_652_port, B2 => n5895, ZN => 
                           n5705);
   U7477 : AOI22_X1 port map( A1 => IF_Regsxreg_file_908_port, A2 => n6167, B1 
                           => IF_Regsxreg_file_140_port, B2 => n6115, ZN => 
                           n5704);
   U7478 : NAND4_X1 port map( A1 => n5707, A2 => n5706, A3 => n5705, A4 => 
                           n5704, ZN => n5708);
   U7479 : AOI211_X1 port map( C1 => n6267, C2 => n5710, A => n5709, B => n5708
                           , ZN => n5711);
   U7480 : AOI21_X1 port map( B1 => n5712, B2 => n5711, A => n5968, ZN => 
                           IF_RegsxN607);
   U7481 : AOI22_X1 port map( A1 => IF_Regsxreg_file_493_port, A2 => n5926, B1 
                           => IF_Regsxreg_file_461_port, B2 => n6155, ZN => 
                           n5715);
   U7482 : AOI22_X1 port map( A1 => IF_Regsxreg_file_749_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_589_port, B2 => n6151, ZN => 
                           n5714);
   U7483 : AOI22_X1 port map( A1 => IF_Regsxreg_file_845_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_333_port, B2 => n6161, ZN => 
                           n5713);
   U7484 : NAND3_X1 port map( A1 => n5715, A2 => n5714, A3 => n5713, ZN => 
                           n5716);
   U7485 : AOI21_X1 port map( B1 => IF_Regsxreg_file_269_port, B2 => n5952, A 
                           => n5716, ZN => n5733);
   U7486 : AOI22_X1 port map( A1 => IF_Regsxreg_file_941_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_45_port, B2 => n6068, ZN => 
                           n5720);
   U7487 : AOI22_X1 port map( A1 => IF_Regsxreg_file_685_port, A2 => n6140, B1 
                           => IF_Regsxreg_file_173_port, B2 => n6139, ZN => 
                           n5719);
   U7488 : AOI22_X1 port map( A1 => IF_Regsxreg_file_429_port, A2 => n6099, B1 
                           => IF_Regsxreg_file_301_port, B2 => n6098, ZN => 
                           n5718);
   U7489 : AOI22_X1 port map( A1 => IF_Regsxreg_file_813_port, A2 => n6067, B1 
                           => IF_Regsxreg_file_557_port, B2 => n6143, ZN => 
                           n5717);
   U7490 : NAND4_X1 port map( A1 => n5720, A2 => n5719, A3 => n5718, A4 => 
                           n5717, ZN => n5731);
   U7491 : AOI22_X1 port map( A1 => IF_Regsxreg_file_621_port, A2 => n6005, B1 
                           => IF_Regsxreg_file_365_port, B2 => n6130, ZN => 
                           n5724);
   U7492 : AOI22_X1 port map( A1 => IF_Regsxreg_file_877_port, A2 => n6128, B1 
                           => IF_Regsxreg_file_237_port, B2 => n6046, ZN => 
                           n5723);
   U7493 : AOI22_X1 port map( A1 => IF_Regsxreg_file_205_port, A2 => n5826, B1 
                           => IF_Regsxreg_file_77_port, B2 => n6149, ZN => 
                           n5722);
   U7494 : AOI22_X1 port map( A1 => IF_Regsxreg_file_109_port, A2 => n6114, B1 
                           => IF_Regsxreg_file_973_port, B2 => n6154, ZN => 
                           n5721);
   U7495 : NAND4_X1 port map( A1 => n5724, A2 => n5723, A3 => n5722, A4 => 
                           n5721, ZN => n5730);
   U7496 : AOI22_X1 port map( A1 => IF_Regsxreg_file_717_port, A2 => n6127, B1 
                           => IF_Regsxreg_file_397_port, B2 => n6163, ZN => 
                           n5728);
   U7497 : AOI22_X1 port map( A1 => IF_Regsxreg_file_13_port, A2 => n6165, B1 
                           => IF_Regsxreg_file_909_port, B2 => n6167, ZN => 
                           n5727);
   U7498 : AOI22_X1 port map( A1 => IF_Regsxreg_file_141_port, A2 => n6115, B1 
                           => IF_Regsxreg_file_525_port, B2 => n6080, ZN => 
                           n5726);
   U7499 : AOI22_X1 port map( A1 => IF_Regsxreg_file_781_port, A2 => n6135, B1 
                           => IF_Regsxreg_file_653_port, B2 => n5895, ZN => 
                           n5725);
   U7500 : NAND4_X1 port map( A1 => n5728, A2 => n5727, A3 => n5726, A4 => 
                           n5725, ZN => n5729);
   U7501 : AOI211_X1 port map( C1 => n6267, C2 => n5731, A => n5730, B => n5729
                           , ZN => n5732);
   U7502 : AOI21_X1 port map( B1 => n5733, B2 => n5732, A => n5968, ZN => 
                           IF_RegsxN608);
   U7503 : AOI22_X1 port map( A1 => IF_Regsxreg_file_494_port, A2 => n6015, B1 
                           => IF_Regsxreg_file_206_port, B2 => n5826, ZN => 
                           n5736);
   U7504 : AOI22_X1 port map( A1 => IF_Regsxreg_file_750_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_878_port, B2 => n6128, ZN => 
                           n5735);
   U7505 : AOI22_X1 port map( A1 => IF_Regsxreg_file_974_port, A2 => n6073, B1 
                           => IF_Regsxreg_file_334_port, B2 => n6161, ZN => 
                           n5734);
   U7506 : NAND3_X1 port map( A1 => n5736, A2 => n5735, A3 => n5734, ZN => 
                           n5737);
   U7507 : AOI21_X1 port map( B1 => IF_Regsxreg_file_654_port, B2 => n6166, A 
                           => n5737, ZN => n5754);
   U7508 : AOI22_X1 port map( A1 => IF_Regsxreg_file_302_port, A2 => n6098, B1 
                           => IF_Regsxreg_file_430_port, B2 => n6136, ZN => 
                           n5741);
   U7509 : AOI22_X1 port map( A1 => IF_Regsxreg_file_814_port, A2 => n6137, B1 
                           => IF_Regsxreg_file_46_port, B2 => n6068, ZN => 
                           n5740);
   U7510 : AOI22_X1 port map( A1 => IF_Regsxreg_file_174_port, A2 => n6139, B1 
                           => IF_Regsxreg_file_558_port, B2 => n6096, ZN => 
                           n5739);
   U7511 : AOI22_X1 port map( A1 => IF_Regsxreg_file_942_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_686_port, B2 => n6140, ZN => 
                           n5738);
   U7512 : NAND4_X1 port map( A1 => n5741, A2 => n5740, A3 => n5739, A4 => 
                           n5738, ZN => n5752);
   U7513 : AOI22_X1 port map( A1 => IF_Regsxreg_file_718_port, A2 => n6109, B1 
                           => IF_Regsxreg_file_110_port, B2 => n6129, ZN => 
                           n5745);
   U7514 : AOI22_X1 port map( A1 => IF_Regsxreg_file_366_port, A2 => n6108, B1 
                           => IF_Regsxreg_file_238_port, B2 => n6046, ZN => 
                           n5744);
   U7515 : AOI22_X1 port map( A1 => IF_Regsxreg_file_78_port, A2 => n6062, B1 
                           => IF_Regsxreg_file_622_port, B2 => n6153, ZN => 
                           n5743);
   U7516 : AOI22_X1 port map( A1 => IF_Regsxreg_file_462_port, A2 => n6155, B1 
                           => IF_Regsxreg_file_590_port, B2 => n6151, ZN => 
                           n5742);
   U7517 : NAND4_X1 port map( A1 => n5745, A2 => n5744, A3 => n5743, A4 => 
                           n5742, ZN => n5751);
   U7518 : AOI22_X1 port map( A1 => IF_Regsxreg_file_846_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_782_port, B2 => n6051, ZN => 
                           n5749);
   U7519 : AOI22_X1 port map( A1 => IF_Regsxreg_file_526_port, A2 => n6080, B1 
                           => IF_Regsxreg_file_910_port, B2 => n6167, ZN => 
                           n5748);
   U7520 : AOI22_X1 port map( A1 => IF_Regsxreg_file_14_port, A2 => n6165, B1 
                           => IF_Regsxreg_file_270_port, B2 => n5952, ZN => 
                           n5747);
   U7521 : AOI22_X1 port map( A1 => IF_Regsxreg_file_142_port, A2 => n6115, B1 
                           => IF_Regsxreg_file_398_port, B2 => n6163, ZN => 
                           n5746);
   U7522 : NAND4_X1 port map( A1 => n5749, A2 => n5748, A3 => n5747, A4 => 
                           n5746, ZN => n5750);
   U7523 : AOI211_X1 port map( C1 => n6267, C2 => n5752, A => n5751, B => n5750
                           , ZN => n5753);
   U7524 : AOI21_X1 port map( B1 => n5754, B2 => n5753, A => n5968, ZN => 
                           IF_RegsxN609);
   U7525 : AOI22_X1 port map( A1 => IF_Regsxreg_file_495_port, A2 => n5926, B1 
                           => IF_Regsxreg_file_207_port, B2 => n6125, ZN => 
                           n5757);
   U7526 : AOI22_X1 port map( A1 => IF_Regsxreg_file_111_port, A2 => n6129, B1 
                           => IF_Regsxreg_file_79_port, B2 => n6149, ZN => 
                           n5756);
   U7527 : AOI22_X1 port map( A1 => IF_Regsxreg_file_751_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_463_port, B2 => n6155, ZN => 
                           n5755);
   U7528 : NAND3_X1 port map( A1 => n5757, A2 => n5756, A3 => n5755, ZN => 
                           n5758);
   U7529 : AOI21_X1 port map( B1 => IF_Regsxreg_file_527_port, B2 => n6162, A 
                           => n5758, ZN => n5775);
   U7530 : AOI22_X1 port map( A1 => IF_Regsxreg_file_943_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_815_port, B2 => n6067, ZN => 
                           n5762);
   U7531 : AOI22_X1 port map( A1 => IF_Regsxreg_file_687_port, A2 => n6140, B1 
                           => IF_Regsxreg_file_303_port, B2 => n6098, ZN => 
                           n5761);
   U7532 : AOI22_X1 port map( A1 => IF_Regsxreg_file_175_port, A2 => n6097, B1 
                           => IF_Regsxreg_file_431_port, B2 => n6136, ZN => 
                           n5760);
   U7533 : AOI22_X1 port map( A1 => IF_Regsxreg_file_47_port, A2 => n6068, B1 
                           => IF_Regsxreg_file_559_port, B2 => n6143, ZN => 
                           n5759);
   U7534 : NAND4_X1 port map( A1 => n5762, A2 => n5761, A3 => n5760, A4 => 
                           n5759, ZN => n5773);
   U7535 : AOI22_X1 port map( A1 => IF_Regsxreg_file_975_port, A2 => n6073, B1 
                           => IF_Regsxreg_file_719_port, B2 => n6127, ZN => 
                           n5766);
   U7536 : AOI22_X1 port map( A1 => IF_Regsxreg_file_623_port, A2 => n6005, B1 
                           => IF_Regsxreg_file_847_port, B2 => n6105, ZN => 
                           n5765);
   U7537 : AOI22_X1 port map( A1 => IF_Regsxreg_file_879_port, A2 => n6107, B1 
                           => IF_Regsxreg_file_335_port, B2 => n6161, ZN => 
                           n5764);
   U7538 : AOI22_X1 port map( A1 => IF_Regsxreg_file_591_port, A2 => n6074, B1 
                           => IF_Regsxreg_file_239_port, B2 => n6152, ZN => 
                           n5763);
   U7539 : NAND4_X1 port map( A1 => n5766, A2 => n5765, A3 => n5764, A4 => 
                           n5763, ZN => n5772);
   U7540 : AOI22_X1 port map( A1 => IF_Regsxreg_file_367_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_911_port, B2 => n5996, ZN => 
                           n5770);
   U7541 : AOI22_X1 port map( A1 => IF_Regsxreg_file_399_port, A2 => n6163, B1 
                           => IF_Regsxreg_file_143_port, B2 => n6115, ZN => 
                           n5769);
   U7542 : AOI22_X1 port map( A1 => IF_Regsxreg_file_271_port, A2 => n5952, B1 
                           => IF_Regsxreg_file_15_port, B2 => n6165, ZN => 
                           n5768);
   U7543 : AOI22_X1 port map( A1 => IF_Regsxreg_file_655_port, A2 => n6166, B1 
                           => IF_Regsxreg_file_783_port, B2 => n6051, ZN => 
                           n5767);
   U7544 : NAND4_X1 port map( A1 => n5770, A2 => n5769, A3 => n5768, A4 => 
                           n5767, ZN => n5771);
   U7545 : AOI211_X1 port map( C1 => n6267, C2 => n5773, A => n5772, B => n5771
                           , ZN => n5774);
   U7546 : AOI21_X1 port map( B1 => n5775, B2 => n5774, A => n5968, ZN => 
                           IF_RegsxN610);
   U7547 : AOI22_X1 port map( A1 => IF_Regsxreg_file_752_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_496_port, B2 => n5926, ZN => 
                           n5778);
   U7548 : AOI22_X1 port map( A1 => IF_Regsxreg_file_368_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_464_port, B2 => n6155, ZN => 
                           n5777);
   U7549 : AOI22_X1 port map( A1 => IF_Regsxreg_file_848_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_592_port, B2 => n6151, ZN => 
                           n5776);
   U7550 : NAND3_X1 port map( A1 => n5778, A2 => n5777, A3 => n5776, ZN => 
                           n5779);
   U7551 : AOI21_X1 port map( B1 => IF_Regsxreg_file_16_port, B2 => n6052, A =>
                           n5779, ZN => n5796);
   U7552 : AOI22_X1 port map( A1 => IF_Regsxreg_file_432_port, A2 => n6099, B1 
                           => IF_Regsxreg_file_176_port, B2 => n6097, ZN => 
                           n5783);
   U7553 : AOI22_X1 port map( A1 => IF_Regsxreg_file_688_port, A2 => n6041, B1 
                           => IF_Regsxreg_file_816_port, B2 => n6067, ZN => 
                           n5782);
   U7554 : AOI22_X1 port map( A1 => IF_Regsxreg_file_560_port, A2 => n6143, B1 
                           => IF_Regsxreg_file_48_port, B2 => n6068, ZN => 
                           n5781);
   U7555 : AOI22_X1 port map( A1 => IF_Regsxreg_file_304_port, A2 => n6141, B1 
                           => IF_Regsxreg_file_944_port, B2 => n5886, ZN => 
                           n5780);
   U7556 : NAND4_X1 port map( A1 => n5783, A2 => n5782, A3 => n5781, A4 => 
                           n5780, ZN => n5794);
   U7557 : AOI22_X1 port map( A1 => IF_Regsxreg_file_720_port, A2 => n6127, B1 
                           => IF_Regsxreg_file_240_port, B2 => n6152, ZN => 
                           n5787);
   U7558 : AOI22_X1 port map( A1 => IF_Regsxreg_file_80_port, A2 => n6149, B1 
                           => IF_Regsxreg_file_336_port, B2 => n6161, ZN => 
                           n5786);
   U7559 : AOI22_X1 port map( A1 => IF_Regsxreg_file_880_port, A2 => n6107, B1 
                           => IF_Regsxreg_file_624_port, B2 => n6005, ZN => 
                           n5785);
   U7560 : AOI22_X1 port map( A1 => IF_Regsxreg_file_208_port, A2 => n5826, B1 
                           => IF_Regsxreg_file_976_port, B2 => n6073, ZN => 
                           n5784);
   U7561 : NAND4_X1 port map( A1 => n5787, A2 => n5786, A3 => n5785, A4 => 
                           n5784, ZN => n5793);
   U7562 : AOI22_X1 port map( A1 => IF_Regsxreg_file_112_port, A2 => n6129, B1 
                           => IF_Regsxreg_file_656_port, B2 => n5895, ZN => 
                           n5791);
   U7563 : AOI22_X1 port map( A1 => IF_Regsxreg_file_144_port, A2 => n6115, B1 
                           => IF_Regsxreg_file_784_port, B2 => n6051, ZN => 
                           n5790);
   U7564 : AOI22_X1 port map( A1 => IF_Regsxreg_file_272_port, A2 => n5952, B1 
                           => IF_Regsxreg_file_912_port, B2 => n5996, ZN => 
                           n5789);
   U7565 : AOI22_X1 port map( A1 => IF_Regsxreg_file_528_port, A2 => n6080, B1 
                           => IF_Regsxreg_file_400_port, B2 => n6163, ZN => 
                           n5788);
   U7566 : NAND4_X1 port map( A1 => n5791, A2 => n5790, A3 => n5789, A4 => 
                           n5788, ZN => n5792);
   U7567 : AOI211_X1 port map( C1 => n6267, C2 => n5794, A => n5793, B => n5792
                           , ZN => n5795);
   U7568 : AOI21_X1 port map( B1 => n5796, B2 => n5795, A => n5968, ZN => 
                           IF_RegsxN611);
   U7569 : AOI22_X1 port map( A1 => IF_Regsxreg_file_497_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_337_port, B2 => n6161, ZN => 
                           n5799);
   U7570 : AOI22_X1 port map( A1 => IF_Regsxreg_file_721_port, A2 => n6127, B1 
                           => IF_Regsxreg_file_369_port, B2 => n6130, ZN => 
                           n5798);
   U7571 : AOI22_X1 port map( A1 => IF_Regsxreg_file_625_port, A2 => n6153, B1 
                           => IF_Regsxreg_file_977_port, B2 => n6154, ZN => 
                           n5797);
   U7572 : NAND3_X1 port map( A1 => n5799, A2 => n5798, A3 => n5797, ZN => 
                           n5800);
   U7573 : AOI21_X1 port map( B1 => IF_Regsxreg_file_529_port, B2 => n6162, A 
                           => n5800, ZN => n5817);
   U7574 : AOI22_X1 port map( A1 => IF_Regsxreg_file_305_port, A2 => n6098, B1 
                           => IF_Regsxreg_file_689_port, B2 => n6041, ZN => 
                           n5804);
   U7575 : AOI22_X1 port map( A1 => IF_Regsxreg_file_817_port, A2 => n6067, B1 
                           => IF_Regsxreg_file_433_port, B2 => n6136, ZN => 
                           n5803);
   U7576 : AOI22_X1 port map( A1 => IF_Regsxreg_file_177_port, A2 => n6139, B1 
                           => IF_Regsxreg_file_945_port, B2 => n5886, ZN => 
                           n5802);
   U7577 : AOI22_X1 port map( A1 => IF_Regsxreg_file_561_port, A2 => n6143, B1 
                           => IF_Regsxreg_file_49_port, B2 => n6068, ZN => 
                           n5801);
   U7578 : NAND4_X1 port map( A1 => n5804, A2 => n5803, A3 => n5802, A4 => 
                           n5801, ZN => n5815);
   U7579 : AOI22_X1 port map( A1 => IF_Regsxreg_file_881_port, A2 => n6128, B1 
                           => IF_Regsxreg_file_113_port, B2 => n6129, ZN => 
                           n5808);
   U7580 : AOI22_X1 port map( A1 => IF_Regsxreg_file_753_port, A2 => n6150, B1 
                           => IF_Regsxreg_file_241_port, B2 => n6152, ZN => 
                           n5807);
   U7581 : AOI22_X1 port map( A1 => IF_Regsxreg_file_849_port, A2 => n6148, B1 
                           => IF_Regsxreg_file_465_port, B2 => n6106, ZN => 
                           n5806);
   U7582 : AOI22_X1 port map( A1 => IF_Regsxreg_file_81_port, A2 => n6062, B1 
                           => IF_Regsxreg_file_209_port, B2 => n6125, ZN => 
                           n5805);
   U7583 : NAND4_X1 port map( A1 => n5808, A2 => n5807, A3 => n5806, A4 => 
                           n5805, ZN => n5814);
   U7584 : AOI22_X1 port map( A1 => IF_Regsxreg_file_593_port, A2 => n6151, B1 
                           => IF_Regsxreg_file_913_port, B2 => n5996, ZN => 
                           n5812);
   U7585 : AOI22_X1 port map( A1 => IF_Regsxreg_file_273_port, A2 => n5952, B1 
                           => IF_Regsxreg_file_145_port, B2 => n6164, ZN => 
                           n5811);
   U7586 : AOI22_X1 port map( A1 => IF_Regsxreg_file_17_port, A2 => n6052, B1 
                           => IF_Regsxreg_file_401_port, B2 => n6163, ZN => 
                           n5810);
   U7587 : AOI22_X1 port map( A1 => IF_Regsxreg_file_657_port, A2 => n6166, B1 
                           => IF_Regsxreg_file_785_port, B2 => n6051, ZN => 
                           n5809);
   U7588 : NAND4_X1 port map( A1 => n5812, A2 => n5811, A3 => n5810, A4 => 
                           n5809, ZN => n5813);
   U7589 : AOI211_X1 port map( C1 => n6267, C2 => n5815, A => n5814, B => n5813
                           , ZN => n5816);
   U7590 : AOI21_X1 port map( B1 => n5817, B2 => n5816, A => n5968, ZN => 
                           IF_RegsxN612);
   U7591 : AOI22_X1 port map( A1 => IF_Regsxreg_file_498_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_338_port, B2 => n6161, ZN => 
                           n5820);
   U7592 : AOI22_X1 port map( A1 => IF_Regsxreg_file_466_port, A2 => n6106, B1 
                           => IF_Regsxreg_file_626_port, B2 => n6005, ZN => 
                           n5819);
   U7593 : AOI22_X1 port map( A1 => IF_Regsxreg_file_242_port, A2 => n6152, B1 
                           => IF_Regsxreg_file_594_port, B2 => n6151, ZN => 
                           n5818);
   U7594 : NAND3_X1 port map( A1 => n5820, A2 => n5819, A3 => n5818, ZN => 
                           n5821);
   U7595 : AOI21_X1 port map( B1 => IF_Regsxreg_file_402_port, B2 => n6163, A 
                           => n5821, ZN => n5839);
   U7596 : AOI22_X1 port map( A1 => IF_Regsxreg_file_178_port, A2 => n6139, B1 
                           => IF_Regsxreg_file_562_port, B2 => n6096, ZN => 
                           n5825);
   U7597 : AOI22_X1 port map( A1 => IF_Regsxreg_file_818_port, A2 => n6067, B1 
                           => IF_Regsxreg_file_690_port, B2 => n6041, ZN => 
                           n5824);
   U7598 : AOI22_X1 port map( A1 => IF_Regsxreg_file_946_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_434_port, B2 => n6136, ZN => 
                           n5823);
   U7599 : AOI22_X1 port map( A1 => IF_Regsxreg_file_306_port, A2 => n6141, B1 
                           => IF_Regsxreg_file_50_port, B2 => n6068, ZN => 
                           n5822);
   U7600 : NAND4_X1 port map( A1 => n5825, A2 => n5824, A3 => n5823, A4 => 
                           n5822, ZN => n5837);
   U7601 : AOI22_X1 port map( A1 => IF_Regsxreg_file_882_port, A2 => n6128, B1 
                           => IF_Regsxreg_file_722_port, B2 => n6127, ZN => 
                           n5830);
   U7602 : AOI22_X1 port map( A1 => IF_Regsxreg_file_82_port, A2 => n6062, B1 
                           => IF_Regsxreg_file_850_port, B2 => n6105, ZN => 
                           n5829);
   U7603 : AOI22_X1 port map( A1 => IF_Regsxreg_file_210_port, A2 => n5826, B1 
                           => IF_Regsxreg_file_114_port, B2 => n6129, ZN => 
                           n5828);
   U7604 : AOI22_X1 port map( A1 => IF_Regsxreg_file_978_port, A2 => n6073, B1 
                           => IF_Regsxreg_file_370_port, B2 => n6130, ZN => 
                           n5827);
   U7605 : NAND4_X1 port map( A1 => n5830, A2 => n5829, A3 => n5828, A4 => 
                           n5827, ZN => n5836);
   U7606 : AOI22_X1 port map( A1 => IF_Regsxreg_file_754_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_658_port, B2 => n5895, ZN => 
                           n5834);
   U7607 : AOI22_X1 port map( A1 => IF_Regsxreg_file_530_port, A2 => n6080, B1 
                           => IF_Regsxreg_file_914_port, B2 => n5996, ZN => 
                           n5833);
   U7608 : AOI22_X1 port map( A1 => IF_Regsxreg_file_786_port, A2 => n6135, B1 
                           => IF_Regsxreg_file_18_port, B2 => n6165, ZN => 
                           n5832);
   U7609 : AOI22_X1 port map( A1 => IF_Regsxreg_file_146_port, A2 => n6115, B1 
                           => IF_Regsxreg_file_274_port, B2 => n5952, ZN => 
                           n5831);
   U7610 : NAND4_X1 port map( A1 => n5834, A2 => n5833, A3 => n5832, A4 => 
                           n5831, ZN => n5835);
   U7611 : AOI211_X1 port map( C1 => n6267, C2 => n5837, A => n5836, B => n5835
                           , ZN => n5838);
   U7612 : AOI21_X1 port map( B1 => n5839, B2 => n5838, A => n5968, ZN => 
                           IF_RegsxN613);
   U7613 : AOI22_X1 port map( A1 => IF_Regsxreg_file_339_port, A2 => n6161, B1 
                           => IF_Regsxreg_file_499_port, B2 => n5926, ZN => 
                           n5842);
   U7614 : AOI22_X1 port map( A1 => IF_Regsxreg_file_371_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_83_port, B2 => n6062, ZN => 
                           n5841);
   U7615 : AOI22_X1 port map( A1 => IF_Regsxreg_file_755_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_243_port, B2 => n6152, ZN => 
                           n5840);
   U7616 : NAND3_X1 port map( A1 => n5842, A2 => n5841, A3 => n5840, ZN => 
                           n5843);
   U7617 : AOI21_X1 port map( B1 => IF_Regsxreg_file_403_port, B2 => n6163, A 
                           => n5843, ZN => n5860);
   U7618 : AOI22_X1 port map( A1 => IF_Regsxreg_file_947_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_435_port, B2 => n6136, ZN => 
                           n5847);
   U7619 : AOI22_X1 port map( A1 => IF_Regsxreg_file_179_port, A2 => n6139, B1 
                           => IF_Regsxreg_file_563_port, B2 => n6096, ZN => 
                           n5846);
   U7620 : AOI22_X1 port map( A1 => IF_Regsxreg_file_307_port, A2 => n6141, B1 
                           => IF_Regsxreg_file_819_port, B2 => n6137, ZN => 
                           n5845);
   U7621 : AOI22_X1 port map( A1 => IF_Regsxreg_file_51_port, A2 => n6068, B1 
                           => IF_Regsxreg_file_691_port, B2 => n6140, ZN => 
                           n5844);
   U7622 : NAND4_X1 port map( A1 => n5847, A2 => n5846, A3 => n5845, A4 => 
                           n5844, ZN => n5858);
   U7623 : AOI22_X1 port map( A1 => IF_Regsxreg_file_595_port, A2 => n6151, B1 
                           => IF_Regsxreg_file_883_port, B2 => n6128, ZN => 
                           n5851);
   U7624 : AOI22_X1 port map( A1 => IF_Regsxreg_file_467_port, A2 => n6106, B1 
                           => IF_Regsxreg_file_115_port, B2 => n6129, ZN => 
                           n5850);
   U7625 : AOI22_X1 port map( A1 => IF_Regsxreg_file_851_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_211_port, B2 => n6125, ZN => 
                           n5849);
   U7626 : AOI22_X1 port map( A1 => IF_Regsxreg_file_723_port, A2 => n6109, B1 
                           => IF_Regsxreg_file_627_port, B2 => n6153, ZN => 
                           n5848);
   U7627 : NAND4_X1 port map( A1 => n5851, A2 => n5850, A3 => n5849, A4 => 
                           n5848, ZN => n5857);
   U7628 : AOI22_X1 port map( A1 => IF_Regsxreg_file_979_port, A2 => n6073, B1 
                           => IF_Regsxreg_file_659_port, B2 => n5895, ZN => 
                           n5855);
   U7629 : AOI22_X1 port map( A1 => IF_Regsxreg_file_147_port, A2 => n6115, B1 
                           => IF_Regsxreg_file_531_port, B2 => n6080, ZN => 
                           n5854);
   U7630 : AOI22_X1 port map( A1 => IF_Regsxreg_file_19_port, A2 => n6052, B1 
                           => IF_Regsxreg_file_915_port, B2 => n5996, ZN => 
                           n5853);
   U7631 : AOI22_X1 port map( A1 => IF_Regsxreg_file_275_port, A2 => n6160, B1 
                           => IF_Regsxreg_file_787_port, B2 => n6051, ZN => 
                           n5852);
   U7632 : NAND4_X1 port map( A1 => n5855, A2 => n5854, A3 => n5853, A4 => 
                           n5852, ZN => n5856);
   U7633 : AOI211_X1 port map( C1 => n6267, C2 => n5858, A => n5857, B => n5856
                           , ZN => n5859);
   U7634 : AOI21_X1 port map( B1 => n5860, B2 => n5859, A => n5968, ZN => 
                           IF_RegsxN614);
   U7635 : AOI22_X1 port map( A1 => IF_Regsxreg_file_500_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_468_port, B2 => n6155, ZN => 
                           n5863);
   U7636 : AOI22_X1 port map( A1 => IF_Regsxreg_file_372_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_724_port, B2 => n6127, ZN => 
                           n5862);
   U7637 : AOI22_X1 port map( A1 => IF_Regsxreg_file_244_port, A2 => n6152, B1 
                           => IF_Regsxreg_file_628_port, B2 => n6153, ZN => 
                           n5861);
   U7638 : NAND3_X1 port map( A1 => n5863, A2 => n5862, A3 => n5861, ZN => 
                           n5864);
   U7639 : AOI21_X1 port map( B1 => IF_Regsxreg_file_276_port, B2 => n5952, A 
                           => n5864, ZN => n5881);
   U7640 : AOI22_X1 port map( A1 => IF_Regsxreg_file_308_port, A2 => n6098, B1 
                           => IF_Regsxreg_file_820_port, B2 => n6137, ZN => 
                           n5868);
   U7641 : AOI22_X1 port map( A1 => IF_Regsxreg_file_564_port, A2 => n6143, B1 
                           => IF_Regsxreg_file_948_port, B2 => n5886, ZN => 
                           n5867);
   U7642 : AOI22_X1 port map( A1 => IF_Regsxreg_file_52_port, A2 => n6142, B1 
                           => IF_Regsxreg_file_180_port, B2 => n6097, ZN => 
                           n5866);
   U7643 : AOI22_X1 port map( A1 => IF_Regsxreg_file_692_port, A2 => n6041, B1 
                           => IF_Regsxreg_file_436_port, B2 => n6136, ZN => 
                           n5865);
   U7644 : NAND4_X1 port map( A1 => n5868, A2 => n5867, A3 => n5866, A4 => 
                           n5865, ZN => n5879);
   U7645 : AOI22_X1 port map( A1 => IF_Regsxreg_file_212_port, A2 => n6125, B1 
                           => IF_Regsxreg_file_756_port, B2 => n6091, ZN => 
                           n5872);
   U7646 : AOI22_X1 port map( A1 => IF_Regsxreg_file_884_port, A2 => n6107, B1 
                           => IF_Regsxreg_file_84_port, B2 => n6149, ZN => 
                           n5871);
   U7647 : AOI22_X1 port map( A1 => IF_Regsxreg_file_116_port, A2 => n6114, B1 
                           => IF_Regsxreg_file_596_port, B2 => n6151, ZN => 
                           n5870);
   U7648 : AOI22_X1 port map( A1 => IF_Regsxreg_file_980_port, A2 => n6073, B1 
                           => IF_Regsxreg_file_852_port, B2 => n6105, ZN => 
                           n5869);
   U7649 : NAND4_X1 port map( A1 => n5872, A2 => n5871, A3 => n5870, A4 => 
                           n5869, ZN => n5878);
   U7650 : AOI22_X1 port map( A1 => IF_Regsxreg_file_340_port, A2 => n6104, B1 
                           => IF_Regsxreg_file_660_port, B2 => n5895, ZN => 
                           n5876);
   U7651 : AOI22_X1 port map( A1 => IF_Regsxreg_file_532_port, A2 => n6162, B1 
                           => IF_Regsxreg_file_788_port, B2 => n6051, ZN => 
                           n5875);
   U7652 : AOI22_X1 port map( A1 => IF_Regsxreg_file_404_port, A2 => n6079, B1 
                           => IF_Regsxreg_file_916_port, B2 => n5996, ZN => 
                           n5874);
   U7653 : AOI22_X1 port map( A1 => IF_Regsxreg_file_20_port, A2 => n6052, B1 
                           => IF_Regsxreg_file_148_port, B2 => n6164, ZN => 
                           n5873);
   U7654 : NAND4_X1 port map( A1 => n5876, A2 => n5875, A3 => n5874, A4 => 
                           n5873, ZN => n5877);
   U7655 : AOI211_X1 port map( C1 => n6267, C2 => n5879, A => n5878, B => n5877
                           , ZN => n5880);
   U7656 : AOI21_X1 port map( B1 => n5881, B2 => n5880, A => n5968, ZN => 
                           IF_RegsxN615);
   U7657 : AOI22_X1 port map( A1 => IF_Regsxreg_file_501_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_629_port, B2 => n6153, ZN => 
                           n5884);
   U7658 : AOI22_X1 port map( A1 => IF_Regsxreg_file_981_port, A2 => n6073, B1 
                           => IF_Regsxreg_file_245_port, B2 => n6152, ZN => 
                           n5883);
   U7659 : AOI22_X1 port map( A1 => IF_Regsxreg_file_757_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_373_port, B2 => n6108, ZN => 
                           n5882);
   U7660 : NAND3_X1 port map( A1 => n5884, A2 => n5883, A3 => n5882, ZN => 
                           n5885);
   U7661 : AOI21_X1 port map( B1 => IF_Regsxreg_file_917_port, B2 => n5996, A 
                           => n5885, ZN => n5904);
   U7662 : AOI22_X1 port map( A1 => IF_Regsxreg_file_821_port, A2 => n6137, B1 
                           => IF_Regsxreg_file_949_port, B2 => n5886, ZN => 
                           n5890);
   U7663 : AOI22_X1 port map( A1 => IF_Regsxreg_file_693_port, A2 => n6041, B1 
                           => IF_Regsxreg_file_437_port, B2 => n6136, ZN => 
                           n5889);
   U7664 : AOI22_X1 port map( A1 => IF_Regsxreg_file_565_port, A2 => n6143, B1 
                           => IF_Regsxreg_file_53_port, B2 => n6142, ZN => 
                           n5888);
   U7665 : AOI22_X1 port map( A1 => IF_Regsxreg_file_309_port, A2 => n6141, B1 
                           => IF_Regsxreg_file_181_port, B2 => n6139, ZN => 
                           n5887);
   U7666 : NAND4_X1 port map( A1 => n5890, A2 => n5889, A3 => n5888, A4 => 
                           n5887, ZN => n5902);
   U7667 : AOI22_X1 port map( A1 => IF_Regsxreg_file_85_port, A2 => n6149, B1 
                           => IF_Regsxreg_file_597_port, B2 => n6074, ZN => 
                           n5894);
   U7668 : AOI22_X1 port map( A1 => IF_Regsxreg_file_341_port, A2 => n6104, B1 
                           => IF_Regsxreg_file_853_port, B2 => n6105, ZN => 
                           n5893);
   U7669 : AOI22_X1 port map( A1 => IF_Regsxreg_file_885_port, A2 => n6107, B1 
                           => IF_Regsxreg_file_213_port, B2 => n6125, ZN => 
                           n5892);
   U7670 : AOI22_X1 port map( A1 => IF_Regsxreg_file_117_port, A2 => n6114, B1 
                           => IF_Regsxreg_file_469_port, B2 => n6106, ZN => 
                           n5891);
   U7671 : NAND4_X1 port map( A1 => n5894, A2 => n5893, A3 => n5892, A4 => 
                           n5891, ZN => n5901);
   U7672 : AOI22_X1 port map( A1 => IF_Regsxreg_file_725_port, A2 => n6127, B1 
                           => IF_Regsxreg_file_533_port, B2 => n6080, ZN => 
                           n5899);
   U7673 : AOI22_X1 port map( A1 => IF_Regsxreg_file_149_port, A2 => n6115, B1 
                           => IF_Regsxreg_file_21_port, B2 => n6165, ZN => 
                           n5898);
   U7674 : AOI22_X1 port map( A1 => IF_Regsxreg_file_277_port, A2 => n6160, B1 
                           => IF_Regsxreg_file_661_port, B2 => n5895, ZN => 
                           n5897);
   U7675 : AOI22_X1 port map( A1 => IF_Regsxreg_file_789_port, A2 => n6135, B1 
                           => IF_Regsxreg_file_405_port, B2 => n6163, ZN => 
                           n5896);
   U7676 : NAND4_X1 port map( A1 => n5899, A2 => n5898, A3 => n5897, A4 => 
                           n5896, ZN => n5900);
   U7677 : AOI211_X1 port map( C1 => n6267, C2 => n5902, A => n5901, B => n5900
                           , ZN => n5903);
   U7678 : AOI21_X1 port map( B1 => n5904, B2 => n5903, A => n5968, ZN => 
                           IF_RegsxN616);
   U7679 : AOI22_X1 port map( A1 => IF_Regsxreg_file_502_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_726_port, B2 => n6127, ZN => 
                           n5907);
   U7680 : AOI22_X1 port map( A1 => IF_Regsxreg_file_758_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_86_port, B2 => n6149, ZN => 
                           n5906);
   U7681 : AOI22_X1 port map( A1 => IF_Regsxreg_file_374_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_630_port, B2 => n6153, ZN => 
                           n5905);
   U7682 : NAND3_X1 port map( A1 => n5907, A2 => n5906, A3 => n5905, ZN => 
                           n5908);
   U7683 : AOI21_X1 port map( B1 => IF_Regsxreg_file_790_port, B2 => n6135, A 
                           => n5908, ZN => n5925);
   U7684 : AOI22_X1 port map( A1 => IF_Regsxreg_file_310_port, A2 => n6098, B1 
                           => IF_Regsxreg_file_54_port, B2 => n6142, ZN => 
                           n5912);
   U7685 : AOI22_X1 port map( A1 => IF_Regsxreg_file_182_port, A2 => n6139, B1 
                           => IF_Regsxreg_file_438_port, B2 => n6136, ZN => 
                           n5911);
   U7686 : AOI22_X1 port map( A1 => IF_Regsxreg_file_822_port, A2 => n6067, B1 
                           => IF_Regsxreg_file_950_port, B2 => n6138, ZN => 
                           n5910);
   U7687 : AOI22_X1 port map( A1 => IF_Regsxreg_file_566_port, A2 => n6143, B1 
                           => IF_Regsxreg_file_694_port, B2 => n6140, ZN => 
                           n5909);
   U7688 : NAND4_X1 port map( A1 => n5912, A2 => n5911, A3 => n5910, A4 => 
                           n5909, ZN => n5923);
   U7689 : AOI22_X1 port map( A1 => IF_Regsxreg_file_118_port, A2 => n6129, B1 
                           => IF_Regsxreg_file_214_port, B2 => n6125, ZN => 
                           n5916);
   U7690 : AOI22_X1 port map( A1 => IF_Regsxreg_file_854_port, A2 => n6148, B1 
                           => IF_Regsxreg_file_342_port, B2 => n6104, ZN => 
                           n5915);
   U7691 : AOI22_X1 port map( A1 => IF_Regsxreg_file_246_port, A2 => n6046, B1 
                           => IF_Regsxreg_file_886_port, B2 => n6128, ZN => 
                           n5914);
   U7692 : AOI22_X1 port map( A1 => IF_Regsxreg_file_598_port, A2 => n6074, B1 
                           => IF_Regsxreg_file_470_port, B2 => n6106, ZN => 
                           n5913);
   U7693 : NAND4_X1 port map( A1 => n5916, A2 => n5915, A3 => n5914, A4 => 
                           n5913, ZN => n5922);
   U7694 : AOI22_X1 port map( A1 => IF_Regsxreg_file_982_port, A2 => n6073, B1 
                           => IF_Regsxreg_file_534_port, B2 => n6162, ZN => 
                           n5920);
   U7695 : AOI22_X1 port map( A1 => IF_Regsxreg_file_918_port, A2 => n5996, B1 
                           => IF_Regsxreg_file_150_port, B2 => n6164, ZN => 
                           n5919);
   U7696 : AOI22_X1 port map( A1 => IF_Regsxreg_file_278_port, A2 => n6160, B1 
                           => IF_Regsxreg_file_406_port, B2 => n6163, ZN => 
                           n5918);
   U7697 : AOI22_X1 port map( A1 => IF_Regsxreg_file_662_port, A2 => n6166, B1 
                           => IF_Regsxreg_file_22_port, B2 => n6165, ZN => 
                           n5917);
   U7698 : NAND4_X1 port map( A1 => n5920, A2 => n5919, A3 => n5918, A4 => 
                           n5917, ZN => n5921);
   U7699 : AOI211_X1 port map( C1 => n6267, C2 => n5923, A => n5922, B => n5921
                           , ZN => n5924);
   U7700 : AOI21_X1 port map( B1 => n5925, B2 => n5924, A => n5968, ZN => 
                           IF_RegsxN617);
   U7701 : AOI22_X1 port map( A1 => IF_Regsxreg_file_343_port, A2 => n6161, B1 
                           => IF_Regsxreg_file_503_port, B2 => n5926, ZN => 
                           n5929);
   U7702 : AOI22_X1 port map( A1 => IF_Regsxreg_file_119_port, A2 => n6129, B1 
                           => IF_Regsxreg_file_247_port, B2 => n6152, ZN => 
                           n5928);
   U7703 : AOI22_X1 port map( A1 => IF_Regsxreg_file_855_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_983_port, B2 => n6090, ZN => 
                           n5927);
   U7704 : NAND3_X1 port map( A1 => n5929, A2 => n5928, A3 => n5927, ZN => 
                           n5930);
   U7705 : AOI21_X1 port map( B1 => IF_Regsxreg_file_279_port, B2 => n5952, A 
                           => n5930, ZN => n5947);
   U7706 : AOI22_X1 port map( A1 => IF_Regsxreg_file_439_port, A2 => n6099, B1 
                           => IF_Regsxreg_file_567_port, B2 => n6096, ZN => 
                           n5934);
   U7707 : AOI22_X1 port map( A1 => IF_Regsxreg_file_951_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_183_port, B2 => n6097, ZN => 
                           n5933);
   U7708 : AOI22_X1 port map( A1 => IF_Regsxreg_file_823_port, A2 => n6067, B1 
                           => IF_Regsxreg_file_55_port, B2 => n6142, ZN => 
                           n5932);
   U7709 : AOI22_X1 port map( A1 => IF_Regsxreg_file_311_port, A2 => n6141, B1 
                           => IF_Regsxreg_file_695_port, B2 => n6140, ZN => 
                           n5931);
   U7710 : NAND4_X1 port map( A1 => n5934, A2 => n5933, A3 => n5932, A4 => 
                           n5931, ZN => n5945);
   U7711 : AOI22_X1 port map( A1 => IF_Regsxreg_file_887_port, A2 => n6128, B1 
                           => IF_Regsxreg_file_727_port, B2 => n6127, ZN => 
                           n5938);
   U7712 : AOI22_X1 port map( A1 => IF_Regsxreg_file_375_port, A2 => n6108, B1 
                           => IF_Regsxreg_file_471_port, B2 => n6106, ZN => 
                           n5937);
   U7713 : AOI22_X1 port map( A1 => IF_Regsxreg_file_759_port, A2 => n6150, B1 
                           => IF_Regsxreg_file_631_port, B2 => n6153, ZN => 
                           n5936);
   U7714 : AOI22_X1 port map( A1 => IF_Regsxreg_file_87_port, A2 => n6062, B1 
                           => IF_Regsxreg_file_215_port, B2 => n6125, ZN => 
                           n5935);
   U7715 : NAND4_X1 port map( A1 => n5938, A2 => n5937, A3 => n5936, A4 => 
                           n5935, ZN => n5944);
   U7716 : AOI22_X1 port map( A1 => IF_Regsxreg_file_919_port, A2 => n5996, B1 
                           => IF_Regsxreg_file_599_port, B2 => n6074, ZN => 
                           n5942);
   U7717 : AOI22_X1 port map( A1 => IF_Regsxreg_file_791_port, A2 => n6135, B1 
                           => IF_Regsxreg_file_407_port, B2 => n6079, ZN => 
                           n5941);
   U7718 : AOI22_X1 port map( A1 => IF_Regsxreg_file_663_port, A2 => n6166, B1 
                           => IF_Regsxreg_file_535_port, B2 => n6162, ZN => 
                           n5940);
   U7719 : AOI22_X1 port map( A1 => IF_Regsxreg_file_23_port, A2 => n6052, B1 
                           => IF_Regsxreg_file_151_port, B2 => n6164, ZN => 
                           n5939);
   U7720 : NAND4_X1 port map( A1 => n5942, A2 => n5941, A3 => n5940, A4 => 
                           n5939, ZN => n5943);
   U7721 : AOI211_X1 port map( C1 => n6267, C2 => n5945, A => n5944, B => n5943
                           , ZN => n5946);
   U7722 : AOI21_X1 port map( B1 => n5947, B2 => n5946, A => n5968, ZN => 
                           IF_RegsxN618);
   U7723 : AOI22_X1 port map( A1 => IF_Regsxreg_file_504_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_728_port, B2 => n6127, ZN => 
                           n5950);
   U7724 : AOI22_X1 port map( A1 => IF_Regsxreg_file_216_port, A2 => n6125, B1 
                           => IF_Regsxreg_file_472_port, B2 => n6106, ZN => 
                           n5949);
   U7725 : AOI22_X1 port map( A1 => IF_Regsxreg_file_856_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_760_port, B2 => n6150, ZN => 
                           n5948);
   U7726 : NAND3_X1 port map( A1 => n5950, A2 => n5949, A3 => n5948, ZN => 
                           n5951);
   U7727 : AOI21_X1 port map( B1 => IF_Regsxreg_file_280_port, B2 => n5952, A 
                           => n5951, ZN => n5970);
   U7728 : AOI22_X1 port map( A1 => IF_Regsxreg_file_184_port, A2 => n6139, B1 
                           => IF_Regsxreg_file_440_port, B2 => n6136, ZN => 
                           n5956);
   U7729 : AOI22_X1 port map( A1 => IF_Regsxreg_file_696_port, A2 => n6140, B1 
                           => IF_Regsxreg_file_312_port, B2 => n6098, ZN => 
                           n5955);
   U7730 : AOI22_X1 port map( A1 => IF_Regsxreg_file_952_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_56_port, B2 => n6142, ZN => 
                           n5954);
   U7731 : AOI22_X1 port map( A1 => IF_Regsxreg_file_824_port, A2 => n6067, B1 
                           => IF_Regsxreg_file_568_port, B2 => n6096, ZN => 
                           n5953);
   U7732 : NAND4_X1 port map( A1 => n5956, A2 => n5955, A3 => n5954, A4 => 
                           n5953, ZN => n5967);
   U7733 : AOI22_X1 port map( A1 => IF_Regsxreg_file_344_port, A2 => n6104, B1 
                           => IF_Regsxreg_file_600_port, B2 => n6074, ZN => 
                           n5960);
   U7734 : AOI22_X1 port map( A1 => IF_Regsxreg_file_120_port, A2 => n6114, B1 
                           => IF_Regsxreg_file_632_port, B2 => n6153, ZN => 
                           n5959);
   U7735 : AOI22_X1 port map( A1 => IF_Regsxreg_file_248_port, A2 => n6046, B1 
                           => IF_Regsxreg_file_88_port, B2 => n6062, ZN => 
                           n5958);
   U7736 : AOI22_X1 port map( A1 => IF_Regsxreg_file_376_port, A2 => n6108, B1 
                           => IF_Regsxreg_file_888_port, B2 => n6128, ZN => 
                           n5957);
   U7737 : NAND4_X1 port map( A1 => n5960, A2 => n5959, A3 => n5958, A4 => 
                           n5957, ZN => n5966);
   U7738 : AOI22_X1 port map( A1 => IF_Regsxreg_file_984_port, A2 => n6073, B1 
                           => IF_Regsxreg_file_664_port, B2 => n6166, ZN => 
                           n5964);
   U7739 : AOI22_X1 port map( A1 => IF_Regsxreg_file_536_port, A2 => n6080, B1 
                           => IF_Regsxreg_file_408_port, B2 => n6079, ZN => 
                           n5963);
   U7740 : AOI22_X1 port map( A1 => IF_Regsxreg_file_792_port, A2 => n6135, B1 
                           => IF_Regsxreg_file_152_port, B2 => n6164, ZN => 
                           n5962);
   U7741 : AOI22_X1 port map( A1 => IF_Regsxreg_file_24_port, A2 => n6052, B1 
                           => IF_Regsxreg_file_920_port, B2 => n6167, ZN => 
                           n5961);
   U7742 : NAND4_X1 port map( A1 => n5964, A2 => n5963, A3 => n5962, A4 => 
                           n5961, ZN => n5965);
   U7743 : AOI211_X1 port map( C1 => n6267, C2 => n5967, A => n5966, B => n5965
                           , ZN => n5969);
   U7744 : CLKBUF_X1 port map( A => n5968, Z => n6175);
   U7745 : AOI21_X1 port map( B1 => n5970, B2 => n5969, A => n6175, ZN => 
                           IF_RegsxN619);
   U7746 : AOI22_X1 port map( A1 => IF_Regsxreg_file_505_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_377_port, B2 => n6108, ZN => 
                           n5973);
   U7747 : AOI22_X1 port map( A1 => IF_Regsxreg_file_633_port, A2 => n6153, B1 
                           => IF_Regsxreg_file_249_port, B2 => n6152, ZN => 
                           n5972);
   U7748 : AOI22_X1 port map( A1 => IF_Regsxreg_file_889_port, A2 => n6128, B1 
                           => IF_Regsxreg_file_121_port, B2 => n6114, ZN => 
                           n5971);
   U7749 : NAND3_X1 port map( A1 => n5973, A2 => n5972, A3 => n5971, ZN => 
                           n5974);
   U7750 : AOI21_X1 port map( B1 => IF_Regsxreg_file_665_port, B2 => n6166, A 
                           => n5974, ZN => n5991);
   U7751 : AOI22_X1 port map( A1 => IF_Regsxreg_file_825_port, A2 => n6137, B1 
                           => IF_Regsxreg_file_697_port, B2 => n6140, ZN => 
                           n5978);
   U7752 : AOI22_X1 port map( A1 => IF_Regsxreg_file_57_port, A2 => n6068, B1 
                           => IF_Regsxreg_file_953_port, B2 => n6138, ZN => 
                           n5977);
   U7753 : AOI22_X1 port map( A1 => IF_Regsxreg_file_185_port, A2 => n6139, B1 
                           => IF_Regsxreg_file_313_port, B2 => n6098, ZN => 
                           n5976);
   U7754 : AOI22_X1 port map( A1 => IF_Regsxreg_file_441_port, A2 => n6099, B1 
                           => IF_Regsxreg_file_569_port, B2 => n6096, ZN => 
                           n5975);
   U7755 : NAND4_X1 port map( A1 => n5978, A2 => n5977, A3 => n5976, A4 => 
                           n5975, ZN => n5989);
   U7756 : AOI22_X1 port map( A1 => IF_Regsxreg_file_217_port, A2 => n6125, B1 
                           => IF_Regsxreg_file_761_port, B2 => n6150, ZN => 
                           n5982);
   U7757 : AOI22_X1 port map( A1 => IF_Regsxreg_file_857_port, A2 => n6148, B1 
                           => IF_Regsxreg_file_473_port, B2 => n6106, ZN => 
                           n5981);
   U7758 : AOI22_X1 port map( A1 => IF_Regsxreg_file_729_port, A2 => n6109, B1 
                           => IF_Regsxreg_file_89_port, B2 => n6062, ZN => 
                           n5980);
   U7759 : AOI22_X1 port map( A1 => IF_Regsxreg_file_601_port, A2 => n6074, B1 
                           => IF_Regsxreg_file_345_port, B2 => n6161, ZN => 
                           n5979);
   U7760 : NAND4_X1 port map( A1 => n5982, A2 => n5981, A3 => n5980, A4 => 
                           n5979, ZN => n5988);
   U7761 : AOI22_X1 port map( A1 => IF_Regsxreg_file_985_port, A2 => n6073, B1 
                           => IF_Regsxreg_file_537_port, B2 => n6162, ZN => 
                           n5986);
   U7762 : AOI22_X1 port map( A1 => IF_Regsxreg_file_153_port, A2 => n6115, B1 
                           => IF_Regsxreg_file_793_port, B2 => n6051, ZN => 
                           n5985);
   U7763 : AOI22_X1 port map( A1 => IF_Regsxreg_file_921_port, A2 => n6167, B1 
                           => IF_Regsxreg_file_409_port, B2 => n6079, ZN => 
                           n5984);
   U7764 : AOI22_X1 port map( A1 => IF_Regsxreg_file_281_port, A2 => n6160, B1 
                           => IF_Regsxreg_file_25_port, B2 => n6052, ZN => 
                           n5983);
   U7765 : NAND4_X1 port map( A1 => n5986, A2 => n5985, A3 => n5984, A4 => 
                           n5983, ZN => n5987);
   U7766 : AOI211_X1 port map( C1 => n6267, C2 => n5989, A => n5988, B => n5987
                           , ZN => n5990);
   U7767 : AOI21_X1 port map( B1 => n5991, B2 => n5990, A => n6175, ZN => 
                           IF_RegsxN620);
   U7768 : AOI22_X1 port map( A1 => IF_Regsxreg_file_506_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_730_port, B2 => n6127, ZN => 
                           n5994);
   U7769 : AOI22_X1 port map( A1 => IF_Regsxreg_file_90_port, A2 => n6149, B1 
                           => IF_Regsxreg_file_890_port, B2 => n6107, ZN => 
                           n5993);
   U7770 : AOI22_X1 port map( A1 => IF_Regsxreg_file_474_port, A2 => n6106, B1 
                           => IF_Regsxreg_file_346_port, B2 => n6104, ZN => 
                           n5992);
   U7771 : NAND3_X1 port map( A1 => n5994, A2 => n5993, A3 => n5992, ZN => 
                           n5995);
   U7772 : AOI21_X1 port map( B1 => IF_Regsxreg_file_922_port, B2 => n5996, A 
                           => n5995, ZN => n6014);
   U7773 : AOI22_X1 port map( A1 => IF_Regsxreg_file_698_port, A2 => n6140, B1 
                           => IF_Regsxreg_file_826_port, B2 => n6137, ZN => 
                           n6000);
   U7774 : AOI22_X1 port map( A1 => IF_Regsxreg_file_570_port, A2 => n6143, B1 
                           => IF_Regsxreg_file_442_port, B2 => n6136, ZN => 
                           n5999);
   U7775 : AOI22_X1 port map( A1 => IF_Regsxreg_file_58_port, A2 => n6142, B1 
                           => IF_Regsxreg_file_314_port, B2 => n6098, ZN => 
                           n5998);
   U7776 : AOI22_X1 port map( A1 => IF_Regsxreg_file_954_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_186_port, B2 => n6139, ZN => 
                           n5997);
   U7777 : NAND4_X1 port map( A1 => n6000, A2 => n5999, A3 => n5998, A4 => 
                           n5997, ZN => n6012);
   U7778 : AOI22_X1 port map( A1 => IF_Regsxreg_file_986_port, A2 => n6073, B1 
                           => IF_Regsxreg_file_122_port, B2 => n6114, ZN => 
                           n6004);
   U7779 : AOI22_X1 port map( A1 => IF_Regsxreg_file_858_port, A2 => n6148, B1 
                           => IF_Regsxreg_file_250_port, B2 => n6152, ZN => 
                           n6003);
   U7780 : AOI22_X1 port map( A1 => IF_Regsxreg_file_762_port, A2 => n6150, B1 
                           => IF_Regsxreg_file_602_port, B2 => n6151, ZN => 
                           n6002);
   U7781 : AOI22_X1 port map( A1 => IF_Regsxreg_file_378_port, A2 => n6108, B1 
                           => IF_Regsxreg_file_218_port, B2 => n6125, ZN => 
                           n6001);
   U7782 : NAND4_X1 port map( A1 => n6004, A2 => n6003, A3 => n6002, A4 => 
                           n6001, ZN => n6011);
   U7783 : AOI22_X1 port map( A1 => IF_Regsxreg_file_634_port, A2 => n6005, B1 
                           => IF_Regsxreg_file_794_port, B2 => n6051, ZN => 
                           n6009);
   U7784 : AOI22_X1 port map( A1 => IF_Regsxreg_file_26_port, A2 => n6165, B1 
                           => IF_Regsxreg_file_154_port, B2 => n6164, ZN => 
                           n6008);
   U7785 : AOI22_X1 port map( A1 => IF_Regsxreg_file_410_port, A2 => n6079, B1 
                           => IF_Regsxreg_file_666_port, B2 => n6166, ZN => 
                           n6007);
   U7786 : AOI22_X1 port map( A1 => IF_Regsxreg_file_282_port, A2 => n6160, B1 
                           => IF_Regsxreg_file_538_port, B2 => n6162, ZN => 
                           n6006);
   U7787 : NAND4_X1 port map( A1 => n6009, A2 => n6008, A3 => n6007, A4 => 
                           n6006, ZN => n6010);
   U7788 : AOI211_X1 port map( C1 => n6267, C2 => n6012, A => n6011, B => n6010
                           , ZN => n6013);
   U7789 : AOI21_X1 port map( B1 => n6014, B2 => n6013, A => n6175, ZN => 
                           IF_RegsxN621);
   U7790 : AOI22_X1 port map( A1 => IF_Regsxreg_file_507_port, A2 => n6015, B1 
                           => IF_Regsxreg_file_603_port, B2 => n6074, ZN => 
                           n6018);
   U7791 : AOI22_X1 port map( A1 => IF_Regsxreg_file_891_port, A2 => n6128, B1 
                           => IF_Regsxreg_file_635_port, B2 => n6153, ZN => 
                           n6017);
   U7792 : AOI22_X1 port map( A1 => IF_Regsxreg_file_251_port, A2 => n6152, B1 
                           => IF_Regsxreg_file_219_port, B2 => n6125, ZN => 
                           n6016);
   U7793 : NAND3_X1 port map( A1 => n6018, A2 => n6017, A3 => n6016, ZN => 
                           n6019);
   U7794 : AOI21_X1 port map( B1 => IF_Regsxreg_file_155_port, B2 => n6164, A 
                           => n6019, ZN => n6036);
   U7795 : AOI22_X1 port map( A1 => IF_Regsxreg_file_315_port, A2 => n6098, B1 
                           => IF_Regsxreg_file_827_port, B2 => n6137, ZN => 
                           n6023);
   U7796 : AOI22_X1 port map( A1 => IF_Regsxreg_file_443_port, A2 => n6099, B1 
                           => IF_Regsxreg_file_955_port, B2 => n6138, ZN => 
                           n6022);
   U7797 : AOI22_X1 port map( A1 => IF_Regsxreg_file_699_port, A2 => n6041, B1 
                           => IF_Regsxreg_file_187_port, B2 => n6097, ZN => 
                           n6021);
   U7798 : AOI22_X1 port map( A1 => IF_Regsxreg_file_571_port, A2 => n6096, B1 
                           => IF_Regsxreg_file_59_port, B2 => n6068, ZN => 
                           n6020);
   U7799 : NAND4_X1 port map( A1 => n6023, A2 => n6022, A3 => n6021, A4 => 
                           n6020, ZN => n6034);
   U7800 : AOI22_X1 port map( A1 => IF_Regsxreg_file_347_port, A2 => n6104, B1 
                           => IF_Regsxreg_file_987_port, B2 => n6073, ZN => 
                           n6027);
   U7801 : AOI22_X1 port map( A1 => IF_Regsxreg_file_859_port, A2 => n6148, B1 
                           => IF_Regsxreg_file_475_port, B2 => n6106, ZN => 
                           n6026);
   U7802 : AOI22_X1 port map( A1 => IF_Regsxreg_file_123_port, A2 => n6114, B1 
                           => IF_Regsxreg_file_379_port, B2 => n6130, ZN => 
                           n6025);
   U7803 : AOI22_X1 port map( A1 => IF_Regsxreg_file_731_port, A2 => n6109, B1 
                           => IF_Regsxreg_file_91_port, B2 => n6149, ZN => 
                           n6024);
   U7804 : NAND4_X1 port map( A1 => n6027, A2 => n6026, A3 => n6025, A4 => 
                           n6024, ZN => n6033);
   U7805 : AOI22_X1 port map( A1 => IF_Regsxreg_file_763_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_795_port, B2 => n6051, ZN => 
                           n6031);
   U7806 : AOI22_X1 port map( A1 => IF_Regsxreg_file_27_port, A2 => n6165, B1 
                           => IF_Regsxreg_file_539_port, B2 => n6162, ZN => 
                           n6030);
   U7807 : AOI22_X1 port map( A1 => IF_Regsxreg_file_667_port, A2 => n6166, B1 
                           => IF_Regsxreg_file_923_port, B2 => n6167, ZN => 
                           n6029);
   U7808 : AOI22_X1 port map( A1 => IF_Regsxreg_file_283_port, A2 => n6160, B1 
                           => IF_Regsxreg_file_411_port, B2 => n6163, ZN => 
                           n6028);
   U7809 : NAND4_X1 port map( A1 => n6031, A2 => n6030, A3 => n6029, A4 => 
                           n6028, ZN => n6032);
   U7810 : AOI211_X1 port map( C1 => n6267, C2 => n6034, A => n6033, B => n6032
                           , ZN => n6035);
   U7811 : AOI21_X1 port map( B1 => n6036, B2 => n6035, A => n6175, ZN => 
                           IF_RegsxN622);
   U7812 : AOI22_X1 port map( A1 => IF_Regsxreg_file_508_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_476_port, B2 => n6106, ZN => 
                           n6039);
   U7813 : AOI22_X1 port map( A1 => IF_Regsxreg_file_732_port, A2 => n6127, B1 
                           => IF_Regsxreg_file_636_port, B2 => n6153, ZN => 
                           n6038);
   U7814 : AOI22_X1 port map( A1 => IF_Regsxreg_file_348_port, A2 => n6161, B1 
                           => IF_Regsxreg_file_124_port, B2 => n6114, ZN => 
                           n6037);
   U7815 : NAND3_X1 port map( A1 => n6039, A2 => n6038, A3 => n6037, ZN => 
                           n6040);
   U7816 : AOI21_X1 port map( B1 => IF_Regsxreg_file_412_port, B2 => n6163, A 
                           => n6040, ZN => n6061);
   U7817 : AOI22_X1 port map( A1 => IF_Regsxreg_file_572_port, A2 => n6143, B1 
                           => IF_Regsxreg_file_316_port, B2 => n6098, ZN => 
                           n6045);
   U7818 : AOI22_X1 port map( A1 => IF_Regsxreg_file_60_port, A2 => n6068, B1 
                           => IF_Regsxreg_file_444_port, B2 => n6099, ZN => 
                           n6044);
   U7819 : AOI22_X1 port map( A1 => IF_Regsxreg_file_956_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_828_port, B2 => n6137, ZN => 
                           n6043);
   U7820 : AOI22_X1 port map( A1 => IF_Regsxreg_file_700_port, A2 => n6041, B1 
                           => IF_Regsxreg_file_188_port, B2 => n6097, ZN => 
                           n6042);
   U7821 : NAND4_X1 port map( A1 => n6045, A2 => n6044, A3 => n6043, A4 => 
                           n6042, ZN => n6059);
   U7822 : AOI22_X1 port map( A1 => IF_Regsxreg_file_380_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_604_port, B2 => n6074, ZN => 
                           n6050);
   U7823 : AOI22_X1 port map( A1 => IF_Regsxreg_file_988_port, A2 => n6073, B1 
                           => IF_Regsxreg_file_860_port, B2 => n6148, ZN => 
                           n6049);
   U7824 : AOI22_X1 port map( A1 => IF_Regsxreg_file_764_port, A2 => n6150, B1 
                           => IF_Regsxreg_file_92_port, B2 => n6149, ZN => 
                           n6048);
   U7825 : AOI22_X1 port map( A1 => IF_Regsxreg_file_252_port, A2 => n6046, B1 
                           => IF_Regsxreg_file_892_port, B2 => n6128, ZN => 
                           n6047);
   U7826 : NAND4_X1 port map( A1 => n6050, A2 => n6049, A3 => n6048, A4 => 
                           n6047, ZN => n6058);
   U7827 : AOI22_X1 port map( A1 => IF_Regsxreg_file_220_port, A2 => n6125, B1 
                           => IF_Regsxreg_file_796_port, B2 => n6051, ZN => 
                           n6056);
   U7828 : AOI22_X1 port map( A1 => IF_Regsxreg_file_668_port, A2 => n6166, B1 
                           => IF_Regsxreg_file_28_port, B2 => n6052, ZN => 
                           n6055);
   U7829 : AOI22_X1 port map( A1 => IF_Regsxreg_file_540_port, A2 => n6080, B1 
                           => IF_Regsxreg_file_156_port, B2 => n6164, ZN => 
                           n6054);
   U7830 : AOI22_X1 port map( A1 => IF_Regsxreg_file_924_port, A2 => n6167, B1 
                           => IF_Regsxreg_file_284_port, B2 => n6160, ZN => 
                           n6053);
   U7831 : NAND4_X1 port map( A1 => n6056, A2 => n6055, A3 => n6054, A4 => 
                           n6053, ZN => n6057);
   U7832 : AOI211_X1 port map( C1 => n6267, C2 => n6059, A => n6058, B => n6057
                           , ZN => n6060);
   U7833 : AOI21_X1 port map( B1 => n6061, B2 => n6060, A => n6175, ZN => 
                           IF_RegsxN623);
   U7834 : AOI22_X1 port map( A1 => IF_Regsxreg_file_509_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_93_port, B2 => n6062, ZN => 
                           n6065);
   U7835 : AOI22_X1 port map( A1 => IF_Regsxreg_file_893_port, A2 => n6128, B1 
                           => IF_Regsxreg_file_125_port, B2 => n6114, ZN => 
                           n6064);
   U7836 : AOI22_X1 port map( A1 => IF_Regsxreg_file_637_port, A2 => n6153, B1 
                           => IF_Regsxreg_file_733_port, B2 => n6127, ZN => 
                           n6063);
   U7837 : NAND3_X1 port map( A1 => n6065, A2 => n6064, A3 => n6063, ZN => 
                           n6066);
   U7838 : AOI21_X1 port map( B1 => IF_Regsxreg_file_157_port, B2 => n6115, A 
                           => n6066, ZN => n6089);
   U7839 : AOI22_X1 port map( A1 => IF_Regsxreg_file_701_port, A2 => n6140, B1 
                           => IF_Regsxreg_file_317_port, B2 => n6098, ZN => 
                           n6072);
   U7840 : AOI22_X1 port map( A1 => IF_Regsxreg_file_957_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_189_port, B2 => n6097, ZN => 
                           n6071);
   U7841 : AOI22_X1 port map( A1 => IF_Regsxreg_file_829_port, A2 => n6067, B1 
                           => IF_Regsxreg_file_573_port, B2 => n6096, ZN => 
                           n6070);
   U7842 : AOI22_X1 port map( A1 => IF_Regsxreg_file_61_port, A2 => n6068, B1 
                           => IF_Regsxreg_file_445_port, B2 => n6099, ZN => 
                           n6069);
   U7843 : NAND4_X1 port map( A1 => n6072, A2 => n6071, A3 => n6070, A4 => 
                           n6069, ZN => n6087);
   U7844 : AOI22_X1 port map( A1 => IF_Regsxreg_file_861_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_221_port, B2 => n6125, ZN => 
                           n6078);
   U7845 : AOI22_X1 port map( A1 => IF_Regsxreg_file_253_port, A2 => n6152, B1 
                           => IF_Regsxreg_file_349_port, B2 => n6104, ZN => 
                           n6077);
   U7846 : AOI22_X1 port map( A1 => IF_Regsxreg_file_605_port, A2 => n6074, B1 
                           => IF_Regsxreg_file_989_port, B2 => n6073, ZN => 
                           n6076);
   U7847 : AOI22_X1 port map( A1 => IF_Regsxreg_file_765_port, A2 => n6150, B1 
                           => IF_Regsxreg_file_477_port, B2 => n6106, ZN => 
                           n6075);
   U7848 : NAND4_X1 port map( A1 => n6078, A2 => n6077, A3 => n6076, A4 => 
                           n6075, ZN => n6086);
   U7849 : AOI22_X1 port map( A1 => IF_Regsxreg_file_381_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_669_port, B2 => n6166, ZN => 
                           n6084);
   U7850 : AOI22_X1 port map( A1 => IF_Regsxreg_file_29_port, A2 => n6165, B1 
                           => IF_Regsxreg_file_925_port, B2 => n6167, ZN => 
                           n6083);
   U7851 : AOI22_X1 port map( A1 => IF_Regsxreg_file_797_port, A2 => n6135, B1 
                           => IF_Regsxreg_file_413_port, B2 => n6079, ZN => 
                           n6082);
   U7852 : AOI22_X1 port map( A1 => IF_Regsxreg_file_541_port, A2 => n6080, B1 
                           => IF_Regsxreg_file_285_port, B2 => n6160, ZN => 
                           n6081);
   U7853 : NAND4_X1 port map( A1 => n6084, A2 => n6083, A3 => n6082, A4 => 
                           n6081, ZN => n6085);
   U7854 : AOI211_X1 port map( C1 => n6267, C2 => n6087, A => n6086, B => n6085
                           , ZN => n6088);
   U7855 : AOI21_X1 port map( B1 => n6089, B2 => n6088, A => n6175, ZN => 
                           IF_RegsxN624);
   U7856 : AOI22_X1 port map( A1 => IF_Regsxreg_file_510_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_222_port, B2 => n6125, ZN => 
                           n6094);
   U7857 : AOI22_X1 port map( A1 => IF_Regsxreg_file_766_port, A2 => n6091, B1 
                           => IF_Regsxreg_file_990_port, B2 => n6090, ZN => 
                           n6093);
   U7858 : AOI22_X1 port map( A1 => IF_Regsxreg_file_94_port, A2 => n6149, B1 
                           => IF_Regsxreg_file_254_port, B2 => n6152, ZN => 
                           n6092);
   U7859 : NAND3_X1 port map( A1 => n6094, A2 => n6093, A3 => n6092, ZN => 
                           n6095);
   U7860 : AOI21_X1 port map( B1 => IF_Regsxreg_file_414_port, B2 => n6163, A 
                           => n6095, ZN => n6124);
   U7861 : AOI22_X1 port map( A1 => IF_Regsxreg_file_830_port, A2 => n6137, B1 
                           => IF_Regsxreg_file_702_port, B2 => n6140, ZN => 
                           n6103);
   U7862 : AOI22_X1 port map( A1 => IF_Regsxreg_file_958_port, A2 => n6138, B1 
                           => IF_Regsxreg_file_62_port, B2 => n6142, ZN => 
                           n6102);
   U7863 : AOI22_X1 port map( A1 => IF_Regsxreg_file_190_port, A2 => n6097, B1 
                           => IF_Regsxreg_file_574_port, B2 => n6096, ZN => 
                           n6101);
   U7864 : AOI22_X1 port map( A1 => IF_Regsxreg_file_446_port, A2 => n6099, B1 
                           => IF_Regsxreg_file_318_port, B2 => n6098, ZN => 
                           n6100);
   U7865 : NAND4_X1 port map( A1 => n6103, A2 => n6102, A3 => n6101, A4 => 
                           n6100, ZN => n6122);
   U7866 : AOI22_X1 port map( A1 => IF_Regsxreg_file_862_port, A2 => n6105, B1 
                           => IF_Regsxreg_file_350_port, B2 => n6104, ZN => 
                           n6113);
   U7867 : AOI22_X1 port map( A1 => IF_Regsxreg_file_894_port, A2 => n6107, B1 
                           => IF_Regsxreg_file_478_port, B2 => n6106, ZN => 
                           n6112);
   U7868 : AOI22_X1 port map( A1 => IF_Regsxreg_file_382_port, A2 => n6108, B1 
                           => IF_Regsxreg_file_606_port, B2 => n6151, ZN => 
                           n6111);
   U7869 : AOI22_X1 port map( A1 => IF_Regsxreg_file_734_port, A2 => n6109, B1 
                           => IF_Regsxreg_file_638_port, B2 => n6153, ZN => 
                           n6110);
   U7870 : NAND4_X1 port map( A1 => n6113, A2 => n6112, A3 => n6111, A4 => 
                           n6110, ZN => n6121);
   U7871 : AOI22_X1 port map( A1 => IF_Regsxreg_file_926_port, A2 => n6167, B1 
                           => IF_Regsxreg_file_126_port, B2 => n6114, ZN => 
                           n6119);
   U7872 : AOI22_X1 port map( A1 => IF_Regsxreg_file_30_port, A2 => n6165, B1 
                           => IF_Regsxreg_file_286_port, B2 => n6160, ZN => 
                           n6118);
   U7873 : AOI22_X1 port map( A1 => IF_Regsxreg_file_798_port, A2 => n6135, B1 
                           => IF_Regsxreg_file_542_port, B2 => n6162, ZN => 
                           n6117);
   U7874 : AOI22_X1 port map( A1 => IF_Regsxreg_file_158_port, A2 => n6115, B1 
                           => IF_Regsxreg_file_670_port, B2 => n6166, ZN => 
                           n6116);
   U7875 : NAND4_X1 port map( A1 => n6119, A2 => n6118, A3 => n6117, A4 => 
                           n6116, ZN => n6120);
   U7876 : AOI211_X1 port map( C1 => n6267, C2 => n6122, A => n6121, B => n6120
                           , ZN => n6123);
   U7877 : AOI21_X1 port map( B1 => n6124, B2 => n6123, A => n6175, ZN => 
                           IF_RegsxN625);
   U7878 : AOI22_X1 port map( A1 => IF_Regsxreg_file_511_port, A2 => n6126, B1 
                           => IF_Regsxreg_file_223_port, B2 => n6125, ZN => 
                           n6133);
   U7879 : AOI22_X1 port map( A1 => IF_Regsxreg_file_895_port, A2 => n6128, B1 
                           => IF_Regsxreg_file_735_port, B2 => n6127, ZN => 
                           n6132);
   U7880 : AOI22_X1 port map( A1 => IF_Regsxreg_file_383_port, A2 => n6130, B1 
                           => IF_Regsxreg_file_127_port, B2 => n6129, ZN => 
                           n6131);
   U7881 : NAND3_X1 port map( A1 => n6133, A2 => n6132, A3 => n6131, ZN => 
                           n6134);
   U7882 : AOI21_X1 port map( B1 => IF_Regsxreg_file_799_port, B2 => n6135, A 
                           => n6134, ZN => n6177);
   U7883 : AOI22_X1 port map( A1 => IF_Regsxreg_file_831_port, A2 => n6137, B1 
                           => IF_Regsxreg_file_447_port, B2 => n6136, ZN => 
                           n6147);
   U7884 : AOI22_X1 port map( A1 => IF_Regsxreg_file_191_port, A2 => n6139, B1 
                           => IF_Regsxreg_file_959_port, B2 => n6138, ZN => 
                           n6146);
   U7885 : AOI22_X1 port map( A1 => IF_Regsxreg_file_319_port, A2 => n6141, B1 
                           => IF_Regsxreg_file_703_port, B2 => n6140, ZN => 
                           n6145);
   U7886 : AOI22_X1 port map( A1 => IF_Regsxreg_file_575_port, A2 => n6143, B1 
                           => IF_Regsxreg_file_63_port, B2 => n6142, ZN => 
                           n6144);
   U7887 : NAND4_X1 port map( A1 => n6147, A2 => n6146, A3 => n6145, A4 => 
                           n6144, ZN => n6174);
   U7888 : AOI22_X1 port map( A1 => IF_Regsxreg_file_95_port, A2 => n6149, B1 
                           => IF_Regsxreg_file_863_port, B2 => n6148, ZN => 
                           n6159);
   U7889 : AOI22_X1 port map( A1 => IF_Regsxreg_file_607_port, A2 => n6151, B1 
                           => IF_Regsxreg_file_767_port, B2 => n6150, ZN => 
                           n6158);
   U7890 : AOI22_X1 port map( A1 => IF_Regsxreg_file_639_port, A2 => n6153, B1 
                           => IF_Regsxreg_file_255_port, B2 => n6152, ZN => 
                           n6157);
   U7891 : AOI22_X1 port map( A1 => IF_Regsxreg_file_479_port, A2 => n6155, B1 
                           => IF_Regsxreg_file_991_port, B2 => n6154, ZN => 
                           n6156);
   U7892 : NAND4_X1 port map( A1 => n6159, A2 => n6158, A3 => n6157, A4 => 
                           n6156, ZN => n6173);
   U7893 : AOI22_X1 port map( A1 => IF_Regsxreg_file_351_port, A2 => n6161, B1 
                           => IF_Regsxreg_file_287_port, B2 => n6160, ZN => 
                           n6171);
   U7894 : AOI22_X1 port map( A1 => IF_Regsxreg_file_415_port, A2 => n6163, B1 
                           => IF_Regsxreg_file_543_port, B2 => n6162, ZN => 
                           n6170);
   U7895 : AOI22_X1 port map( A1 => IF_Regsxreg_file_31_port, A2 => n6165, B1 
                           => IF_Regsxreg_file_159_port, B2 => n6164, ZN => 
                           n6169);
   U7896 : AOI22_X1 port map( A1 => IF_Regsxreg_file_927_port, A2 => n6167, B1 
                           => IF_Regsxreg_file_671_port, B2 => n6166, ZN => 
                           n6168);
   U7897 : NAND4_X1 port map( A1 => n6171, A2 => n6170, A3 => n6169, A4 => 
                           n6168, ZN => n6172);
   U7898 : AOI211_X1 port map( C1 => n6267, C2 => n6174, A => n6173, B => n6172
                           , ZN => n6176);
   U7899 : AOI21_X1 port map( B1 => n6177, B2 => n6176, A => n6175, ZN => 
                           IF_RegsxN626);
   U7900 : OAI21_X1 port map( B1 => CtlToRegs_port_req, B2 => n6237, A => n6178
                           , ZN => IF_RegsxN594);
   U7901 : INV_X1 port map( A => n6179, ZN => n6181);
   U7902 : OAI211_X1 port map( C1 => n6182, C2 => n6181, A => 
                           CtlToDec_port_notify, B => n6180, ZN => n6183);
   U7903 : OAI21_X1 port map( B1 => n6185, B2 => n6184, A => n6183, ZN => n2946
                           );
   U7904 : AOI21_X1 port map( B1 => MemToCtl_port_notify_port, B2 => n6187, A 
                           => n6186, ZN => n6188);
   U7905 : NOR2_X1 port map( A1 => rst, A2 => n6188, ZN => n2944);
   clk_gate_IF_ALUxALUtoCtl_port_reg : SNPS_CLOCK_GATE_HIGH_CPU_0 port map( CLK
                           => clk, EN => IF_ALUxN937, ENCLK => net2468144);
   clk_gate_IF_CPathxCtlToALU_port_op2_sel_reg : SNPS_CLOCK_GATE_HIGH_CPU_54 
                           port map( CLK => clk, EN => IF_CPathxN2396, ENCLK =>
                           net2468149);
   clk_gate_IF_CPathxCtlToRegs_port_src2_reg : SNPS_CLOCK_GATE_HIGH_CPU_53 port
                           map( CLK => clk, EN => IF_CPathxN2394, ENCLK => 
                           net2468154);
   clk_gate_IF_CPathxCtlToDec_port_reg : SNPS_CLOCK_GATE_HIGH_CPU_52 port map( 
                           CLK => clk, EN => IF_CPathxN2393, ENCLK => 
                           net2468159);
   clk_gate_IF_CPathxCtlToMem_port_req_reg : SNPS_CLOCK_GATE_HIGH_CPU_51 port 
                           map( CLK => clk, EN => IF_CPathxN2316, ENCLK => 
                           net2468164);
   clk_gate_IF_CPathxwb_sel_signal_reg : SNPS_CLOCK_GATE_HIGH_CPU_50 port map( 
                           CLK => clk, EN => IF_CPathxN2310, ENCLK => 
                           net2468169);
   clk_gate_IF_CPathxpc_reg_signal_reg : SNPS_CLOCK_GATE_HIGH_CPU_49 port map( 
                           CLK => clk, EN => IF_CPathxN2274, ENCLK => 
                           net2468174);
   clk_gate_IF_CPathxpc_next_signal_reg : SNPS_CLOCK_GATE_HIGH_CPU_48 port map(
                           CLK => clk, EN => IF_CPathxN1859, ENCLK => 
                           net2468179);
   clk_gate_IF_CPathxmemoryAccess_signal_mask_reg : SNPS_CLOCK_GATE_HIGH_CPU_47
                           port map( CLK => clk, EN => IF_CPathxN2235, ENCLK =>
                           net2468184);
   clk_gate_IF_CPathxMemToCtl_data_signal_reg : SNPS_CLOCK_GATE_HIGH_CPU_46 
                           port map( CLK => clk, EN => IF_CPathxN2201, ENCLK =>
                           net2468189);
   clk_gate_IF_CPathxDecToCtl_data_signal_rd_addr_reg : 
                           SNPS_CLOCK_GATE_HIGH_CPU_45 port map( CLK => clk, EN
                           => IF_CPathxN2157, ENCLK => net2468194);
   clk_gate_IF_CPathxRegsToCtl_data_signal_contents2_reg : 
                           SNPS_CLOCK_GATE_HIGH_CPU_44 port map( CLK => clk, EN
                           => IF_CPathxN2091, ENCLK => net2468199);
   clk_gate_IF_CPathxCtlToRegs_data_signal_src2_reg : 
                           SNPS_CLOCK_GATE_HIGH_CPU_43 port map( CLK => clk, EN
                           => IF_CPathxN2078, ENCLK => net2468204);
   clk_gate_IF_CPathxCtlToRegs_port_req_reg : SNPS_CLOCK_GATE_HIGH_CPU_42 port 
                           map( CLK => clk, EN => IF_CPathxN2038, ENCLK => 
                           net2468209);
   clk_gate_IF_CPathxCtlToRegs_port_dst_data_reg : SNPS_CLOCK_GATE_HIGH_CPU_41 
                           port map( CLK => clk, EN => IF_CPathxN2044, ENCLK =>
                           net2468214);
   clk_gate_IF_CPathxCtlToRegs_data_signal_dst_reg : 
                           SNPS_CLOCK_GATE_HIGH_CPU_40 port map( CLK => clk, EN
                           => IF_CPathxN2032, ENCLK => net2468219);
   clk_gate_IF_CPathxCtlToALU_port_reg2_contents_reg : 
                           SNPS_CLOCK_GATE_HIGH_CPU_39 port map( CLK => clk, EN
                           => IF_CPathxN1935, ENCLK => net2468224);
   clk_gate_IF_CPathxCtlToALU_data_signal_op2_sel_reg : 
                           SNPS_CLOCK_GATE_HIGH_CPU_38 port map( CLK => clk, EN
                           => IF_CPathxN1930, ENCLK => net2468229);
   clk_gate_IF_CPathxCtlToALU_data_signal_alu_fun_reg : 
                           SNPS_CLOCK_GATE_HIGH_CPU_37 port map( CLK => clk, EN
                           => IF_CPathxN1892, ENCLK => net2468234);
   clk_gate_IF_CPathxsection_reg : SNPS_CLOCK_GATE_HIGH_CPU_36 port map( CLK =>
                           clk, EN => IF_CPathxN1854, ENCLK => net2468239);
   clk_gate_IF_DecoderxDecToCtl_port_rs2_addr_reg : SNPS_CLOCK_GATE_HIGH_CPU_34
                           port map( CLK => clk, EN => IF_DecoderxN596, ENCLK 
                           => net2468249);
   clk_gate_IF_DecoderxDecToCtl_port_imm_reg : SNPS_CLOCK_GATE_HIGH_CPU_33 port
                           map( CLK => clk, EN => IF_DecoderxN552, ENCLK => 
                           net2468254);
   clk_gate_IF_Regsxreg_file_regx31x : SNPS_CLOCK_GATE_HIGH_CPU_32 port map( 
                           CLK => clk, EN => IF_RegsxN659, ENCLK => net2468259)
                           ;
   clk_gate_IF_Regsxreg_file_regx30x : SNPS_CLOCK_GATE_HIGH_CPU_31 port map( 
                           CLK => clk, EN => IF_RegsxN692, ENCLK => net2468264)
                           ;
   clk_gate_IF_Regsxreg_file_regx29x : SNPS_CLOCK_GATE_HIGH_CPU_30 port map( 
                           CLK => clk, EN => IF_RegsxN693, ENCLK => net2468269)
                           ;
   clk_gate_IF_Regsxreg_file_regx28x : SNPS_CLOCK_GATE_HIGH_CPU_29 port map( 
                           CLK => clk, EN => IF_RegsxN694, ENCLK => net2468274)
                           ;
   clk_gate_IF_Regsxreg_file_regx27x : SNPS_CLOCK_GATE_HIGH_CPU_28 port map( 
                           CLK => clk, EN => IF_RegsxN695, ENCLK => net2468279)
                           ;
   clk_gate_IF_Regsxreg_file_regx26x : SNPS_CLOCK_GATE_HIGH_CPU_27 port map( 
                           CLK => clk, EN => IF_RegsxN696, ENCLK => net2468284)
                           ;
   clk_gate_IF_Regsxreg_file_regx25x : SNPS_CLOCK_GATE_HIGH_CPU_26 port map( 
                           CLK => clk, EN => IF_RegsxN697, ENCLK => net2468289)
                           ;
   clk_gate_IF_Regsxreg_file_regx24x : SNPS_CLOCK_GATE_HIGH_CPU_25 port map( 
                           CLK => clk, EN => IF_RegsxN698, ENCLK => net2468294)
                           ;
   clk_gate_IF_Regsxreg_file_regx23x : SNPS_CLOCK_GATE_HIGH_CPU_24 port map( 
                           CLK => clk, EN => IF_RegsxN699, ENCLK => net2468299)
                           ;
   clk_gate_IF_Regsxreg_file_regx22x : SNPS_CLOCK_GATE_HIGH_CPU_23 port map( 
                           CLK => clk, EN => IF_RegsxN700, ENCLK => net2468304)
                           ;
   clk_gate_IF_Regsxreg_file_regx21x : SNPS_CLOCK_GATE_HIGH_CPU_22 port map( 
                           CLK => clk, EN => IF_RegsxN701, ENCLK => net2468309)
                           ;
   clk_gate_IF_Regsxreg_file_regx20x : SNPS_CLOCK_GATE_HIGH_CPU_21 port map( 
                           CLK => clk, EN => IF_RegsxN702, ENCLK => net2468314)
                           ;
   clk_gate_IF_Regsxreg_file_regx19x : SNPS_CLOCK_GATE_HIGH_CPU_20 port map( 
                           CLK => clk, EN => IF_RegsxN703, ENCLK => net2468319)
                           ;
   clk_gate_IF_Regsxreg_file_regx18x : SNPS_CLOCK_GATE_HIGH_CPU_19 port map( 
                           CLK => clk, EN => IF_RegsxN704, ENCLK => net2468324)
                           ;
   clk_gate_IF_Regsxreg_file_regx17x : SNPS_CLOCK_GATE_HIGH_CPU_18 port map( 
                           CLK => clk, EN => IF_RegsxN705, ENCLK => net2468329)
                           ;
   clk_gate_IF_Regsxreg_file_regx16x : SNPS_CLOCK_GATE_HIGH_CPU_17 port map( 
                           CLK => clk, EN => IF_RegsxN706, ENCLK => net2468334)
                           ;
   clk_gate_IF_Regsxreg_file_regx15x : SNPS_CLOCK_GATE_HIGH_CPU_16 port map( 
                           CLK => clk, EN => IF_RegsxN707, ENCLK => net2468339)
                           ;
   clk_gate_IF_Regsxreg_file_regx14x : SNPS_CLOCK_GATE_HIGH_CPU_15 port map( 
                           CLK => clk, EN => IF_RegsxN708, ENCLK => net2468344)
                           ;
   clk_gate_IF_Regsxreg_file_regx13x : SNPS_CLOCK_GATE_HIGH_CPU_14 port map( 
                           CLK => clk, EN => IF_RegsxN709, ENCLK => net2468349)
                           ;
   clk_gate_IF_Regsxreg_file_regx12x : SNPS_CLOCK_GATE_HIGH_CPU_13 port map( 
                           CLK => clk, EN => IF_RegsxN710, ENCLK => net2468354)
                           ;
   clk_gate_IF_Regsxreg_file_regx11x : SNPS_CLOCK_GATE_HIGH_CPU_12 port map( 
                           CLK => clk, EN => IF_RegsxN711, ENCLK => net2468359)
                           ;
   clk_gate_IF_Regsxreg_file_regx10x : SNPS_CLOCK_GATE_HIGH_CPU_11 port map( 
                           CLK => clk, EN => IF_RegsxN712, ENCLK => net2468364)
                           ;
   clk_gate_IF_Regsxreg_file_regx9x : SNPS_CLOCK_GATE_HIGH_CPU_10 port map( CLK
                           => clk, EN => IF_RegsxN713, ENCLK => net2468369);
   clk_gate_IF_Regsxreg_file_regx8x : SNPS_CLOCK_GATE_HIGH_CPU_9 port map( CLK 
                           => clk, EN => IF_RegsxN714, ENCLK => net2468374);
   clk_gate_IF_Regsxreg_file_regx7x : SNPS_CLOCK_GATE_HIGH_CPU_8 port map( CLK 
                           => clk, EN => IF_RegsxN715, ENCLK => net2468379);
   clk_gate_IF_Regsxreg_file_regx6x : SNPS_CLOCK_GATE_HIGH_CPU_7 port map( CLK 
                           => clk, EN => IF_RegsxN716, ENCLK => net2468384);
   clk_gate_IF_Regsxreg_file_regx5x : SNPS_CLOCK_GATE_HIGH_CPU_6 port map( CLK 
                           => clk, EN => IF_RegsxN717, ENCLK => net2468389);
   clk_gate_IF_Regsxreg_file_regx4x : SNPS_CLOCK_GATE_HIGH_CPU_5 port map( CLK 
                           => clk, EN => IF_RegsxN718, ENCLK => net2468394);
   clk_gate_IF_Regsxreg_file_regx3x : SNPS_CLOCK_GATE_HIGH_CPU_4 port map( CLK 
                           => clk, EN => IF_RegsxN719, ENCLK => net2468399);
   clk_gate_IF_Regsxreg_file_regx2x : SNPS_CLOCK_GATE_HIGH_CPU_3 port map( CLK 
                           => clk, EN => IF_RegsxN720, ENCLK => net2468404);
   clk_gate_IF_Regsxreg_file_regx1x : SNPS_CLOCK_GATE_HIGH_CPU_2 port map( CLK 
                           => clk, EN => IF_RegsxN721, ENCLK => net2468409);
   clk_gate_IF_RegsxRegsToCtl_port_contents2_reg : SNPS_CLOCK_GATE_HIGH_CPU_1 
                           port map( CLK => clk, EN => IF_RegsxN594, ENCLK => 
                           net2468414);

end SYN_CPU_arch;
