library ieee;
use IEEE.numeric_std.all;

package TestBasic10_types is
type TestBasic10_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic10_types;
