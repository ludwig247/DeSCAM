library ieee;
use IEEE.numeric_std.all;

package TestBasic4_types is
type TestBasic4_SECTIONS is (run);
end package TestBasic4_types;
