library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave4_types is
type TestMasterSlave4_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave4_types;
