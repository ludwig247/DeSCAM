library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave12_types is
type TestMasterSlave12_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave12_types;
