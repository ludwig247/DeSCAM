package testbasic9_types;

	typedef enum logic {
		run
	} TestBasic9_SECTIONS;

endpackage
