library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestMasterSlave4_types is
type Sections is (SECTION_A, SECTION_B);
end package TestMasterSlave4_types;