library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestGlobal2_types is
-- No local datatypes implemented!


end package TestGlobal2_types;