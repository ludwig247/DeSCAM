library ieee;
use IEEE.numeric_std.all;

package TestBasic5_types is
end package TestBasic5_types;