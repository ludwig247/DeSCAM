library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestArray4_types is
end package TestArray4_types;