library ieee;
use IEEE.numeric_std.all;

package TestBasic20_types is
type TestBasic20_SECTIONS is (SECTION_A, SECTION_B);
type color_t is (GREEN, RED, YELLOW);
end package TestBasic20_types;
