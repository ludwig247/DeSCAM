package testbasic10_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic10_SECTIONS;

endpackage
