package testmasterslave2_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave2_SECTIONS;

endpackage
