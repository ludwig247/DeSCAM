package testbasic8_types;

	typedef enum logic {
		run
	} TestBasic8_SECTIONS;

endpackage
