library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave6_types is
type TestMasterSlave6_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave6_types;

