package testmasterslave4_types;

	import scam_model_types::*;
	typedef enum logic {
		section_a,
		section_b
	} Sections;

endpackage