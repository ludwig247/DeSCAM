library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestMasterSlave18_types is
-- No local datatypes implemented!


end package TestMasterSlave18_types;