package testarray2_types;

	import scam_model_types::*;
endpackage