library ieee;
use IEEE.numeric_std.all;

package TestBasic21_types is
type TestBasic21_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic21_types;
