library ieee;
use IEEE.numeric_std.all;

package TestBasic13_types is
type TestBasic13_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic13_types;
