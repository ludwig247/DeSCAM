library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestFunction2_types is
end package TestFunction2_types;