package testbasic4_types;

	import scam_model_types::*;
endpackage