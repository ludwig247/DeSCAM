package testarray0_types;

	 import top_level_types::*;
endpackage