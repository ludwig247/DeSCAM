package SCAM_Model_types is
subtype bool is Boolean;
subtype int is Integer;
type ALUfuncType is (ALU_ADD,ALU_AND,ALU_COPY1,ALU_OR,ALU_SLL,ALU_SLT,ALU_SLTU,ALU_SRA,ALU_SRL,ALU_SUB,ALU_X,ALU_XOR);
type AmoInstrType is (AMO_ADD,AMO_AND,AMO_LR,AMO_MAX,AMO_MAXU,AMO_MIN,AMO_MINU,AMO_OR,AMO_SC,AMO_SWAP,AMO_UNKNOWN,AMO_XOR);
type EncType is (ENC_A,ENC_B,ENC_ERR,ENC_I_I,ENC_I_J,ENC_I_L,ENC_I_M,ENC_I_S,ENC_J,ENC_R,ENC_S,ENC_U);
type ISA_SECTIONS is (execute,fetch);
type InstrType_Complete is (INSTR_ADD,INSTR_ADDI,INSTR_AND,INSTR_ANDI,INSTR_AUIPC,INSTR_BEQ,INSTR_BGE,INSTR_BGEU,INSTR_BLT,INSTR_BLTU,INSTR_BNE,INSTR_CSRRC,INSTR_CSRRCI,INSTR_CSRRS,INSTR_CSRRSI,INSTR_CSRRW,INSTR_CSRRWI,INSTR_FENCE,INSTR_FENCEI,INSTR_JAL,INSTR_JALR,INSTR_LB,INSTR_LBU,INSTR_LH,INSTR_LHU,INSTR_LUI,INSTR_LW,INSTR_OR,INSTR_ORI,INSTR_PRIV,INSTR_SB,INSTR_SH,INSTR_SLL,INSTR_SLLI,INSTR_SLT,INSTR_SLTI,INSTR_SLTU,INSTR_SLTUI,INSTR_SRA,INSTR_SRAI,INSTR_SRL,INSTR_SRLI,INSTR_SUB,INSTR_SW,INSTR_UNKNOWN,INSTR_XOR,INSTR_XORI);
type LR_SC is (LR,NONE,SC);
type ME_AccessType is (ME_RD,ME_WR,ME_X);
type ME_MaskType is (MT_B,MT_BU,MT_H,MT_HU,MT_W,MT_X);
type MMUaccessType is (FETCH,LOAD,STORE);
type PrivInstrType is (INSTR_EBREAK,INSTR_ECALL,INSTR_MRET,INSTR_PRIV_UNKNOWN,INSTR_SFENCEVMA,INSTR_SRET,INSTR_URET,INSTR_WFI);
type CSRfileType is record
	mcause: unsigned;
	mcounteren: unsigned;
	mcycleh: unsigned;
	mcyclel: unsigned;
	medeleg: unsigned;
	mepc: unsigned;
	mideleg: unsigned;
	mie: unsigned;
	minstreth: unsigned;
	minstretl: unsigned;
	mip: unsigned;
	misa: unsigned;
	mscratch: unsigned;
	mstatus: unsigned;
	mtimeh: unsigned;
	mtimel: unsigned;
	mtval: unsigned;
	mtvec: unsigned;
	satp: unsigned;
	scause: unsigned;
	scounteren: unsigned;
	sedeleg: unsigned;
	sepc: unsigned;
	sideleg: unsigned;
	sscratch: unsigned;
	stval: unsigned;
	stvec: unsigned;
	ucause: unsigned;
	uepc: unsigned;
	uscratch: unsigned;
	utval: unsigned;
	utvec: unsigned;
end record;
type CUtoME_IF is record
	addrIn: unsigned;
	dataIn: unsigned;
	mask: ME_MaskType;
	req: ME_AccessType;
end record;
type MEtoCU_IF is record
	loadedData: unsigned;
end record;
type MMU_in is record
	accesstype: MMUaccessType;
	data: unsigned;
	exception_in: unsigned;
	lrsc: LR_SC;
	mask: ME_MaskType;
	mstatus: unsigned;
	prv: unsigned;
	reset_lrsc: unsigned;
	satp: unsigned;
	v_addr: unsigned;
end record;
type MMU_return is record
	data: unsigned;
	exception: unsigned;
	sc_success: unsigned;
end record;
type RegfileType is record
	reg_file_01: unsigned;
	reg_file_02: unsigned;
	reg_file_03: unsigned;
	reg_file_04: unsigned;
	reg_file_05: unsigned;
	reg_file_06: unsigned;
	reg_file_07: unsigned;
	reg_file_08: unsigned;
	reg_file_09: unsigned;
	reg_file_10: unsigned;
	reg_file_11: unsigned;
	reg_file_12: unsigned;
	reg_file_13: unsigned;
	reg_file_14: unsigned;
	reg_file_15: unsigned;
	reg_file_16: unsigned;
	reg_file_17: unsigned;
	reg_file_18: unsigned;
	reg_file_19: unsigned;
	reg_file_20: unsigned;
	reg_file_21: unsigned;
	reg_file_22: unsigned;
	reg_file_23: unsigned;
	reg_file_24: unsigned;
	reg_file_25: unsigned;
	reg_file_26: unsigned;
	reg_file_27: unsigned;
	reg_file_28: unsigned;
	reg_file_29: unsigned;
	reg_file_30: unsigned;
	reg_file_31: unsigned;
end record;
type RegfileWriteType is record
	dst: unsigned;
	dstData: unsigned;
	exception: unsigned;
end record;
end package SCAM_Model_types;
