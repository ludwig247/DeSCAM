library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestArray5_types is
end package TestArray5_types;