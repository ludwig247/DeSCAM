library ieee;
use IEEE.numeric_std.all;
use work.SCAM_Model_types.all;

package TestBasic3_types is
end package TestBasic3_types;