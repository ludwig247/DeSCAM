package testfunction2_types;

	typedef enum logic {
		run
	} TestFunction2_SECTIONS;

endpackage
