library ieee ;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all; 
use work.SCAM_Model_types.all;

entity ISA is
port(	
	clk:		in std_logic;
	rst:		in std_logic;
	ecall_isa_Port:		in bool;
	ecall_isa_Port_sync:	 in bool;
	ecall_isa_Port_notify:	 out bool;
	fromMemoryPort:		in MMU_return;
	fromMemoryPort_sync:	 in bool;
	fromMemoryPort_notify:	 out bool;
	fromRegsPort:		in RegfileType;
	fromRegsPort_sync:	 in bool;
	fromRegsPort_notify:	 out bool;
	isa_ecall_Port:		out bool;
	isa_ecall_Port_sync:	 in bool;
	isa_ecall_Port_notify:	 out bool;
	mip_isa_Port:		in unsigned;
	mip_isa_Port_sync:	 in bool;
	mip_isa_Port_notify:	 out bool;
	toMemoryPort:		out MMU_in;
	toMemoryPort_sync:	 in bool;
	toMemoryPort_notify:	 out bool;
	toRegsPort:		out RegfileWriteType;
	toRegsPort_sync:	 in bool;
	toRegsPort_notify:	 out bool);
end ISA;

architecture ISA_arch of ISA is
signal section: ISA_SECTIONS;
			 signal aluOp1_signal:unsigned(31 down to 0);
			 signal aluOp2_signal:unsigned(31 down to 0);
			 signal aluResult_signal:unsigned(31 down to 0);
			 signal csrfile_signal:CSRfileType;
			 signal encodedInstr_signal:unsigned(31 down to 0);
			 signal exception_signal:unsigned(31 down to 0);
			 signal fromMemoryData_signal:MEtoCU_IF;
			 signal from_mmu_signal:MMU_return;
			 signal isaREQ_signal:bool;
			 signal lastPc_signal:unsigned(31 down to 0);
			 signal lr_sc_signal:unsigned(31 down to 0);
			 signal mip_tmp_signal:unsigned(31 down to 0);
			 signal pcReg_signal:unsigned(31 down to 0);
			 signal pending_signal:unsigned(31 down to 0);
			 signal prv_signal:unsigned(31 down to 0);
			 signal regfile_signal:RegfileType;
			 signal regfileWrite_signal:RegfileWriteType;
			 signal sysRES_signal:bool;
			 signal target_prv_signal:unsigned(31 down to 0);
			 signal toMemoryData_signal:CUtoME_IF;
			 signal to_mmu_signal:MMU_in;
			 signal write_signal:unsigned(31 down to 0);
			 signal xcause_signal:unsigned(31 down to 0);
			 signal xstatus_mask_signal:unsigned(31 down to 0);
			 signal xtval_signal:unsigned(31 down to 0);
			 signal xtvec_signal:unsigned(31 down to 0);
begin
	 process(clk)
	 begin
	 if(clk='1' and clk'event) then
		 if rst = '1' then
			 section <=fetch;
			aluOp1_signal:= (others => 0);
			aluOp2_signal:= (others => 0);
			aluResult_signal:= (others => 0);
			csrfile_signal.mcause<=0;
			csrfile_signal.mcounteren<=0;
			csrfile_signal.mcycleh<=0;
			csrfile_signal.mcyclel<=0;
			csrfile_signal.medeleg<=0;
			csrfile_signal.mepc<=0;
			csrfile_signal.mideleg<=0;
			csrfile_signal.mie<=0;
			csrfile_signal.minstreth<=0;
			csrfile_signal.minstretl<=0;
			csrfile_signal.mip<=0;
			csrfile_signal.misa<=0;
			csrfile_signal.mscratch<=0;
			csrfile_signal.mstatus<=0;
			csrfile_signal.mtimeh<=0;
			csrfile_signal.mtimel<=0;
			csrfile_signal.mtval<=0;
			csrfile_signal.mtvec<=0;
			csrfile_signal.satp<=0;
			csrfile_signal.scause<=0;
			csrfile_signal.scounteren<=0;
			csrfile_signal.sedeleg<=0;
			csrfile_signal.sepc<=0;
			csrfile_signal.sideleg<=0;
			csrfile_signal.sscratch<=0;
			csrfile_signal.stval<=0;
			csrfile_signal.stvec<=0;
			csrfile_signal.ucause<=0;
			csrfile_signal.uepc<=0;
			csrfile_signal.uscratch<=0;
			csrfile_signal.utval<=0;
			csrfile_signal.utvec<=0;
			encodedInstr_signal:= (others => 0);
			exception_signal:= (others => 0);
			fromMemoryData_signal.loadedData<=0;
			from_mmu_signal.data<=0;
			from_mmu_signal.exception<=0;
			from_mmu_signal.sc_success<=0;
			isaREQ_signal<=false;
			lastPc_signal:= (others => 0);
			lr_sc_signal:= (others => 0);
			mip_tmp_signal:= (others => 0);
			pcReg_signal:= (others => 0);
			pending_signal:= (others => 0);
			prv_signal:= (others => 3);
			regfile_signal.reg_file_01<=0;
			regfile_signal.reg_file_02<=0;
			regfile_signal.reg_file_03<=0;
			regfile_signal.reg_file_04<=0;
			regfile_signal.reg_file_05<=0;
			regfile_signal.reg_file_06<=0;
			regfile_signal.reg_file_07<=0;
			regfile_signal.reg_file_08<=0;
			regfile_signal.reg_file_09<=0;
			regfile_signal.reg_file_10<=0;
			regfile_signal.reg_file_11<=0;
			regfile_signal.reg_file_12<=0;
			regfile_signal.reg_file_13<=0;
			regfile_signal.reg_file_14<=0;
			regfile_signal.reg_file_15<=0;
			regfile_signal.reg_file_16<=0;
			regfile_signal.reg_file_17<=0;
			regfile_signal.reg_file_18<=0;
			regfile_signal.reg_file_19<=0;
			regfile_signal.reg_file_20<=0;
			regfile_signal.reg_file_21<=0;
			regfile_signal.reg_file_22<=0;
			regfile_signal.reg_file_23<=0;
			regfile_signal.reg_file_24<=0;
			regfile_signal.reg_file_25<=0;
			regfile_signal.reg_file_26<=0;
			regfile_signal.reg_file_27<=0;
			regfile_signal.reg_file_28<=0;
			regfile_signal.reg_file_29<=0;
			regfile_signal.reg_file_30<=0;
			regfile_signal.reg_file_31<=0;
			regfileWrite_signal.dst<=0;
			regfileWrite_signal.dstData<=0;
			regfileWrite_signal.exception<=0;
			sysRES_signal<=true;
			target_prv_signal:= (others => 0);
			toMemoryData_signal.addrIn<=0;
			toMemoryData_signal.dataIn<=0;
			toMemoryData_signal.mask<=MT_B;
			toMemoryData_signal.req<=ME_RD;
			to_mmu_signal.accesstype<=FETCH;
			to_mmu_signal.data<=0;
			to_mmu_signal.exception_in<=0;
			to_mmu_signal.lrsc<=LR;
			to_mmu_signal.mask<=MT_B;
			to_mmu_signal.mstatus<=0;
			to_mmu_signal.prv<=0;
			to_mmu_signal.reset_lrsc<=0;
			to_mmu_signal.satp<=0;
			to_mmu_signal.v_addr<=0;
			write_signal:= (others => 0);
			xcause_signal:= (others => 0);
			xstatus_mask_signal:= (others => 0);
			xtval_signal:= (others => 0);
			xtvec_signal:= (others => 0);
			ecall_isa_Port_notify <= false;
			fromMemoryPort_notify <= false;
			isa_ecall_Port_notify <= false;
			toMemoryPort_notify <= true;
			toRegsPort_notify <= false;
		 else
		 if section = execute then
		 -- FILL OUT HERE;
		 end if;
		 if section = fetch then
		 -- FILL OUT HERE;
		 end if;
		 end if;
	 end if;
	 end process;
end ISA_arch;
