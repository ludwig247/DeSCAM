library ieee;
use IEEE.numeric_std.all;

package TestBasic12_types is
type TestBasic12_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic12_types;
