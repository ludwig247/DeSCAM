library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestBasic6_types is
end package TestBasic6_types;