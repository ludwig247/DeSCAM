library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave11_types is
type TestMasterSlave11_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave11_types;
