package testmasterslave4_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave4_SECTIONS;

endpackage
