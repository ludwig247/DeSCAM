package testmasterslave0_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave0_SECTIONS;

endpackage
