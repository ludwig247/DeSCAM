library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestArray0_types is
end package TestArray0_types;