package SCAM_Model_types is
subtype bool is Boolean;
subtype int is Integer;
type baudgen_SECTIONS is (RUN);
end package SCAM_Model_types;
