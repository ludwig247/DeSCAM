library ieee;
use IEEE.numeric_std.all;

package TestBasic22_types is
type TestBasic22_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic22_types;
