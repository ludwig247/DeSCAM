library ieee;
use IEEE.numeric_std.all;

package TestBasic2_types is
type TestBasic2_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic2_types;
