library ieee;
use IEEE.numeric_std.all;

package TestBasic18_types is
type TestBasic18_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic18_types;
