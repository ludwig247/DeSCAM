package testbasic17_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic17_SECTIONS;

endpackage
