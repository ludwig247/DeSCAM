library ieee;
use IEEE.numeric_std.all;

package TestBasic17_types is
type TestBasic17_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic17_types;
