library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestBasic0_types is
type Sections is (SECTION_A, SECTION_B);
end package TestBasic0_types;