library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave2_types is
type TestMasterSlave2_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave2_types;
