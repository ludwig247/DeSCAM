package testbasic8_types;

endpackage