library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave8_types is
type TestMasterSlave8_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave8_types;

