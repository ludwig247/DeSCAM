library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package top_level_types is
subtype bool is Boolean;
type int_2 is array(1 downto 0) of signed(31 downto 0);
end package top_level_types;