import top_level_types::*;
import isa_new_types::*;

module ISA_new (
	input logic clk,
	input logic rst,
	input MEtoCU_IF fromMemoryPort,
	input logic fromMemoryPort_sync,
	output logic fromMemoryPort_notify,
	input unsigned_32 fromRegsPort,
	output CUtoME_IF toMemoryPort,
	input logic toMemoryPort_sync,
	output logic toMemoryPort_notify,
	output RegfileWriteType toRegsPort,
	output logic toRegsPort_notify
	);
	
	bit[31:0] pcReg_signal;
	Phases phase;

	always_ff @(posedge clk, posedge rst) begin
		bit[31:0] encodedInstr;
		EncType opcode;
		logic[31:0] aluOp1;
		logic[31:0] aluOp2;
		logic[31:0] aluResult;
		
		if (rst) begin
			phase <= fetch_ph;
			pcReg_signal = 0;
			toRegsPort.dst <= 0;
			toRegsPort.dstdata <= 0;
			fromMemoryPort_notify <= 1'b0;
			toMemoryPort_notify <= 1'b1;
			toRegsPort_notify <= 1'b0;
			toMemoryPort.addrin <= 1'b0;
			toMemoryPort.datain <= 32'b0;
			toMemoryPort.mask <= mt_w;
			toMemoryPort.req <= me_rd;
		end 
		else begin
			case (phase)
				fetch_ph: begin
			
					toRegsPort_notify <= 1'b0;

					if (toMemoryPort_sync == 1'b1) begin
						toMemoryPort_notify <= 1'b0;
						fromMemoryPort_notify <= 1'b1;
						phase <= execute_ph;
					end
				end
				execute_ph: begin
					if(fromMemoryPort_sync == 1'b1) begin
						fromMemoryPort_notify <= 1'b0;
						toMemoryPort_notify <= 1'b1;

						encodedInstr = fromMemoryPort.loadeddata;
						opcode = get_enc_type(encodedInstr);
						aluOp1 = fromRegsPort[encodedInstr[19:15]]; //rs1 = encodedInstr[19:15]
						aluOp2 = fromRegsPort[encodedInstr[24:20]]; //rs2 = encodedInstr[24:20]
						aluResult = get_alu_result(get_alu_funct(get_instr_type(encodedInstr)), aluOp1, aluOp2);

						if (opcode == enc_r || opcode == enc_i_i) begin
							toRegsPort.dst <= encodedInstr[11:7]; //rd = encodedInstr[11:7]
							toRegsPort.dstdata <= aluResult;
							toRegsPort_notify <= 1'b1;

							pcReg_signal += 4;
							toMemoryPort.addrin <= pcReg_signal;

							phase <= fetch_ph;
						end
						else if (opcode == enc_b) begin
							pcReg_signal = branch_PC_calculation(encodedInstr, aluResult, pcReg_signal);
							toMemoryPort.addrin <= pcReg_signal;
							phase <= fetch_ph;	
						end	
						else if (opcode == enc_s || opcode == enc_i_l) begin	
							aluOp2 = get_immediate(encodedInstr);
							aluResult = get_alu_result(alu_add, aluOp1, aluOp2);
							toMemoryPort.mask <= get_memory_mask(get_instr_type(encodedInstr));
							toMemoryPort.addrin <= aluResult;

							if(opcode == enc_s) begin
								toMemoryPort.req <= me_wr;
								toMemoryPort.datain <= aluOp2;
								phase <= Store;
							end
							else begin	
								toMemoryPort.datain <= 1'b0;
								toMemoryPort.req <= me_rd;
								toRegsPort.dst <= encodedInstr[11:7]; //rd = encodedInstr[11:7]
								phase <= Load_req;
							end
						end
						else if (opcode == enc_u) begin
							toRegsPort.dst <= encodedInstr[11:7]; //rd = encodedInstr[11:7]
							toRegsPort.dstdata <= get_Enc_U_ALU_result(encodedInstr, pcReg_signal);
							toRegsPort_notify <= 1'b1;
	
							pcReg_signal += 4;
						
							toMemoryPort.addrin <= pcReg_signal;

							phase <= fetch_ph;
						end
						else if (opcode == enc_j || opcode == enc_i_j) begin
							toRegsPort.dst <= encodedInstr[11:7]; //rd = encodedInstr[11:7]
							toRegsPort.dstdata <= pcReg_signal + 4;
							toRegsPort_notify <= 1'b1;
							if(opcode == enc_i_j) pcReg_signal = aluOp1 + get_immediate(encodedInstr);
							else pcReg_signal += get_immediate(encodedInstr);
		
							toMemoryPort.addrin <= pcReg_signal;
		
							phase <= fetch_ph;
						end
						else phase <= fetch_ph;
					end
				end
				Store: begin
					if (toMemoryPort_sync == 1'b1) begin
						toMemoryPort_notify <= 1'b0;
						fromMemoryPort_notify <= 1'b1;
					
						phase <= Store_done;
					end
				end
				Store_done: begin
					if (fromMemoryPort_sync == 1'b1) begin
						fromMemoryPort_notify <= 1'b0;
				
						pcReg_signal = pcReg_signal + 4;

						toMemoryPort_notify <= 1'b1;
						toMemoryPort.addrin <= pcReg_signal;
						toMemoryPort.datain <= 32'b0;
						toMemoryPort.mask   <= mt_w;
						toMemoryPort.req    <= me_rd;
					
						phase <= fetch_ph;
					end
				end
				Load_req: begin
					if (toMemoryPort_sync == 1'b1) begin
						toMemoryPort_notify <= 1'b0;
						fromMemoryPort_notify <= 1'b1;
					
						phase <= Load_done;
					end
				end
				Load_done: begin
					if (fromMemoryPort_sync == 1'b1) begin
						fromMemoryPort_notify <= 1'b0;
	
						toRegsPort.dstdata <= fromMemoryPort.loadeddata;
						toRegsPort_notify  <= 1'b1;

						pcReg_signal = pcReg_signal + 4;

						toMemoryPort_notify <= 1'b1;
						toMemoryPort.addrin <= pcReg_signal;
						toMemoryPort.datain <= 32'b0;
						toMemoryPort.mask   <= mt_w;
						toMemoryPort.req    <= me_rd;
					
						phase <= fetch_ph;
					end
				end
			endcase
		end
	end
endmodule