library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave0_types is
type TestMasterSlave0_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave0_types;
