package testbasic7_types;

	 import top_level_types::*;
endpackage