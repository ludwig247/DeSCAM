package testbasic16_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic16_SECTIONS;

endpackage
