package testfunction0_types;

	typedef enum logic {
		run
	} TestFunction0_SECTIONS;

endpackage
