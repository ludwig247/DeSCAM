library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave5_types is
type TestMasterSlave5_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave5_types;
