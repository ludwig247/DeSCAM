package testarray0_types;

	import scam_model_types::*;
endpackage