package testbasic5_types;

	typedef enum logic {
		run
	} TestBasic5_SECTIONS;

endpackage
