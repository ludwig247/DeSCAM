library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestTernary01_types is
-- No local datatypes implemented!


end package TestTernary01_types;