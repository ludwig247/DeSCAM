module Bus( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_master_in_sync, // @[:@6.4]
  input         io_master_out_sync, // @[:@6.4]
  input         io_slave_in0_sync, // @[:@6.4]
  input         io_slave_in1_sync, // @[:@6.4]
  input         io_slave_in2_sync, // @[:@6.4]
  input         io_slave_in3_sync, // @[:@6.4]
  input         io_slave_out0_sync, // @[:@6.4]
  input         io_slave_out1_sync, // @[:@6.4]
  input         io_slave_out2_sync, // @[:@6.4]
  input         io_slave_out3_sync, // @[:@6.4]
  output        io_master_in_notify, // @[:@6.4]
  output        io_master_out_notify, // @[:@6.4]
  output        io_slave_in0_notify, // @[:@6.4]
  output        io_slave_in1_notify, // @[:@6.4]
  output        io_slave_in2_notify, // @[:@6.4]
  output        io_slave_in3_notify, // @[:@6.4]
  output        io_slave_out0_notify, // @[:@6.4]
  output        io_slave_out1_notify, // @[:@6.4]
  output        io_slave_out2_notify, // @[:@6.4]
  output        io_slave_out3_notify, // @[:@6.4]
  input  [31:0] io_master_in_addr, // @[:@6.4]
  input  [31:0] io_master_in_data, // @[:@6.4]
  input  [31:0] io_master_in_trans_type, // @[:@6.4]
  output [31:0] io_master_out_ack, // @[:@6.4]
  output [31:0] io_master_out_data, // @[:@6.4]
  input  [31:0] io_slave_in0_ack, // @[:@6.4]
  input  [31:0] io_slave_in0_data, // @[:@6.4]
  input  [31:0] io_slave_in1_ack, // @[:@6.4]
  input  [31:0] io_slave_in1_data, // @[:@6.4]
  input  [31:0] io_slave_in2_ack, // @[:@6.4]
  input  [31:0] io_slave_in2_data, // @[:@6.4]
  input  [31:0] io_slave_in3_ack, // @[:@6.4]
  input  [31:0] io_slave_in3_data, // @[:@6.4]
  output [31:0] io_slave_out0_addr, // @[:@6.4]
  output [31:0] io_slave_out0_data, // @[:@6.4]
  output [31:0] io_slave_out0_trans_type, // @[:@6.4]
  output [31:0] io_slave_out1_addr, // @[:@6.4]
  output [31:0] io_slave_out1_data, // @[:@6.4]
  output [31:0] io_slave_out1_trans_type, // @[:@6.4]
  output [31:0] io_slave_out2_addr, // @[:@6.4]
  output [31:0] io_slave_out2_data, // @[:@6.4]
  output [31:0] io_slave_out2_trans_type, // @[:@6.4]
  output [31:0] io_slave_out3_addr, // @[:@6.4]
  output [31:0] io_slave_out3_data, // @[:@6.4]
  output [31:0] io_slave_out3_trans_type // @[:@6.4]
);
  reg  master_in_notify_r; // @[Bus.scala 50:37:@8.4]
  reg [31:0] _RAND_0;
  reg  master_out_notify_r; // @[Bus.scala 51:38:@9.4]
  reg [31:0] _RAND_1;
  reg  slave_in0_notify_r; // @[Bus.scala 52:37:@10.4]
  reg [31:0] _RAND_2;
  reg  slave_in1_notify_r; // @[Bus.scala 53:37:@11.4]
  reg [31:0] _RAND_3;
  reg  slave_in2_notify_r; // @[Bus.scala 54:37:@12.4]
  reg [31:0] _RAND_4;
  reg  slave_in3_notify_r; // @[Bus.scala 55:37:@13.4]
  reg [31:0] _RAND_5;
  reg  slave_out0_notify_r; // @[Bus.scala 56:38:@14.4]
  reg [31:0] _RAND_6;
  reg  slave_out1_notify_r; // @[Bus.scala 57:38:@15.4]
  reg [31:0] _RAND_7;
  reg  slave_out2_notify_r; // @[Bus.scala 58:38:@16.4]
  reg [31:0] _RAND_8;
  reg  slave_out3_notify_r; // @[Bus.scala 59:38:@17.4]
  reg [31:0] _RAND_9;
  reg [31:0] master_out_r_ack; // @[Bus.scala 60:31:@18.4]
  reg [31:0] _RAND_10;
  reg [31:0] master_out_r_data; // @[Bus.scala 60:31:@18.4]
  reg [31:0] _RAND_11;
  reg [31:0] slave_out0_r_addr; // @[Bus.scala 61:31:@19.4]
  reg [31:0] _RAND_12;
  reg [31:0] slave_out0_r_data; // @[Bus.scala 61:31:@19.4]
  reg [31:0] _RAND_13;
  reg [31:0] slave_out0_r_trans_type; // @[Bus.scala 61:31:@19.4]
  reg [31:0] _RAND_14;
  reg [31:0] slave_out1_r_addr; // @[Bus.scala 62:31:@20.4]
  reg [31:0] _RAND_15;
  reg [31:0] slave_out1_r_data; // @[Bus.scala 62:31:@20.4]
  reg [31:0] _RAND_16;
  reg [31:0] slave_out1_r_trans_type; // @[Bus.scala 62:31:@20.4]
  reg [31:0] _RAND_17;
  reg [31:0] slave_out2_r_addr; // @[Bus.scala 63:31:@21.4]
  reg [31:0] _RAND_18;
  reg [31:0] slave_out2_r_data; // @[Bus.scala 63:31:@21.4]
  reg [31:0] _RAND_19;
  reg [31:0] slave_out2_r_trans_type; // @[Bus.scala 63:31:@21.4]
  reg [31:0] _RAND_20;
  reg [31:0] slave_out3_r_addr; // @[Bus.scala 64:31:@22.4]
  reg [31:0] _RAND_21;
  reg [31:0] slave_out3_r_data; // @[Bus.scala 64:31:@22.4]
  reg [31:0] _RAND_22;
  reg [31:0] slave_out3_r_trans_type; // @[Bus.scala 64:31:@22.4]
  reg [31:0] _RAND_23;
  reg [31:0] req_signal_r_addr; // @[Bus.scala 65:31:@23.4]
  reg [31:0] _RAND_24;
  reg [31:0] req_signal_r_data; // @[Bus.scala 65:31:@23.4]
  reg [31:0] _RAND_25;
  reg [31:0] req_signal_r_trans_type; // @[Bus.scala 65:31:@23.4]
  reg [31:0] _RAND_26;
  reg [31:0] resp_signal_r_ack; // @[Bus.scala 66:32:@24.4]
  reg [31:0] _RAND_27;
  reg [31:0] resp_signal_r_data; // @[Bus.scala 66:32:@24.4]
  reg [31:0] _RAND_28;
  reg [3:0] state_r; // @[Bus.scala 67:26:@25.4]
  reg [31:0] _RAND_29;
  wire  _T_97; // @[Bus.scala 92:30:@46.6]
  wire  _T_98; // @[Bus.scala 93:44:@48.8]
  wire  _T_100; // @[Bus.scala 93:30:@49.8]
  wire  _T_102; // @[Bus.scala 94:57:@51.10]
  wire  _T_104; // @[Bus.scala 95:65:@53.12]
  wire [3:0] _GEN_0; // @[Bus.scala 96:73:@55.14]
  wire [31:0] _GEN_1; // @[Bus.scala 96:73:@55.14]
  wire [31:0] _GEN_2; // @[Bus.scala 96:73:@55.14]
  wire [31:0] _GEN_3; // @[Bus.scala 96:73:@55.14]
  wire [31:0] _GEN_6; // @[Bus.scala 96:73:@55.14]
  wire [31:0] _GEN_7; // @[Bus.scala 96:73:@55.14]
  wire [31:0] _GEN_8; // @[Bus.scala 96:73:@55.14]
  wire  _GEN_9; // @[Bus.scala 96:73:@55.14]
  wire  _GEN_10; // @[Bus.scala 96:73:@55.14]
  wire  _GEN_11; // @[Bus.scala 96:73:@55.14]
  wire  _GEN_12; // @[Bus.scala 96:73:@55.14]
  wire  _GEN_13; // @[Bus.scala 96:73:@55.14]
  wire  _GEN_14; // @[Bus.scala 96:73:@55.14]
  wire  _GEN_15; // @[Bus.scala 96:73:@55.14]
  wire  _GEN_16; // @[Bus.scala 96:73:@55.14]
  wire  _GEN_17; // @[Bus.scala 96:73:@55.14]
  wire  _GEN_18; // @[Bus.scala 96:73:@55.14]
  wire [3:0] _GEN_19; // @[Bus.scala 95:80:@54.12]
  wire [31:0] _GEN_20; // @[Bus.scala 95:80:@54.12]
  wire [31:0] _GEN_21; // @[Bus.scala 95:80:@54.12]
  wire [31:0] _GEN_22; // @[Bus.scala 95:80:@54.12]
  wire [31:0] _GEN_25; // @[Bus.scala 95:80:@54.12]
  wire [31:0] _GEN_26; // @[Bus.scala 95:80:@54.12]
  wire [31:0] _GEN_27; // @[Bus.scala 95:80:@54.12]
  wire  _GEN_28; // @[Bus.scala 95:80:@54.12]
  wire  _GEN_29; // @[Bus.scala 95:80:@54.12]
  wire  _GEN_30; // @[Bus.scala 95:80:@54.12]
  wire  _GEN_31; // @[Bus.scala 95:80:@54.12]
  wire  _GEN_32; // @[Bus.scala 95:80:@54.12]
  wire  _GEN_33; // @[Bus.scala 95:80:@54.12]
  wire  _GEN_34; // @[Bus.scala 95:80:@54.12]
  wire  _GEN_35; // @[Bus.scala 95:80:@54.12]
  wire  _GEN_36; // @[Bus.scala 95:80:@54.12]
  wire  _GEN_37; // @[Bus.scala 95:80:@54.12]
  wire [3:0] _GEN_38; // @[Bus.scala 94:72:@52.10]
  wire [31:0] _GEN_39; // @[Bus.scala 94:72:@52.10]
  wire [31:0] _GEN_40; // @[Bus.scala 94:72:@52.10]
  wire [31:0] _GEN_41; // @[Bus.scala 94:72:@52.10]
  wire [31:0] _GEN_44; // @[Bus.scala 94:72:@52.10]
  wire [31:0] _GEN_45; // @[Bus.scala 94:72:@52.10]
  wire [31:0] _GEN_46; // @[Bus.scala 94:72:@52.10]
  wire  _GEN_47; // @[Bus.scala 94:72:@52.10]
  wire  _GEN_48; // @[Bus.scala 94:72:@52.10]
  wire  _GEN_49; // @[Bus.scala 94:72:@52.10]
  wire  _GEN_50; // @[Bus.scala 94:72:@52.10]
  wire  _GEN_51; // @[Bus.scala 94:72:@52.10]
  wire  _GEN_52; // @[Bus.scala 94:72:@52.10]
  wire  _GEN_53; // @[Bus.scala 94:72:@52.10]
  wire  _GEN_54; // @[Bus.scala 94:72:@52.10]
  wire  _GEN_55; // @[Bus.scala 94:72:@52.10]
  wire  _GEN_56; // @[Bus.scala 94:72:@52.10]
  wire [3:0] _GEN_57; // @[Bus.scala 93:74:@50.8]
  wire [31:0] _GEN_58; // @[Bus.scala 93:74:@50.8]
  wire [31:0] _GEN_59; // @[Bus.scala 93:74:@50.8]
  wire [31:0] _GEN_60; // @[Bus.scala 93:74:@50.8]
  wire [31:0] _GEN_63; // @[Bus.scala 93:74:@50.8]
  wire [31:0] _GEN_64; // @[Bus.scala 93:74:@50.8]
  wire [31:0] _GEN_65; // @[Bus.scala 93:74:@50.8]
  wire  _GEN_66; // @[Bus.scala 93:74:@50.8]
  wire  _GEN_67; // @[Bus.scala 93:74:@50.8]
  wire  _GEN_68; // @[Bus.scala 93:74:@50.8]
  wire  _GEN_69; // @[Bus.scala 93:74:@50.8]
  wire  _GEN_70; // @[Bus.scala 93:74:@50.8]
  wire  _GEN_71; // @[Bus.scala 93:74:@50.8]
  wire  _GEN_72; // @[Bus.scala 93:74:@50.8]
  wire  _GEN_73; // @[Bus.scala 93:74:@50.8]
  wire  _GEN_74; // @[Bus.scala 93:74:@50.8]
  wire  _GEN_75; // @[Bus.scala 93:74:@50.8]
  wire [3:0] _GEN_76; // @[Bus.scala 92:41:@47.6]
  wire [31:0] _GEN_77; // @[Bus.scala 92:41:@47.6]
  wire [31:0] _GEN_78; // @[Bus.scala 92:41:@47.6]
  wire [31:0] _GEN_79; // @[Bus.scala 92:41:@47.6]
  wire [31:0] _GEN_82; // @[Bus.scala 92:41:@47.6]
  wire [31:0] _GEN_83; // @[Bus.scala 92:41:@47.6]
  wire [31:0] _GEN_84; // @[Bus.scala 92:41:@47.6]
  wire  _GEN_85; // @[Bus.scala 92:41:@47.6]
  wire  _GEN_86; // @[Bus.scala 92:41:@47.6]
  wire  _GEN_87; // @[Bus.scala 92:41:@47.6]
  wire  _GEN_88; // @[Bus.scala 92:41:@47.6]
  wire  _GEN_89; // @[Bus.scala 92:41:@47.6]
  wire  _GEN_90; // @[Bus.scala 92:41:@47.6]
  wire  _GEN_91; // @[Bus.scala 92:41:@47.6]
  wire  _GEN_92; // @[Bus.scala 92:41:@47.6]
  wire  _GEN_93; // @[Bus.scala 92:41:@47.6]
  wire  _GEN_94; // @[Bus.scala 92:41:@47.6]
  wire [3:0] _GEN_95; // @[Bus.scala 125:73:@88.14]
  wire [31:0] _GEN_96; // @[Bus.scala 125:73:@88.14]
  wire [31:0] _GEN_97; // @[Bus.scala 125:73:@88.14]
  wire [31:0] _GEN_98; // @[Bus.scala 125:73:@88.14]
  wire [31:0] _GEN_101; // @[Bus.scala 125:73:@88.14]
  wire [31:0] _GEN_102; // @[Bus.scala 125:73:@88.14]
  wire [31:0] _GEN_103; // @[Bus.scala 125:73:@88.14]
  wire  _GEN_104; // @[Bus.scala 125:73:@88.14]
  wire  _GEN_105; // @[Bus.scala 125:73:@88.14]
  wire  _GEN_106; // @[Bus.scala 125:73:@88.14]
  wire  _GEN_107; // @[Bus.scala 125:73:@88.14]
  wire  _GEN_108; // @[Bus.scala 125:73:@88.14]
  wire  _GEN_109; // @[Bus.scala 125:73:@88.14]
  wire  _GEN_110; // @[Bus.scala 125:73:@88.14]
  wire  _GEN_111; // @[Bus.scala 125:73:@88.14]
  wire  _GEN_112; // @[Bus.scala 125:73:@88.14]
  wire  _GEN_113; // @[Bus.scala 125:73:@88.14]
  wire [3:0] _GEN_114; // @[Bus.scala 124:80:@87.12]
  wire [31:0] _GEN_115; // @[Bus.scala 124:80:@87.12]
  wire [31:0] _GEN_116; // @[Bus.scala 124:80:@87.12]
  wire [31:0] _GEN_117; // @[Bus.scala 124:80:@87.12]
  wire [31:0] _GEN_120; // @[Bus.scala 124:80:@87.12]
  wire [31:0] _GEN_121; // @[Bus.scala 124:80:@87.12]
  wire [31:0] _GEN_122; // @[Bus.scala 124:80:@87.12]
  wire  _GEN_123; // @[Bus.scala 124:80:@87.12]
  wire  _GEN_124; // @[Bus.scala 124:80:@87.12]
  wire  _GEN_125; // @[Bus.scala 124:80:@87.12]
  wire  _GEN_126; // @[Bus.scala 124:80:@87.12]
  wire  _GEN_127; // @[Bus.scala 124:80:@87.12]
  wire  _GEN_128; // @[Bus.scala 124:80:@87.12]
  wire  _GEN_129; // @[Bus.scala 124:80:@87.12]
  wire  _GEN_130; // @[Bus.scala 124:80:@87.12]
  wire  _GEN_131; // @[Bus.scala 124:80:@87.12]
  wire  _GEN_132; // @[Bus.scala 124:80:@87.12]
  wire [3:0] _GEN_133; // @[Bus.scala 123:72:@85.10]
  wire [31:0] _GEN_134; // @[Bus.scala 123:72:@85.10]
  wire [31:0] _GEN_135; // @[Bus.scala 123:72:@85.10]
  wire [31:0] _GEN_136; // @[Bus.scala 123:72:@85.10]
  wire [31:0] _GEN_139; // @[Bus.scala 123:72:@85.10]
  wire [31:0] _GEN_140; // @[Bus.scala 123:72:@85.10]
  wire [31:0] _GEN_141; // @[Bus.scala 123:72:@85.10]
  wire  _GEN_142; // @[Bus.scala 123:72:@85.10]
  wire  _GEN_143; // @[Bus.scala 123:72:@85.10]
  wire  _GEN_144; // @[Bus.scala 123:72:@85.10]
  wire  _GEN_145; // @[Bus.scala 123:72:@85.10]
  wire  _GEN_146; // @[Bus.scala 123:72:@85.10]
  wire  _GEN_147; // @[Bus.scala 123:72:@85.10]
  wire  _GEN_148; // @[Bus.scala 123:72:@85.10]
  wire  _GEN_149; // @[Bus.scala 123:72:@85.10]
  wire  _GEN_150; // @[Bus.scala 123:72:@85.10]
  wire  _GEN_151; // @[Bus.scala 123:72:@85.10]
  wire [3:0] _GEN_152; // @[Bus.scala 122:73:@83.8]
  wire [31:0] _GEN_153; // @[Bus.scala 122:73:@83.8]
  wire [31:0] _GEN_154; // @[Bus.scala 122:73:@83.8]
  wire [31:0] _GEN_155; // @[Bus.scala 122:73:@83.8]
  wire [31:0] _GEN_158; // @[Bus.scala 122:73:@83.8]
  wire [31:0] _GEN_159; // @[Bus.scala 122:73:@83.8]
  wire [31:0] _GEN_160; // @[Bus.scala 122:73:@83.8]
  wire  _GEN_161; // @[Bus.scala 122:73:@83.8]
  wire  _GEN_162; // @[Bus.scala 122:73:@83.8]
  wire  _GEN_163; // @[Bus.scala 122:73:@83.8]
  wire  _GEN_164; // @[Bus.scala 122:73:@83.8]
  wire  _GEN_165; // @[Bus.scala 122:73:@83.8]
  wire  _GEN_166; // @[Bus.scala 122:73:@83.8]
  wire  _GEN_167; // @[Bus.scala 122:73:@83.8]
  wire  _GEN_168; // @[Bus.scala 122:73:@83.8]
  wire  _GEN_169; // @[Bus.scala 122:73:@83.8]
  wire  _GEN_170; // @[Bus.scala 122:73:@83.8]
  wire [3:0] _GEN_171; // @[Bus.scala 121:41:@81.6]
  wire [31:0] _GEN_172; // @[Bus.scala 121:41:@81.6]
  wire [31:0] _GEN_173; // @[Bus.scala 121:41:@81.6]
  wire [31:0] _GEN_174; // @[Bus.scala 121:41:@81.6]
  wire [31:0] _GEN_177; // @[Bus.scala 121:41:@81.6]
  wire [31:0] _GEN_178; // @[Bus.scala 121:41:@81.6]
  wire [31:0] _GEN_179; // @[Bus.scala 121:41:@81.6]
  wire  _GEN_180; // @[Bus.scala 121:41:@81.6]
  wire  _GEN_181; // @[Bus.scala 121:41:@81.6]
  wire  _GEN_182; // @[Bus.scala 121:41:@81.6]
  wire  _GEN_183; // @[Bus.scala 121:41:@81.6]
  wire  _GEN_184; // @[Bus.scala 121:41:@81.6]
  wire  _GEN_185; // @[Bus.scala 121:41:@81.6]
  wire  _GEN_186; // @[Bus.scala 121:41:@81.6]
  wire  _GEN_187; // @[Bus.scala 121:41:@81.6]
  wire  _GEN_188; // @[Bus.scala 121:41:@81.6]
  wire  _GEN_189; // @[Bus.scala 121:41:@81.6]
  wire  _T_138; // @[Bus.scala 152:88:@118.10]
  wire  _T_140; // @[Bus.scala 152:76:@119.10]
  wire  _T_141; // @[Bus.scala 152:73:@120.10]
  wire  _T_143; // @[Bus.scala 152:38:@121.10]
  wire  _T_145; // @[Bus.scala 153:67:@123.12]
  wire  _T_147; // @[Bus.scala 153:97:@124.12]
  wire  _T_149; // @[Bus.scala 153:84:@125.12]
  wire  _T_150; // @[Bus.scala 153:81:@126.12]
  wire  _T_152; // @[Bus.scala 153:46:@127.12]
  wire  _T_154; // @[Bus.scala 154:75:@129.14]
  wire  _T_156; // @[Bus.scala 154:106:@130.14]
  wire  _T_158; // @[Bus.scala 154:93:@131.14]
  wire  _T_159; // @[Bus.scala 154:90:@132.14]
  wire  _T_161; // @[Bus.scala 154:54:@133.14]
  wire  _T_163; // @[Bus.scala 155:83:@135.16]
  wire  _T_165; // @[Bus.scala 155:114:@136.16]
  wire  _T_167; // @[Bus.scala 155:101:@137.16]
  wire  _T_168; // @[Bus.scala 155:98:@138.16]
  wire  _T_170; // @[Bus.scala 155:62:@139.16]
  wire [3:0] _GEN_190; // @[Bus.scala 156:89:@141.18]
  wire [31:0] _GEN_191; // @[Bus.scala 156:89:@141.18]
  wire [31:0] _GEN_192; // @[Bus.scala 156:89:@141.18]
  wire [31:0] _GEN_193; // @[Bus.scala 156:89:@141.18]
  wire [31:0] _GEN_194; // @[Bus.scala 156:89:@141.18]
  wire [31:0] _GEN_195; // @[Bus.scala 156:89:@141.18]
  wire [31:0] _GEN_196; // @[Bus.scala 156:89:@141.18]
  wire [31:0] _GEN_197; // @[Bus.scala 156:89:@141.18]
  wire  _GEN_198; // @[Bus.scala 156:89:@141.18]
  wire  _GEN_199; // @[Bus.scala 156:89:@141.18]
  wire  _GEN_200; // @[Bus.scala 156:89:@141.18]
  wire  _GEN_201; // @[Bus.scala 156:89:@141.18]
  wire  _GEN_202; // @[Bus.scala 156:89:@141.18]
  wire  _GEN_203; // @[Bus.scala 156:89:@141.18]
  wire  _GEN_204; // @[Bus.scala 156:89:@141.18]
  wire  _GEN_205; // @[Bus.scala 156:89:@141.18]
  wire  _GEN_206; // @[Bus.scala 156:89:@141.18]
  wire  _GEN_207; // @[Bus.scala 156:89:@141.18]
  wire [3:0] _GEN_208; // @[Bus.scala 155:138:@140.16]
  wire [31:0] _GEN_209; // @[Bus.scala 155:138:@140.16]
  wire [31:0] _GEN_210; // @[Bus.scala 155:138:@140.16]
  wire [31:0] _GEN_211; // @[Bus.scala 155:138:@140.16]
  wire [31:0] _GEN_212; // @[Bus.scala 155:138:@140.16]
  wire [31:0] _GEN_213; // @[Bus.scala 155:138:@140.16]
  wire [31:0] _GEN_214; // @[Bus.scala 155:138:@140.16]
  wire [31:0] _GEN_215; // @[Bus.scala 155:138:@140.16]
  wire  _GEN_216; // @[Bus.scala 155:138:@140.16]
  wire  _GEN_217; // @[Bus.scala 155:138:@140.16]
  wire  _GEN_218; // @[Bus.scala 155:138:@140.16]
  wire  _GEN_219; // @[Bus.scala 155:138:@140.16]
  wire  _GEN_220; // @[Bus.scala 155:138:@140.16]
  wire  _GEN_221; // @[Bus.scala 155:138:@140.16]
  wire  _GEN_222; // @[Bus.scala 155:138:@140.16]
  wire  _GEN_223; // @[Bus.scala 155:138:@140.16]
  wire  _GEN_224; // @[Bus.scala 155:138:@140.16]
  wire  _GEN_225; // @[Bus.scala 155:138:@140.16]
  wire [3:0] _GEN_226; // @[Bus.scala 154:130:@134.14]
  wire [31:0] _GEN_227; // @[Bus.scala 154:130:@134.14]
  wire [31:0] _GEN_228; // @[Bus.scala 154:130:@134.14]
  wire [31:0] _GEN_229; // @[Bus.scala 154:130:@134.14]
  wire [31:0] _GEN_230; // @[Bus.scala 154:130:@134.14]
  wire [31:0] _GEN_231; // @[Bus.scala 154:130:@134.14]
  wire [31:0] _GEN_232; // @[Bus.scala 154:130:@134.14]
  wire [31:0] _GEN_233; // @[Bus.scala 154:130:@134.14]
  wire  _GEN_234; // @[Bus.scala 154:130:@134.14]
  wire  _GEN_235; // @[Bus.scala 154:130:@134.14]
  wire  _GEN_236; // @[Bus.scala 154:130:@134.14]
  wire  _GEN_237; // @[Bus.scala 154:130:@134.14]
  wire  _GEN_238; // @[Bus.scala 154:130:@134.14]
  wire  _GEN_239; // @[Bus.scala 154:130:@134.14]
  wire  _GEN_240; // @[Bus.scala 154:130:@134.14]
  wire  _GEN_241; // @[Bus.scala 154:130:@134.14]
  wire  _GEN_242; // @[Bus.scala 154:130:@134.14]
  wire  _GEN_243; // @[Bus.scala 154:130:@134.14]
  wire [3:0] _GEN_244; // @[Bus.scala 153:121:@128.12]
  wire [31:0] _GEN_245; // @[Bus.scala 153:121:@128.12]
  wire [31:0] _GEN_246; // @[Bus.scala 153:121:@128.12]
  wire [31:0] _GEN_247; // @[Bus.scala 153:121:@128.12]
  wire [31:0] _GEN_248; // @[Bus.scala 153:121:@128.12]
  wire [31:0] _GEN_249; // @[Bus.scala 153:121:@128.12]
  wire [31:0] _GEN_250; // @[Bus.scala 153:121:@128.12]
  wire [31:0] _GEN_251; // @[Bus.scala 153:121:@128.12]
  wire  _GEN_252; // @[Bus.scala 153:121:@128.12]
  wire  _GEN_253; // @[Bus.scala 153:121:@128.12]
  wire  _GEN_254; // @[Bus.scala 153:121:@128.12]
  wire  _GEN_255; // @[Bus.scala 153:121:@128.12]
  wire  _GEN_256; // @[Bus.scala 153:121:@128.12]
  wire  _GEN_257; // @[Bus.scala 153:121:@128.12]
  wire  _GEN_258; // @[Bus.scala 153:121:@128.12]
  wire  _GEN_259; // @[Bus.scala 153:121:@128.12]
  wire  _GEN_260; // @[Bus.scala 153:121:@128.12]
  wire  _GEN_261; // @[Bus.scala 153:121:@128.12]
  wire [3:0] _GEN_262; // @[Bus.scala 152:112:@122.10]
  wire [31:0] _GEN_263; // @[Bus.scala 152:112:@122.10]
  wire [31:0] _GEN_264; // @[Bus.scala 152:112:@122.10]
  wire [31:0] _GEN_265; // @[Bus.scala 152:112:@122.10]
  wire [31:0] _GEN_266; // @[Bus.scala 152:112:@122.10]
  wire [31:0] _GEN_267; // @[Bus.scala 152:112:@122.10]
  wire [31:0] _GEN_268; // @[Bus.scala 152:112:@122.10]
  wire [31:0] _GEN_269; // @[Bus.scala 152:112:@122.10]
  wire  _GEN_270; // @[Bus.scala 152:112:@122.10]
  wire  _GEN_271; // @[Bus.scala 152:112:@122.10]
  wire  _GEN_272; // @[Bus.scala 152:112:@122.10]
  wire  _GEN_273; // @[Bus.scala 152:112:@122.10]
  wire  _GEN_274; // @[Bus.scala 152:112:@122.10]
  wire  _GEN_275; // @[Bus.scala 152:112:@122.10]
  wire  _GEN_276; // @[Bus.scala 152:112:@122.10]
  wire  _GEN_277; // @[Bus.scala 152:112:@122.10]
  wire  _GEN_278; // @[Bus.scala 152:112:@122.10]
  wire  _GEN_279; // @[Bus.scala 152:112:@122.10]
  wire [3:0] _GEN_280; // @[Bus.scala 151:73:@116.8]
  wire [31:0] _GEN_281; // @[Bus.scala 151:73:@116.8]
  wire [31:0] _GEN_282; // @[Bus.scala 151:73:@116.8]
  wire [31:0] _GEN_283; // @[Bus.scala 151:73:@116.8]
  wire [31:0] _GEN_284; // @[Bus.scala 151:73:@116.8]
  wire [31:0] _GEN_285; // @[Bus.scala 151:73:@116.8]
  wire [31:0] _GEN_286; // @[Bus.scala 151:73:@116.8]
  wire [31:0] _GEN_287; // @[Bus.scala 151:73:@116.8]
  wire  _GEN_288; // @[Bus.scala 151:73:@116.8]
  wire  _GEN_289; // @[Bus.scala 151:73:@116.8]
  wire  _GEN_290; // @[Bus.scala 151:73:@116.8]
  wire  _GEN_291; // @[Bus.scala 151:73:@116.8]
  wire  _GEN_292; // @[Bus.scala 151:73:@116.8]
  wire  _GEN_293; // @[Bus.scala 151:73:@116.8]
  wire  _GEN_294; // @[Bus.scala 151:73:@116.8]
  wire  _GEN_295; // @[Bus.scala 151:73:@116.8]
  wire  _GEN_296; // @[Bus.scala 151:73:@116.8]
  wire  _GEN_297; // @[Bus.scala 151:73:@116.8]
  wire [3:0] _GEN_298; // @[Bus.scala 150:41:@114.6]
  wire [31:0] _GEN_299; // @[Bus.scala 150:41:@114.6]
  wire [31:0] _GEN_300; // @[Bus.scala 150:41:@114.6]
  wire [31:0] _GEN_301; // @[Bus.scala 150:41:@114.6]
  wire [31:0] _GEN_302; // @[Bus.scala 150:41:@114.6]
  wire [31:0] _GEN_303; // @[Bus.scala 150:41:@114.6]
  wire [31:0] _GEN_304; // @[Bus.scala 150:41:@114.6]
  wire [31:0] _GEN_305; // @[Bus.scala 150:41:@114.6]
  wire  _GEN_306; // @[Bus.scala 150:41:@114.6]
  wire  _GEN_307; // @[Bus.scala 150:41:@114.6]
  wire  _GEN_308; // @[Bus.scala 150:41:@114.6]
  wire  _GEN_309; // @[Bus.scala 150:41:@114.6]
  wire  _GEN_310; // @[Bus.scala 150:41:@114.6]
  wire  _GEN_311; // @[Bus.scala 150:41:@114.6]
  wire  _GEN_312; // @[Bus.scala 150:41:@114.6]
  wire  _GEN_313; // @[Bus.scala 150:41:@114.6]
  wire  _GEN_314; // @[Bus.scala 150:41:@114.6]
  wire  _GEN_315; // @[Bus.scala 150:41:@114.6]
  wire  _T_221; // @[Bus.scala 187:76:@193.16]
  wire [3:0] _GEN_316; // @[Bus.scala 188:89:@195.18]
  wire [31:0] _GEN_317; // @[Bus.scala 188:89:@195.18]
  wire [31:0] _GEN_318; // @[Bus.scala 188:89:@195.18]
  wire [31:0] _GEN_319; // @[Bus.scala 188:89:@195.18]
  wire [31:0] _GEN_320; // @[Bus.scala 188:89:@195.18]
  wire [31:0] _GEN_321; // @[Bus.scala 188:89:@195.18]
  wire [31:0] _GEN_322; // @[Bus.scala 188:89:@195.18]
  wire [31:0] _GEN_323; // @[Bus.scala 188:89:@195.18]
  wire  _GEN_324; // @[Bus.scala 188:89:@195.18]
  wire  _GEN_325; // @[Bus.scala 188:89:@195.18]
  wire  _GEN_326; // @[Bus.scala 188:89:@195.18]
  wire  _GEN_327; // @[Bus.scala 188:89:@195.18]
  wire  _GEN_328; // @[Bus.scala 188:89:@195.18]
  wire  _GEN_329; // @[Bus.scala 188:89:@195.18]
  wire  _GEN_330; // @[Bus.scala 188:89:@195.18]
  wire  _GEN_331; // @[Bus.scala 188:89:@195.18]
  wire  _GEN_332; // @[Bus.scala 188:89:@195.18]
  wire  _GEN_333; // @[Bus.scala 188:89:@195.18]
  wire [3:0] _GEN_334; // @[Bus.scala 187:106:@194.16]
  wire [31:0] _GEN_335; // @[Bus.scala 187:106:@194.16]
  wire [31:0] _GEN_336; // @[Bus.scala 187:106:@194.16]
  wire [31:0] _GEN_337; // @[Bus.scala 187:106:@194.16]
  wire [31:0] _GEN_338; // @[Bus.scala 187:106:@194.16]
  wire [31:0] _GEN_339; // @[Bus.scala 187:106:@194.16]
  wire [31:0] _GEN_340; // @[Bus.scala 187:106:@194.16]
  wire [31:0] _GEN_341; // @[Bus.scala 187:106:@194.16]
  wire  _GEN_342; // @[Bus.scala 187:106:@194.16]
  wire  _GEN_343; // @[Bus.scala 187:106:@194.16]
  wire  _GEN_344; // @[Bus.scala 187:106:@194.16]
  wire  _GEN_345; // @[Bus.scala 187:106:@194.16]
  wire  _GEN_346; // @[Bus.scala 187:106:@194.16]
  wire  _GEN_347; // @[Bus.scala 187:106:@194.16]
  wire  _GEN_348; // @[Bus.scala 187:106:@194.16]
  wire  _GEN_349; // @[Bus.scala 187:106:@194.16]
  wire  _GEN_350; // @[Bus.scala 187:106:@194.16]
  wire  _GEN_351; // @[Bus.scala 187:106:@194.16]
  wire [3:0] _GEN_352; // @[Bus.scala 186:130:@192.14]
  wire [31:0] _GEN_353; // @[Bus.scala 186:130:@192.14]
  wire [31:0] _GEN_354; // @[Bus.scala 186:130:@192.14]
  wire [31:0] _GEN_355; // @[Bus.scala 186:130:@192.14]
  wire [31:0] _GEN_356; // @[Bus.scala 186:130:@192.14]
  wire [31:0] _GEN_357; // @[Bus.scala 186:130:@192.14]
  wire [31:0] _GEN_358; // @[Bus.scala 186:130:@192.14]
  wire [31:0] _GEN_359; // @[Bus.scala 186:130:@192.14]
  wire  _GEN_360; // @[Bus.scala 186:130:@192.14]
  wire  _GEN_361; // @[Bus.scala 186:130:@192.14]
  wire  _GEN_362; // @[Bus.scala 186:130:@192.14]
  wire  _GEN_363; // @[Bus.scala 186:130:@192.14]
  wire  _GEN_364; // @[Bus.scala 186:130:@192.14]
  wire  _GEN_365; // @[Bus.scala 186:130:@192.14]
  wire  _GEN_366; // @[Bus.scala 186:130:@192.14]
  wire  _GEN_367; // @[Bus.scala 186:130:@192.14]
  wire  _GEN_368; // @[Bus.scala 186:130:@192.14]
  wire  _GEN_369; // @[Bus.scala 186:130:@192.14]
  wire [3:0] _GEN_370; // @[Bus.scala 185:122:@186.12]
  wire [31:0] _GEN_371; // @[Bus.scala 185:122:@186.12]
  wire [31:0] _GEN_372; // @[Bus.scala 185:122:@186.12]
  wire [31:0] _GEN_373; // @[Bus.scala 185:122:@186.12]
  wire [31:0] _GEN_374; // @[Bus.scala 185:122:@186.12]
  wire [31:0] _GEN_375; // @[Bus.scala 185:122:@186.12]
  wire [31:0] _GEN_376; // @[Bus.scala 185:122:@186.12]
  wire [31:0] _GEN_377; // @[Bus.scala 185:122:@186.12]
  wire  _GEN_378; // @[Bus.scala 185:122:@186.12]
  wire  _GEN_379; // @[Bus.scala 185:122:@186.12]
  wire  _GEN_380; // @[Bus.scala 185:122:@186.12]
  wire  _GEN_381; // @[Bus.scala 185:122:@186.12]
  wire  _GEN_382; // @[Bus.scala 185:122:@186.12]
  wire  _GEN_383; // @[Bus.scala 185:122:@186.12]
  wire  _GEN_384; // @[Bus.scala 185:122:@186.12]
  wire  _GEN_385; // @[Bus.scala 185:122:@186.12]
  wire  _GEN_386; // @[Bus.scala 185:122:@186.12]
  wire  _GEN_387; // @[Bus.scala 185:122:@186.12]
  wire [3:0] _GEN_388; // @[Bus.scala 184:113:@180.10]
  wire [31:0] _GEN_389; // @[Bus.scala 184:113:@180.10]
  wire [31:0] _GEN_390; // @[Bus.scala 184:113:@180.10]
  wire [31:0] _GEN_391; // @[Bus.scala 184:113:@180.10]
  wire [31:0] _GEN_392; // @[Bus.scala 184:113:@180.10]
  wire [31:0] _GEN_393; // @[Bus.scala 184:113:@180.10]
  wire [31:0] _GEN_394; // @[Bus.scala 184:113:@180.10]
  wire [31:0] _GEN_395; // @[Bus.scala 184:113:@180.10]
  wire  _GEN_396; // @[Bus.scala 184:113:@180.10]
  wire  _GEN_397; // @[Bus.scala 184:113:@180.10]
  wire  _GEN_398; // @[Bus.scala 184:113:@180.10]
  wire  _GEN_399; // @[Bus.scala 184:113:@180.10]
  wire  _GEN_400; // @[Bus.scala 184:113:@180.10]
  wire  _GEN_401; // @[Bus.scala 184:113:@180.10]
  wire  _GEN_402; // @[Bus.scala 184:113:@180.10]
  wire  _GEN_403; // @[Bus.scala 184:113:@180.10]
  wire  _GEN_404; // @[Bus.scala 184:113:@180.10]
  wire  _GEN_405; // @[Bus.scala 184:113:@180.10]
  wire [3:0] _GEN_406; // @[Bus.scala 183:104:@174.8]
  wire [31:0] _GEN_407; // @[Bus.scala 183:104:@174.8]
  wire [31:0] _GEN_408; // @[Bus.scala 183:104:@174.8]
  wire [31:0] _GEN_409; // @[Bus.scala 183:104:@174.8]
  wire [31:0] _GEN_410; // @[Bus.scala 183:104:@174.8]
  wire [31:0] _GEN_411; // @[Bus.scala 183:104:@174.8]
  wire [31:0] _GEN_412; // @[Bus.scala 183:104:@174.8]
  wire [31:0] _GEN_413; // @[Bus.scala 183:104:@174.8]
  wire  _GEN_414; // @[Bus.scala 183:104:@174.8]
  wire  _GEN_415; // @[Bus.scala 183:104:@174.8]
  wire  _GEN_416; // @[Bus.scala 183:104:@174.8]
  wire  _GEN_417; // @[Bus.scala 183:104:@174.8]
  wire  _GEN_418; // @[Bus.scala 183:104:@174.8]
  wire  _GEN_419; // @[Bus.scala 183:104:@174.8]
  wire  _GEN_420; // @[Bus.scala 183:104:@174.8]
  wire  _GEN_421; // @[Bus.scala 183:104:@174.8]
  wire  _GEN_422; // @[Bus.scala 183:104:@174.8]
  wire  _GEN_423; // @[Bus.scala 183:104:@174.8]
  wire [3:0] _GEN_424; // @[Bus.scala 182:41:@168.6]
  wire [31:0] _GEN_425; // @[Bus.scala 182:41:@168.6]
  wire [31:0] _GEN_426; // @[Bus.scala 182:41:@168.6]
  wire [31:0] _GEN_427; // @[Bus.scala 182:41:@168.6]
  wire [31:0] _GEN_428; // @[Bus.scala 182:41:@168.6]
  wire [31:0] _GEN_429; // @[Bus.scala 182:41:@168.6]
  wire [31:0] _GEN_430; // @[Bus.scala 182:41:@168.6]
  wire [31:0] _GEN_431; // @[Bus.scala 182:41:@168.6]
  wire  _GEN_432; // @[Bus.scala 182:41:@168.6]
  wire  _GEN_433; // @[Bus.scala 182:41:@168.6]
  wire  _GEN_434; // @[Bus.scala 182:41:@168.6]
  wire  _GEN_435; // @[Bus.scala 182:41:@168.6]
  wire  _GEN_436; // @[Bus.scala 182:41:@168.6]
  wire  _GEN_437; // @[Bus.scala 182:41:@168.6]
  wire  _GEN_438; // @[Bus.scala 182:41:@168.6]
  wire  _GEN_439; // @[Bus.scala 182:41:@168.6]
  wire  _GEN_440; // @[Bus.scala 182:41:@168.6]
  wire  _GEN_441; // @[Bus.scala 182:41:@168.6]
  wire  _T_241; // @[Bus.scala 217:65:@228.12]
  wire [32:0] _T_243; // @[Bus.scala 220:92:@232.16]
  wire [31:0] _T_244; // @[Bus.scala 220:92:@233.16]
  wire [31:0] _T_245; // @[Bus.scala 220:92:@234.16]
  wire [3:0] _GEN_442; // @[Bus.scala 218:73:@230.14]
  wire [31:0] _GEN_443; // @[Bus.scala 218:73:@230.14]
  wire [31:0] _GEN_444; // @[Bus.scala 218:73:@230.14]
  wire [31:0] _GEN_445; // @[Bus.scala 218:73:@230.14]
  wire [31:0] _GEN_446; // @[Bus.scala 218:73:@230.14]
  wire [31:0] _GEN_447; // @[Bus.scala 218:73:@230.14]
  wire [31:0] _GEN_448; // @[Bus.scala 218:73:@230.14]
  wire [31:0] _GEN_449; // @[Bus.scala 218:73:@230.14]
  wire [31:0] _GEN_450; // @[Bus.scala 218:73:@230.14]
  wire  _GEN_451; // @[Bus.scala 218:73:@230.14]
  wire  _GEN_452; // @[Bus.scala 218:73:@230.14]
  wire  _GEN_453; // @[Bus.scala 218:73:@230.14]
  wire  _GEN_454; // @[Bus.scala 218:73:@230.14]
  wire  _GEN_455; // @[Bus.scala 218:73:@230.14]
  wire  _GEN_456; // @[Bus.scala 218:73:@230.14]
  wire  _GEN_457; // @[Bus.scala 218:73:@230.14]
  wire  _GEN_458; // @[Bus.scala 218:73:@230.14]
  wire  _GEN_459; // @[Bus.scala 218:73:@230.14]
  wire  _GEN_460; // @[Bus.scala 218:73:@230.14]
  wire [3:0] _GEN_461; // @[Bus.scala 217:81:@229.12]
  wire [31:0] _GEN_462; // @[Bus.scala 217:81:@229.12]
  wire [31:0] _GEN_463; // @[Bus.scala 217:81:@229.12]
  wire [31:0] _GEN_464; // @[Bus.scala 217:81:@229.12]
  wire [31:0] _GEN_465; // @[Bus.scala 217:81:@229.12]
  wire [31:0] _GEN_466; // @[Bus.scala 217:81:@229.12]
  wire [31:0] _GEN_467; // @[Bus.scala 217:81:@229.12]
  wire [31:0] _GEN_468; // @[Bus.scala 217:81:@229.12]
  wire [31:0] _GEN_469; // @[Bus.scala 217:81:@229.12]
  wire  _GEN_470; // @[Bus.scala 217:81:@229.12]
  wire  _GEN_471; // @[Bus.scala 217:81:@229.12]
  wire  _GEN_472; // @[Bus.scala 217:81:@229.12]
  wire  _GEN_473; // @[Bus.scala 217:81:@229.12]
  wire  _GEN_474; // @[Bus.scala 217:81:@229.12]
  wire  _GEN_475; // @[Bus.scala 217:81:@229.12]
  wire  _GEN_476; // @[Bus.scala 217:81:@229.12]
  wire  _GEN_477; // @[Bus.scala 217:81:@229.12]
  wire  _GEN_478; // @[Bus.scala 217:81:@229.12]
  wire  _GEN_479; // @[Bus.scala 217:81:@229.12]
  wire [3:0] _GEN_480; // @[Bus.scala 216:72:@227.10]
  wire [31:0] _GEN_481; // @[Bus.scala 216:72:@227.10]
  wire [31:0] _GEN_482; // @[Bus.scala 216:72:@227.10]
  wire [31:0] _GEN_483; // @[Bus.scala 216:72:@227.10]
  wire [31:0] _GEN_484; // @[Bus.scala 216:72:@227.10]
  wire [31:0] _GEN_485; // @[Bus.scala 216:72:@227.10]
  wire [31:0] _GEN_486; // @[Bus.scala 216:72:@227.10]
  wire [31:0] _GEN_487; // @[Bus.scala 216:72:@227.10]
  wire [31:0] _GEN_488; // @[Bus.scala 216:72:@227.10]
  wire  _GEN_489; // @[Bus.scala 216:72:@227.10]
  wire  _GEN_490; // @[Bus.scala 216:72:@227.10]
  wire  _GEN_491; // @[Bus.scala 216:72:@227.10]
  wire  _GEN_492; // @[Bus.scala 216:72:@227.10]
  wire  _GEN_493; // @[Bus.scala 216:72:@227.10]
  wire  _GEN_494; // @[Bus.scala 216:72:@227.10]
  wire  _GEN_495; // @[Bus.scala 216:72:@227.10]
  wire  _GEN_496; // @[Bus.scala 216:72:@227.10]
  wire  _GEN_497; // @[Bus.scala 216:72:@227.10]
  wire  _GEN_498; // @[Bus.scala 216:72:@227.10]
  wire [3:0] _GEN_499; // @[Bus.scala 215:74:@225.8]
  wire [31:0] _GEN_500; // @[Bus.scala 215:74:@225.8]
  wire [31:0] _GEN_501; // @[Bus.scala 215:74:@225.8]
  wire [31:0] _GEN_502; // @[Bus.scala 215:74:@225.8]
  wire [31:0] _GEN_503; // @[Bus.scala 215:74:@225.8]
  wire [31:0] _GEN_504; // @[Bus.scala 215:74:@225.8]
  wire [31:0] _GEN_505; // @[Bus.scala 215:74:@225.8]
  wire [31:0] _GEN_506; // @[Bus.scala 215:74:@225.8]
  wire [31:0] _GEN_507; // @[Bus.scala 215:74:@225.8]
  wire  _GEN_508; // @[Bus.scala 215:74:@225.8]
  wire  _GEN_509; // @[Bus.scala 215:74:@225.8]
  wire  _GEN_510; // @[Bus.scala 215:74:@225.8]
  wire  _GEN_511; // @[Bus.scala 215:74:@225.8]
  wire  _GEN_512; // @[Bus.scala 215:74:@225.8]
  wire  _GEN_513; // @[Bus.scala 215:74:@225.8]
  wire  _GEN_514; // @[Bus.scala 215:74:@225.8]
  wire  _GEN_515; // @[Bus.scala 215:74:@225.8]
  wire  _GEN_516; // @[Bus.scala 215:74:@225.8]
  wire  _GEN_517; // @[Bus.scala 215:74:@225.8]
  wire [3:0] _GEN_518; // @[Bus.scala 214:41:@222.6]
  wire [31:0] _GEN_519; // @[Bus.scala 214:41:@222.6]
  wire [31:0] _GEN_520; // @[Bus.scala 214:41:@222.6]
  wire [31:0] _GEN_521; // @[Bus.scala 214:41:@222.6]
  wire [31:0] _GEN_522; // @[Bus.scala 214:41:@222.6]
  wire [31:0] _GEN_523; // @[Bus.scala 214:41:@222.6]
  wire [31:0] _GEN_524; // @[Bus.scala 214:41:@222.6]
  wire [31:0] _GEN_525; // @[Bus.scala 214:41:@222.6]
  wire [31:0] _GEN_526; // @[Bus.scala 214:41:@222.6]
  wire  _GEN_527; // @[Bus.scala 214:41:@222.6]
  wire  _GEN_528; // @[Bus.scala 214:41:@222.6]
  wire  _GEN_529; // @[Bus.scala 214:41:@222.6]
  wire  _GEN_530; // @[Bus.scala 214:41:@222.6]
  wire  _GEN_531; // @[Bus.scala 214:41:@222.6]
  wire  _GEN_532; // @[Bus.scala 214:41:@222.6]
  wire  _GEN_533; // @[Bus.scala 214:41:@222.6]
  wire  _GEN_534; // @[Bus.scala 214:41:@222.6]
  wire  _GEN_535; // @[Bus.scala 214:41:@222.6]
  wire  _GEN_536; // @[Bus.scala 214:41:@222.6]
  wire [3:0] _GEN_537; // @[Bus.scala 247:73:@269.14]
  wire [31:0] _GEN_538; // @[Bus.scala 247:73:@269.14]
  wire [31:0] _GEN_539; // @[Bus.scala 247:73:@269.14]
  wire [31:0] _GEN_540; // @[Bus.scala 247:73:@269.14]
  wire [31:0] _GEN_541; // @[Bus.scala 247:73:@269.14]
  wire [31:0] _GEN_542; // @[Bus.scala 247:73:@269.14]
  wire [31:0] _GEN_543; // @[Bus.scala 247:73:@269.14]
  wire [31:0] _GEN_544; // @[Bus.scala 247:73:@269.14]
  wire [31:0] _GEN_545; // @[Bus.scala 247:73:@269.14]
  wire  _GEN_546; // @[Bus.scala 247:73:@269.14]
  wire  _GEN_547; // @[Bus.scala 247:73:@269.14]
  wire  _GEN_548; // @[Bus.scala 247:73:@269.14]
  wire  _GEN_549; // @[Bus.scala 247:73:@269.14]
  wire  _GEN_550; // @[Bus.scala 247:73:@269.14]
  wire  _GEN_551; // @[Bus.scala 247:73:@269.14]
  wire  _GEN_552; // @[Bus.scala 247:73:@269.14]
  wire  _GEN_553; // @[Bus.scala 247:73:@269.14]
  wire  _GEN_554; // @[Bus.scala 247:73:@269.14]
  wire  _GEN_555; // @[Bus.scala 247:73:@269.14]
  wire [3:0] _GEN_556; // @[Bus.scala 246:81:@268.12]
  wire [31:0] _GEN_557; // @[Bus.scala 246:81:@268.12]
  wire [31:0] _GEN_558; // @[Bus.scala 246:81:@268.12]
  wire [31:0] _GEN_559; // @[Bus.scala 246:81:@268.12]
  wire [31:0] _GEN_560; // @[Bus.scala 246:81:@268.12]
  wire [31:0] _GEN_561; // @[Bus.scala 246:81:@268.12]
  wire [31:0] _GEN_562; // @[Bus.scala 246:81:@268.12]
  wire [31:0] _GEN_563; // @[Bus.scala 246:81:@268.12]
  wire [31:0] _GEN_564; // @[Bus.scala 246:81:@268.12]
  wire  _GEN_565; // @[Bus.scala 246:81:@268.12]
  wire  _GEN_566; // @[Bus.scala 246:81:@268.12]
  wire  _GEN_567; // @[Bus.scala 246:81:@268.12]
  wire  _GEN_568; // @[Bus.scala 246:81:@268.12]
  wire  _GEN_569; // @[Bus.scala 246:81:@268.12]
  wire  _GEN_570; // @[Bus.scala 246:81:@268.12]
  wire  _GEN_571; // @[Bus.scala 246:81:@268.12]
  wire  _GEN_572; // @[Bus.scala 246:81:@268.12]
  wire  _GEN_573; // @[Bus.scala 246:81:@268.12]
  wire  _GEN_574; // @[Bus.scala 246:81:@268.12]
  wire [3:0] _GEN_575; // @[Bus.scala 245:72:@266.10]
  wire [31:0] _GEN_576; // @[Bus.scala 245:72:@266.10]
  wire [31:0] _GEN_577; // @[Bus.scala 245:72:@266.10]
  wire [31:0] _GEN_578; // @[Bus.scala 245:72:@266.10]
  wire [31:0] _GEN_579; // @[Bus.scala 245:72:@266.10]
  wire [31:0] _GEN_580; // @[Bus.scala 245:72:@266.10]
  wire [31:0] _GEN_581; // @[Bus.scala 245:72:@266.10]
  wire [31:0] _GEN_582; // @[Bus.scala 245:72:@266.10]
  wire [31:0] _GEN_583; // @[Bus.scala 245:72:@266.10]
  wire  _GEN_584; // @[Bus.scala 245:72:@266.10]
  wire  _GEN_585; // @[Bus.scala 245:72:@266.10]
  wire  _GEN_586; // @[Bus.scala 245:72:@266.10]
  wire  _GEN_587; // @[Bus.scala 245:72:@266.10]
  wire  _GEN_588; // @[Bus.scala 245:72:@266.10]
  wire  _GEN_589; // @[Bus.scala 245:72:@266.10]
  wire  _GEN_590; // @[Bus.scala 245:72:@266.10]
  wire  _GEN_591; // @[Bus.scala 245:72:@266.10]
  wire  _GEN_592; // @[Bus.scala 245:72:@266.10]
  wire  _GEN_593; // @[Bus.scala 245:72:@266.10]
  wire [3:0] _GEN_594; // @[Bus.scala 244:73:@264.8]
  wire [31:0] _GEN_595; // @[Bus.scala 244:73:@264.8]
  wire [31:0] _GEN_596; // @[Bus.scala 244:73:@264.8]
  wire [31:0] _GEN_597; // @[Bus.scala 244:73:@264.8]
  wire [31:0] _GEN_598; // @[Bus.scala 244:73:@264.8]
  wire [31:0] _GEN_599; // @[Bus.scala 244:73:@264.8]
  wire [31:0] _GEN_600; // @[Bus.scala 244:73:@264.8]
  wire [31:0] _GEN_601; // @[Bus.scala 244:73:@264.8]
  wire [31:0] _GEN_602; // @[Bus.scala 244:73:@264.8]
  wire  _GEN_603; // @[Bus.scala 244:73:@264.8]
  wire  _GEN_604; // @[Bus.scala 244:73:@264.8]
  wire  _GEN_605; // @[Bus.scala 244:73:@264.8]
  wire  _GEN_606; // @[Bus.scala 244:73:@264.8]
  wire  _GEN_607; // @[Bus.scala 244:73:@264.8]
  wire  _GEN_608; // @[Bus.scala 244:73:@264.8]
  wire  _GEN_609; // @[Bus.scala 244:73:@264.8]
  wire  _GEN_610; // @[Bus.scala 244:73:@264.8]
  wire  _GEN_611; // @[Bus.scala 244:73:@264.8]
  wire  _GEN_612; // @[Bus.scala 244:73:@264.8]
  wire [3:0] _GEN_613; // @[Bus.scala 243:41:@262.6]
  wire [31:0] _GEN_614; // @[Bus.scala 243:41:@262.6]
  wire [31:0] _GEN_615; // @[Bus.scala 243:41:@262.6]
  wire [31:0] _GEN_616; // @[Bus.scala 243:41:@262.6]
  wire [31:0] _GEN_617; // @[Bus.scala 243:41:@262.6]
  wire [31:0] _GEN_618; // @[Bus.scala 243:41:@262.6]
  wire [31:0] _GEN_619; // @[Bus.scala 243:41:@262.6]
  wire [31:0] _GEN_620; // @[Bus.scala 243:41:@262.6]
  wire [31:0] _GEN_621; // @[Bus.scala 243:41:@262.6]
  wire  _GEN_622; // @[Bus.scala 243:41:@262.6]
  wire  _GEN_623; // @[Bus.scala 243:41:@262.6]
  wire  _GEN_624; // @[Bus.scala 243:41:@262.6]
  wire  _GEN_625; // @[Bus.scala 243:41:@262.6]
  wire  _GEN_626; // @[Bus.scala 243:41:@262.6]
  wire  _GEN_627; // @[Bus.scala 243:41:@262.6]
  wire  _GEN_628; // @[Bus.scala 243:41:@262.6]
  wire  _GEN_629; // @[Bus.scala 243:41:@262.6]
  wire  _GEN_630; // @[Bus.scala 243:41:@262.6]
  wire  _GEN_631; // @[Bus.scala 243:41:@262.6]
  wire  _T_293; // @[Bus.scala 275:65:@307.12]
  wire [32:0] _T_295; // @[Bus.scala 278:93:@311.16]
  wire [31:0] _T_296; // @[Bus.scala 278:93:@312.16]
  wire [31:0] _T_297; // @[Bus.scala 278:93:@313.16]
  wire [3:0] _GEN_632; // @[Bus.scala 276:73:@309.14]
  wire [31:0] _GEN_633; // @[Bus.scala 276:73:@309.14]
  wire [31:0] _GEN_634; // @[Bus.scala 276:73:@309.14]
  wire [31:0] _GEN_635; // @[Bus.scala 276:73:@309.14]
  wire [31:0] _GEN_636; // @[Bus.scala 276:73:@309.14]
  wire [31:0] _GEN_637; // @[Bus.scala 276:73:@309.14]
  wire [31:0] _GEN_638; // @[Bus.scala 276:73:@309.14]
  wire [31:0] _GEN_639; // @[Bus.scala 276:73:@309.14]
  wire [31:0] _GEN_640; // @[Bus.scala 276:73:@309.14]
  wire  _GEN_641; // @[Bus.scala 276:73:@309.14]
  wire  _GEN_642; // @[Bus.scala 276:73:@309.14]
  wire  _GEN_643; // @[Bus.scala 276:73:@309.14]
  wire  _GEN_644; // @[Bus.scala 276:73:@309.14]
  wire  _GEN_645; // @[Bus.scala 276:73:@309.14]
  wire  _GEN_646; // @[Bus.scala 276:73:@309.14]
  wire  _GEN_647; // @[Bus.scala 276:73:@309.14]
  wire  _GEN_648; // @[Bus.scala 276:73:@309.14]
  wire  _GEN_649; // @[Bus.scala 276:73:@309.14]
  wire  _GEN_650; // @[Bus.scala 276:73:@309.14]
  wire [3:0] _GEN_651; // @[Bus.scala 275:81:@308.12]
  wire [31:0] _GEN_652; // @[Bus.scala 275:81:@308.12]
  wire [31:0] _GEN_653; // @[Bus.scala 275:81:@308.12]
  wire [31:0] _GEN_654; // @[Bus.scala 275:81:@308.12]
  wire [31:0] _GEN_655; // @[Bus.scala 275:81:@308.12]
  wire [31:0] _GEN_656; // @[Bus.scala 275:81:@308.12]
  wire [31:0] _GEN_657; // @[Bus.scala 275:81:@308.12]
  wire [31:0] _GEN_658; // @[Bus.scala 275:81:@308.12]
  wire [31:0] _GEN_659; // @[Bus.scala 275:81:@308.12]
  wire  _GEN_660; // @[Bus.scala 275:81:@308.12]
  wire  _GEN_661; // @[Bus.scala 275:81:@308.12]
  wire  _GEN_662; // @[Bus.scala 275:81:@308.12]
  wire  _GEN_663; // @[Bus.scala 275:81:@308.12]
  wire  _GEN_664; // @[Bus.scala 275:81:@308.12]
  wire  _GEN_665; // @[Bus.scala 275:81:@308.12]
  wire  _GEN_666; // @[Bus.scala 275:81:@308.12]
  wire  _GEN_667; // @[Bus.scala 275:81:@308.12]
  wire  _GEN_668; // @[Bus.scala 275:81:@308.12]
  wire  _GEN_669; // @[Bus.scala 275:81:@308.12]
  wire [3:0] _GEN_670; // @[Bus.scala 274:73:@306.10]
  wire [31:0] _GEN_671; // @[Bus.scala 274:73:@306.10]
  wire [31:0] _GEN_672; // @[Bus.scala 274:73:@306.10]
  wire [31:0] _GEN_673; // @[Bus.scala 274:73:@306.10]
  wire [31:0] _GEN_674; // @[Bus.scala 274:73:@306.10]
  wire [31:0] _GEN_675; // @[Bus.scala 274:73:@306.10]
  wire [31:0] _GEN_676; // @[Bus.scala 274:73:@306.10]
  wire [31:0] _GEN_677; // @[Bus.scala 274:73:@306.10]
  wire [31:0] _GEN_678; // @[Bus.scala 274:73:@306.10]
  wire  _GEN_679; // @[Bus.scala 274:73:@306.10]
  wire  _GEN_680; // @[Bus.scala 274:73:@306.10]
  wire  _GEN_681; // @[Bus.scala 274:73:@306.10]
  wire  _GEN_682; // @[Bus.scala 274:73:@306.10]
  wire  _GEN_683; // @[Bus.scala 274:73:@306.10]
  wire  _GEN_684; // @[Bus.scala 274:73:@306.10]
  wire  _GEN_685; // @[Bus.scala 274:73:@306.10]
  wire  _GEN_686; // @[Bus.scala 274:73:@306.10]
  wire  _GEN_687; // @[Bus.scala 274:73:@306.10]
  wire  _GEN_688; // @[Bus.scala 274:73:@306.10]
  wire [3:0] _GEN_689; // @[Bus.scala 273:74:@304.8]
  wire [31:0] _GEN_690; // @[Bus.scala 273:74:@304.8]
  wire [31:0] _GEN_691; // @[Bus.scala 273:74:@304.8]
  wire [31:0] _GEN_692; // @[Bus.scala 273:74:@304.8]
  wire [31:0] _GEN_693; // @[Bus.scala 273:74:@304.8]
  wire [31:0] _GEN_694; // @[Bus.scala 273:74:@304.8]
  wire [31:0] _GEN_695; // @[Bus.scala 273:74:@304.8]
  wire [31:0] _GEN_696; // @[Bus.scala 273:74:@304.8]
  wire [31:0] _GEN_697; // @[Bus.scala 273:74:@304.8]
  wire  _GEN_698; // @[Bus.scala 273:74:@304.8]
  wire  _GEN_699; // @[Bus.scala 273:74:@304.8]
  wire  _GEN_700; // @[Bus.scala 273:74:@304.8]
  wire  _GEN_701; // @[Bus.scala 273:74:@304.8]
  wire  _GEN_702; // @[Bus.scala 273:74:@304.8]
  wire  _GEN_703; // @[Bus.scala 273:74:@304.8]
  wire  _GEN_704; // @[Bus.scala 273:74:@304.8]
  wire  _GEN_705; // @[Bus.scala 273:74:@304.8]
  wire  _GEN_706; // @[Bus.scala 273:74:@304.8]
  wire  _GEN_707; // @[Bus.scala 273:74:@304.8]
  wire [3:0] _GEN_708; // @[Bus.scala 272:41:@301.6]
  wire [31:0] _GEN_709; // @[Bus.scala 272:41:@301.6]
  wire [31:0] _GEN_710; // @[Bus.scala 272:41:@301.6]
  wire [31:0] _GEN_711; // @[Bus.scala 272:41:@301.6]
  wire [31:0] _GEN_712; // @[Bus.scala 272:41:@301.6]
  wire [31:0] _GEN_713; // @[Bus.scala 272:41:@301.6]
  wire [31:0] _GEN_714; // @[Bus.scala 272:41:@301.6]
  wire [31:0] _GEN_715; // @[Bus.scala 272:41:@301.6]
  wire [31:0] _GEN_716; // @[Bus.scala 272:41:@301.6]
  wire  _GEN_717; // @[Bus.scala 272:41:@301.6]
  wire  _GEN_718; // @[Bus.scala 272:41:@301.6]
  wire  _GEN_719; // @[Bus.scala 272:41:@301.6]
  wire  _GEN_720; // @[Bus.scala 272:41:@301.6]
  wire  _GEN_721; // @[Bus.scala 272:41:@301.6]
  wire  _GEN_722; // @[Bus.scala 272:41:@301.6]
  wire  _GEN_723; // @[Bus.scala 272:41:@301.6]
  wire  _GEN_724; // @[Bus.scala 272:41:@301.6]
  wire  _GEN_725; // @[Bus.scala 272:41:@301.6]
  wire  _GEN_726; // @[Bus.scala 272:41:@301.6]
  wire [3:0] _GEN_727; // @[Bus.scala 305:73:@348.14]
  wire [31:0] _GEN_728; // @[Bus.scala 305:73:@348.14]
  wire [31:0] _GEN_729; // @[Bus.scala 305:73:@348.14]
  wire [31:0] _GEN_730; // @[Bus.scala 305:73:@348.14]
  wire [31:0] _GEN_731; // @[Bus.scala 305:73:@348.14]
  wire [31:0] _GEN_732; // @[Bus.scala 305:73:@348.14]
  wire [31:0] _GEN_733; // @[Bus.scala 305:73:@348.14]
  wire [31:0] _GEN_734; // @[Bus.scala 305:73:@348.14]
  wire [31:0] _GEN_735; // @[Bus.scala 305:73:@348.14]
  wire  _GEN_736; // @[Bus.scala 305:73:@348.14]
  wire  _GEN_737; // @[Bus.scala 305:73:@348.14]
  wire  _GEN_738; // @[Bus.scala 305:73:@348.14]
  wire  _GEN_739; // @[Bus.scala 305:73:@348.14]
  wire  _GEN_740; // @[Bus.scala 305:73:@348.14]
  wire  _GEN_741; // @[Bus.scala 305:73:@348.14]
  wire  _GEN_742; // @[Bus.scala 305:73:@348.14]
  wire  _GEN_743; // @[Bus.scala 305:73:@348.14]
  wire  _GEN_744; // @[Bus.scala 305:73:@348.14]
  wire  _GEN_745; // @[Bus.scala 305:73:@348.14]
  wire [3:0] _GEN_746; // @[Bus.scala 304:81:@347.12]
  wire [31:0] _GEN_747; // @[Bus.scala 304:81:@347.12]
  wire [31:0] _GEN_748; // @[Bus.scala 304:81:@347.12]
  wire [31:0] _GEN_749; // @[Bus.scala 304:81:@347.12]
  wire [31:0] _GEN_750; // @[Bus.scala 304:81:@347.12]
  wire [31:0] _GEN_751; // @[Bus.scala 304:81:@347.12]
  wire [31:0] _GEN_752; // @[Bus.scala 304:81:@347.12]
  wire [31:0] _GEN_753; // @[Bus.scala 304:81:@347.12]
  wire [31:0] _GEN_754; // @[Bus.scala 304:81:@347.12]
  wire  _GEN_755; // @[Bus.scala 304:81:@347.12]
  wire  _GEN_756; // @[Bus.scala 304:81:@347.12]
  wire  _GEN_757; // @[Bus.scala 304:81:@347.12]
  wire  _GEN_758; // @[Bus.scala 304:81:@347.12]
  wire  _GEN_759; // @[Bus.scala 304:81:@347.12]
  wire  _GEN_760; // @[Bus.scala 304:81:@347.12]
  wire  _GEN_761; // @[Bus.scala 304:81:@347.12]
  wire  _GEN_762; // @[Bus.scala 304:81:@347.12]
  wire  _GEN_763; // @[Bus.scala 304:81:@347.12]
  wire  _GEN_764; // @[Bus.scala 304:81:@347.12]
  wire [3:0] _GEN_765; // @[Bus.scala 303:73:@345.10]
  wire [31:0] _GEN_766; // @[Bus.scala 303:73:@345.10]
  wire [31:0] _GEN_767; // @[Bus.scala 303:73:@345.10]
  wire [31:0] _GEN_768; // @[Bus.scala 303:73:@345.10]
  wire [31:0] _GEN_769; // @[Bus.scala 303:73:@345.10]
  wire [31:0] _GEN_770; // @[Bus.scala 303:73:@345.10]
  wire [31:0] _GEN_771; // @[Bus.scala 303:73:@345.10]
  wire [31:0] _GEN_772; // @[Bus.scala 303:73:@345.10]
  wire [31:0] _GEN_773; // @[Bus.scala 303:73:@345.10]
  wire  _GEN_774; // @[Bus.scala 303:73:@345.10]
  wire  _GEN_775; // @[Bus.scala 303:73:@345.10]
  wire  _GEN_776; // @[Bus.scala 303:73:@345.10]
  wire  _GEN_777; // @[Bus.scala 303:73:@345.10]
  wire  _GEN_778; // @[Bus.scala 303:73:@345.10]
  wire  _GEN_779; // @[Bus.scala 303:73:@345.10]
  wire  _GEN_780; // @[Bus.scala 303:73:@345.10]
  wire  _GEN_781; // @[Bus.scala 303:73:@345.10]
  wire  _GEN_782; // @[Bus.scala 303:73:@345.10]
  wire  _GEN_783; // @[Bus.scala 303:73:@345.10]
  wire [3:0] _GEN_784; // @[Bus.scala 302:73:@343.8]
  wire [31:0] _GEN_785; // @[Bus.scala 302:73:@343.8]
  wire [31:0] _GEN_786; // @[Bus.scala 302:73:@343.8]
  wire [31:0] _GEN_787; // @[Bus.scala 302:73:@343.8]
  wire [31:0] _GEN_788; // @[Bus.scala 302:73:@343.8]
  wire [31:0] _GEN_789; // @[Bus.scala 302:73:@343.8]
  wire [31:0] _GEN_790; // @[Bus.scala 302:73:@343.8]
  wire [31:0] _GEN_791; // @[Bus.scala 302:73:@343.8]
  wire [31:0] _GEN_792; // @[Bus.scala 302:73:@343.8]
  wire  _GEN_793; // @[Bus.scala 302:73:@343.8]
  wire  _GEN_794; // @[Bus.scala 302:73:@343.8]
  wire  _GEN_795; // @[Bus.scala 302:73:@343.8]
  wire  _GEN_796; // @[Bus.scala 302:73:@343.8]
  wire  _GEN_797; // @[Bus.scala 302:73:@343.8]
  wire  _GEN_798; // @[Bus.scala 302:73:@343.8]
  wire  _GEN_799; // @[Bus.scala 302:73:@343.8]
  wire  _GEN_800; // @[Bus.scala 302:73:@343.8]
  wire  _GEN_801; // @[Bus.scala 302:73:@343.8]
  wire  _GEN_802; // @[Bus.scala 302:73:@343.8]
  wire [3:0] _GEN_803; // @[Bus.scala 301:41:@341.6]
  wire [31:0] _GEN_804; // @[Bus.scala 301:41:@341.6]
  wire [31:0] _GEN_805; // @[Bus.scala 301:41:@341.6]
  wire [31:0] _GEN_806; // @[Bus.scala 301:41:@341.6]
  wire [31:0] _GEN_807; // @[Bus.scala 301:41:@341.6]
  wire [31:0] _GEN_808; // @[Bus.scala 301:41:@341.6]
  wire [31:0] _GEN_809; // @[Bus.scala 301:41:@341.6]
  wire [31:0] _GEN_810; // @[Bus.scala 301:41:@341.6]
  wire [31:0] _GEN_811; // @[Bus.scala 301:41:@341.6]
  wire  _GEN_812; // @[Bus.scala 301:41:@341.6]
  wire  _GEN_813; // @[Bus.scala 301:41:@341.6]
  wire  _GEN_814; // @[Bus.scala 301:41:@341.6]
  wire  _GEN_815; // @[Bus.scala 301:41:@341.6]
  wire  _GEN_816; // @[Bus.scala 301:41:@341.6]
  wire  _GEN_817; // @[Bus.scala 301:41:@341.6]
  wire  _GEN_818; // @[Bus.scala 301:41:@341.6]
  wire  _GEN_819; // @[Bus.scala 301:41:@341.6]
  wire  _GEN_820; // @[Bus.scala 301:41:@341.6]
  wire  _GEN_821; // @[Bus.scala 301:41:@341.6]
  wire  _T_345; // @[Bus.scala 333:65:@386.12]
  wire [32:0] _T_347; // @[Bus.scala 336:93:@390.16]
  wire [31:0] _T_348; // @[Bus.scala 336:93:@391.16]
  wire [31:0] _T_349; // @[Bus.scala 336:93:@392.16]
  wire [3:0] _GEN_822; // @[Bus.scala 334:73:@388.14]
  wire [31:0] _GEN_823; // @[Bus.scala 334:73:@388.14]
  wire [31:0] _GEN_824; // @[Bus.scala 334:73:@388.14]
  wire [31:0] _GEN_825; // @[Bus.scala 334:73:@388.14]
  wire [31:0] _GEN_826; // @[Bus.scala 334:73:@388.14]
  wire [31:0] _GEN_827; // @[Bus.scala 334:73:@388.14]
  wire [31:0] _GEN_828; // @[Bus.scala 334:73:@388.14]
  wire [31:0] _GEN_829; // @[Bus.scala 334:73:@388.14]
  wire [31:0] _GEN_830; // @[Bus.scala 334:73:@388.14]
  wire  _GEN_831; // @[Bus.scala 334:73:@388.14]
  wire  _GEN_832; // @[Bus.scala 334:73:@388.14]
  wire  _GEN_833; // @[Bus.scala 334:73:@388.14]
  wire  _GEN_834; // @[Bus.scala 334:73:@388.14]
  wire  _GEN_835; // @[Bus.scala 334:73:@388.14]
  wire  _GEN_836; // @[Bus.scala 334:73:@388.14]
  wire  _GEN_837; // @[Bus.scala 334:73:@388.14]
  wire  _GEN_838; // @[Bus.scala 334:73:@388.14]
  wire  _GEN_839; // @[Bus.scala 334:73:@388.14]
  wire  _GEN_840; // @[Bus.scala 334:73:@388.14]
  wire [3:0] _GEN_841; // @[Bus.scala 333:81:@387.12]
  wire [31:0] _GEN_842; // @[Bus.scala 333:81:@387.12]
  wire [31:0] _GEN_843; // @[Bus.scala 333:81:@387.12]
  wire [31:0] _GEN_844; // @[Bus.scala 333:81:@387.12]
  wire [31:0] _GEN_845; // @[Bus.scala 333:81:@387.12]
  wire [31:0] _GEN_846; // @[Bus.scala 333:81:@387.12]
  wire [31:0] _GEN_847; // @[Bus.scala 333:81:@387.12]
  wire [31:0] _GEN_848; // @[Bus.scala 333:81:@387.12]
  wire [31:0] _GEN_849; // @[Bus.scala 333:81:@387.12]
  wire  _GEN_850; // @[Bus.scala 333:81:@387.12]
  wire  _GEN_851; // @[Bus.scala 333:81:@387.12]
  wire  _GEN_852; // @[Bus.scala 333:81:@387.12]
  wire  _GEN_853; // @[Bus.scala 333:81:@387.12]
  wire  _GEN_854; // @[Bus.scala 333:81:@387.12]
  wire  _GEN_855; // @[Bus.scala 333:81:@387.12]
  wire  _GEN_856; // @[Bus.scala 333:81:@387.12]
  wire  _GEN_857; // @[Bus.scala 333:81:@387.12]
  wire  _GEN_858; // @[Bus.scala 333:81:@387.12]
  wire  _GEN_859; // @[Bus.scala 333:81:@387.12]
  wire [3:0] _GEN_860; // @[Bus.scala 332:73:@385.10]
  wire [31:0] _GEN_861; // @[Bus.scala 332:73:@385.10]
  wire [31:0] _GEN_862; // @[Bus.scala 332:73:@385.10]
  wire [31:0] _GEN_863; // @[Bus.scala 332:73:@385.10]
  wire [31:0] _GEN_864; // @[Bus.scala 332:73:@385.10]
  wire [31:0] _GEN_865; // @[Bus.scala 332:73:@385.10]
  wire [31:0] _GEN_866; // @[Bus.scala 332:73:@385.10]
  wire [31:0] _GEN_867; // @[Bus.scala 332:73:@385.10]
  wire [31:0] _GEN_868; // @[Bus.scala 332:73:@385.10]
  wire  _GEN_869; // @[Bus.scala 332:73:@385.10]
  wire  _GEN_870; // @[Bus.scala 332:73:@385.10]
  wire  _GEN_871; // @[Bus.scala 332:73:@385.10]
  wire  _GEN_872; // @[Bus.scala 332:73:@385.10]
  wire  _GEN_873; // @[Bus.scala 332:73:@385.10]
  wire  _GEN_874; // @[Bus.scala 332:73:@385.10]
  wire  _GEN_875; // @[Bus.scala 332:73:@385.10]
  wire  _GEN_876; // @[Bus.scala 332:73:@385.10]
  wire  _GEN_877; // @[Bus.scala 332:73:@385.10]
  wire  _GEN_878; // @[Bus.scala 332:73:@385.10]
  wire [3:0] _GEN_879; // @[Bus.scala 331:74:@383.8]
  wire [31:0] _GEN_880; // @[Bus.scala 331:74:@383.8]
  wire [31:0] _GEN_881; // @[Bus.scala 331:74:@383.8]
  wire [31:0] _GEN_882; // @[Bus.scala 331:74:@383.8]
  wire [31:0] _GEN_883; // @[Bus.scala 331:74:@383.8]
  wire [31:0] _GEN_884; // @[Bus.scala 331:74:@383.8]
  wire [31:0] _GEN_885; // @[Bus.scala 331:74:@383.8]
  wire [31:0] _GEN_886; // @[Bus.scala 331:74:@383.8]
  wire [31:0] _GEN_887; // @[Bus.scala 331:74:@383.8]
  wire  _GEN_888; // @[Bus.scala 331:74:@383.8]
  wire  _GEN_889; // @[Bus.scala 331:74:@383.8]
  wire  _GEN_890; // @[Bus.scala 331:74:@383.8]
  wire  _GEN_891; // @[Bus.scala 331:74:@383.8]
  wire  _GEN_892; // @[Bus.scala 331:74:@383.8]
  wire  _GEN_893; // @[Bus.scala 331:74:@383.8]
  wire  _GEN_894; // @[Bus.scala 331:74:@383.8]
  wire  _GEN_895; // @[Bus.scala 331:74:@383.8]
  wire  _GEN_896; // @[Bus.scala 331:74:@383.8]
  wire  _GEN_897; // @[Bus.scala 331:74:@383.8]
  wire [3:0] _GEN_898; // @[Bus.scala 330:41:@380.6]
  wire [31:0] _GEN_899; // @[Bus.scala 330:41:@380.6]
  wire [31:0] _GEN_900; // @[Bus.scala 330:41:@380.6]
  wire [31:0] _GEN_901; // @[Bus.scala 330:41:@380.6]
  wire [31:0] _GEN_902; // @[Bus.scala 330:41:@380.6]
  wire [31:0] _GEN_903; // @[Bus.scala 330:41:@380.6]
  wire [31:0] _GEN_904; // @[Bus.scala 330:41:@380.6]
  wire [31:0] _GEN_905; // @[Bus.scala 330:41:@380.6]
  wire [31:0] _GEN_906; // @[Bus.scala 330:41:@380.6]
  wire  _GEN_907; // @[Bus.scala 330:41:@380.6]
  wire  _GEN_908; // @[Bus.scala 330:41:@380.6]
  wire  _GEN_909; // @[Bus.scala 330:41:@380.6]
  wire  _GEN_910; // @[Bus.scala 330:41:@380.6]
  wire  _GEN_911; // @[Bus.scala 330:41:@380.6]
  wire  _GEN_912; // @[Bus.scala 330:41:@380.6]
  wire  _GEN_913; // @[Bus.scala 330:41:@380.6]
  wire  _GEN_914; // @[Bus.scala 330:41:@380.6]
  wire  _GEN_915; // @[Bus.scala 330:41:@380.6]
  wire  _GEN_916; // @[Bus.scala 330:41:@380.6]
  wire [3:0] _GEN_917; // @[Bus.scala 363:73:@427.14]
  wire [31:0] _GEN_918; // @[Bus.scala 363:73:@427.14]
  wire [31:0] _GEN_919; // @[Bus.scala 363:73:@427.14]
  wire [31:0] _GEN_920; // @[Bus.scala 363:73:@427.14]
  wire [31:0] _GEN_921; // @[Bus.scala 363:73:@427.14]
  wire [31:0] _GEN_922; // @[Bus.scala 363:73:@427.14]
  wire [31:0] _GEN_923; // @[Bus.scala 363:73:@427.14]
  wire [31:0] _GEN_924; // @[Bus.scala 363:73:@427.14]
  wire [31:0] _GEN_925; // @[Bus.scala 363:73:@427.14]
  wire  _GEN_926; // @[Bus.scala 363:73:@427.14]
  wire  _GEN_927; // @[Bus.scala 363:73:@427.14]
  wire  _GEN_928; // @[Bus.scala 363:73:@427.14]
  wire  _GEN_929; // @[Bus.scala 363:73:@427.14]
  wire  _GEN_930; // @[Bus.scala 363:73:@427.14]
  wire  _GEN_931; // @[Bus.scala 363:73:@427.14]
  wire  _GEN_932; // @[Bus.scala 363:73:@427.14]
  wire  _GEN_933; // @[Bus.scala 363:73:@427.14]
  wire  _GEN_934; // @[Bus.scala 363:73:@427.14]
  wire  _GEN_935; // @[Bus.scala 363:73:@427.14]
  wire [3:0] _GEN_936; // @[Bus.scala 362:81:@426.12]
  wire [31:0] _GEN_937; // @[Bus.scala 362:81:@426.12]
  wire [31:0] _GEN_938; // @[Bus.scala 362:81:@426.12]
  wire [31:0] _GEN_939; // @[Bus.scala 362:81:@426.12]
  wire [31:0] _GEN_940; // @[Bus.scala 362:81:@426.12]
  wire [31:0] _GEN_941; // @[Bus.scala 362:81:@426.12]
  wire [31:0] _GEN_942; // @[Bus.scala 362:81:@426.12]
  wire [31:0] _GEN_943; // @[Bus.scala 362:81:@426.12]
  wire [31:0] _GEN_944; // @[Bus.scala 362:81:@426.12]
  wire  _GEN_945; // @[Bus.scala 362:81:@426.12]
  wire  _GEN_946; // @[Bus.scala 362:81:@426.12]
  wire  _GEN_947; // @[Bus.scala 362:81:@426.12]
  wire  _GEN_948; // @[Bus.scala 362:81:@426.12]
  wire  _GEN_949; // @[Bus.scala 362:81:@426.12]
  wire  _GEN_950; // @[Bus.scala 362:81:@426.12]
  wire  _GEN_951; // @[Bus.scala 362:81:@426.12]
  wire  _GEN_952; // @[Bus.scala 362:81:@426.12]
  wire  _GEN_953; // @[Bus.scala 362:81:@426.12]
  wire  _GEN_954; // @[Bus.scala 362:81:@426.12]
  wire [3:0] _GEN_955; // @[Bus.scala 361:73:@424.10]
  wire [31:0] _GEN_956; // @[Bus.scala 361:73:@424.10]
  wire [31:0] _GEN_957; // @[Bus.scala 361:73:@424.10]
  wire [31:0] _GEN_958; // @[Bus.scala 361:73:@424.10]
  wire [31:0] _GEN_959; // @[Bus.scala 361:73:@424.10]
  wire [31:0] _GEN_960; // @[Bus.scala 361:73:@424.10]
  wire [31:0] _GEN_961; // @[Bus.scala 361:73:@424.10]
  wire [31:0] _GEN_962; // @[Bus.scala 361:73:@424.10]
  wire [31:0] _GEN_963; // @[Bus.scala 361:73:@424.10]
  wire  _GEN_964; // @[Bus.scala 361:73:@424.10]
  wire  _GEN_965; // @[Bus.scala 361:73:@424.10]
  wire  _GEN_966; // @[Bus.scala 361:73:@424.10]
  wire  _GEN_967; // @[Bus.scala 361:73:@424.10]
  wire  _GEN_968; // @[Bus.scala 361:73:@424.10]
  wire  _GEN_969; // @[Bus.scala 361:73:@424.10]
  wire  _GEN_970; // @[Bus.scala 361:73:@424.10]
  wire  _GEN_971; // @[Bus.scala 361:73:@424.10]
  wire  _GEN_972; // @[Bus.scala 361:73:@424.10]
  wire  _GEN_973; // @[Bus.scala 361:73:@424.10]
  wire [3:0] _GEN_974; // @[Bus.scala 360:73:@422.8]
  wire [31:0] _GEN_975; // @[Bus.scala 360:73:@422.8]
  wire [31:0] _GEN_976; // @[Bus.scala 360:73:@422.8]
  wire [31:0] _GEN_977; // @[Bus.scala 360:73:@422.8]
  wire [31:0] _GEN_978; // @[Bus.scala 360:73:@422.8]
  wire [31:0] _GEN_979; // @[Bus.scala 360:73:@422.8]
  wire [31:0] _GEN_980; // @[Bus.scala 360:73:@422.8]
  wire [31:0] _GEN_981; // @[Bus.scala 360:73:@422.8]
  wire [31:0] _GEN_982; // @[Bus.scala 360:73:@422.8]
  wire  _GEN_983; // @[Bus.scala 360:73:@422.8]
  wire  _GEN_984; // @[Bus.scala 360:73:@422.8]
  wire  _GEN_985; // @[Bus.scala 360:73:@422.8]
  wire  _GEN_986; // @[Bus.scala 360:73:@422.8]
  wire  _GEN_987; // @[Bus.scala 360:73:@422.8]
  wire  _GEN_988; // @[Bus.scala 360:73:@422.8]
  wire  _GEN_989; // @[Bus.scala 360:73:@422.8]
  wire  _GEN_990; // @[Bus.scala 360:73:@422.8]
  wire  _GEN_991; // @[Bus.scala 360:73:@422.8]
  wire  _GEN_992; // @[Bus.scala 360:73:@422.8]
  wire [3:0] _GEN_993; // @[Bus.scala 359:41:@420.6]
  wire [31:0] _GEN_994; // @[Bus.scala 359:41:@420.6]
  wire [31:0] _GEN_995; // @[Bus.scala 359:41:@420.6]
  wire [31:0] _GEN_996; // @[Bus.scala 359:41:@420.6]
  wire [31:0] _GEN_997; // @[Bus.scala 359:41:@420.6]
  wire [31:0] _GEN_998; // @[Bus.scala 359:41:@420.6]
  wire [31:0] _GEN_999; // @[Bus.scala 359:41:@420.6]
  wire [31:0] _GEN_1000; // @[Bus.scala 359:41:@420.6]
  wire [31:0] _GEN_1001; // @[Bus.scala 359:41:@420.6]
  wire  _GEN_1002; // @[Bus.scala 359:41:@420.6]
  wire  _GEN_1003; // @[Bus.scala 359:41:@420.6]
  wire  _GEN_1004; // @[Bus.scala 359:41:@420.6]
  wire  _GEN_1005; // @[Bus.scala 359:41:@420.6]
  wire  _GEN_1006; // @[Bus.scala 359:41:@420.6]
  wire  _GEN_1007; // @[Bus.scala 359:41:@420.6]
  wire  _GEN_1008; // @[Bus.scala 359:41:@420.6]
  wire  _GEN_1009; // @[Bus.scala 359:41:@420.6]
  wire  _GEN_1010; // @[Bus.scala 359:41:@420.6]
  wire  _GEN_1011; // @[Bus.scala 359:41:@420.6]
  wire  _T_390; // @[Bus.scala 388:30:@458.6]
  wire [3:0] _GEN_1012; // @[Bus.scala 389:50:@460.8]
  wire [31:0] _GEN_1013; // @[Bus.scala 389:50:@460.8]
  wire [31:0] _GEN_1014; // @[Bus.scala 389:50:@460.8]
  wire [31:0] _GEN_1015; // @[Bus.scala 389:50:@460.8]
  wire [31:0] _GEN_1016; // @[Bus.scala 389:50:@460.8]
  wire [31:0] _GEN_1017; // @[Bus.scala 389:50:@460.8]
  wire  _GEN_1018; // @[Bus.scala 389:50:@460.8]
  wire  _GEN_1019; // @[Bus.scala 389:50:@460.8]
  wire  _GEN_1020; // @[Bus.scala 389:50:@460.8]
  wire  _GEN_1021; // @[Bus.scala 389:50:@460.8]
  wire  _GEN_1022; // @[Bus.scala 389:50:@460.8]
  wire  _GEN_1023; // @[Bus.scala 389:50:@460.8]
  wire  _GEN_1024; // @[Bus.scala 389:50:@460.8]
  wire  _GEN_1025; // @[Bus.scala 389:50:@460.8]
  wire  _GEN_1026; // @[Bus.scala 389:50:@460.8]
  wire  _GEN_1027; // @[Bus.scala 389:50:@460.8]
  wire [3:0] _GEN_1028; // @[Bus.scala 388:41:@459.6]
  wire [31:0] _GEN_1029; // @[Bus.scala 388:41:@459.6]
  wire [31:0] _GEN_1030; // @[Bus.scala 388:41:@459.6]
  wire [31:0] _GEN_1031; // @[Bus.scala 388:41:@459.6]
  wire [31:0] _GEN_1032; // @[Bus.scala 388:41:@459.6]
  wire [31:0] _GEN_1033; // @[Bus.scala 388:41:@459.6]
  wire  _GEN_1034; // @[Bus.scala 388:41:@459.6]
  wire  _GEN_1035; // @[Bus.scala 388:41:@459.6]
  wire  _GEN_1036; // @[Bus.scala 388:41:@459.6]
  wire  _GEN_1037; // @[Bus.scala 388:41:@459.6]
  wire  _GEN_1038; // @[Bus.scala 388:41:@459.6]
  wire  _GEN_1039; // @[Bus.scala 388:41:@459.6]
  wire  _GEN_1040; // @[Bus.scala 388:41:@459.6]
  wire  _GEN_1041; // @[Bus.scala 388:41:@459.6]
  wire  _GEN_1042; // @[Bus.scala 388:41:@459.6]
  wire  _GEN_1043; // @[Bus.scala 388:41:@459.6]
  wire  _T_401; // @[Bus.scala 408:30:@479.6]
  wire  _T_402; // @[Bus.scala 409:45:@481.8]
  wire  _T_404; // @[Bus.scala 409:30:@482.8]
  wire [3:0] _GEN_1044; // @[Bus.scala 410:57:@484.10]
  wire [31:0] _GEN_1045; // @[Bus.scala 410:57:@484.10]
  wire [31:0] _GEN_1046; // @[Bus.scala 410:57:@484.10]
  wire [31:0] _GEN_1047; // @[Bus.scala 410:57:@484.10]
  wire [31:0] _GEN_1048; // @[Bus.scala 410:57:@484.10]
  wire [31:0] _GEN_1049; // @[Bus.scala 410:57:@484.10]
  wire [31:0] _GEN_1050; // @[Bus.scala 410:57:@484.10]
  wire [31:0] _GEN_1051; // @[Bus.scala 410:57:@484.10]
  wire  _GEN_1052; // @[Bus.scala 410:57:@484.10]
  wire  _GEN_1053; // @[Bus.scala 410:57:@484.10]
  wire  _GEN_1054; // @[Bus.scala 410:57:@484.10]
  wire  _GEN_1055; // @[Bus.scala 410:57:@484.10]
  wire  _GEN_1056; // @[Bus.scala 410:57:@484.10]
  wire  _GEN_1057; // @[Bus.scala 410:57:@484.10]
  wire  _GEN_1058; // @[Bus.scala 410:57:@484.10]
  wire  _GEN_1059; // @[Bus.scala 410:57:@484.10]
  wire  _GEN_1060; // @[Bus.scala 410:57:@484.10]
  wire  _GEN_1061; // @[Bus.scala 410:57:@484.10]
  wire [3:0] _GEN_1062; // @[Bus.scala 409:75:@483.8]
  wire [31:0] _GEN_1063; // @[Bus.scala 409:75:@483.8]
  wire [31:0] _GEN_1064; // @[Bus.scala 409:75:@483.8]
  wire [31:0] _GEN_1065; // @[Bus.scala 409:75:@483.8]
  wire [31:0] _GEN_1066; // @[Bus.scala 409:75:@483.8]
  wire [31:0] _GEN_1067; // @[Bus.scala 409:75:@483.8]
  wire [31:0] _GEN_1068; // @[Bus.scala 409:75:@483.8]
  wire [31:0] _GEN_1069; // @[Bus.scala 409:75:@483.8]
  wire  _GEN_1070; // @[Bus.scala 409:75:@483.8]
  wire  _GEN_1071; // @[Bus.scala 409:75:@483.8]
  wire  _GEN_1072; // @[Bus.scala 409:75:@483.8]
  wire  _GEN_1073; // @[Bus.scala 409:75:@483.8]
  wire  _GEN_1074; // @[Bus.scala 409:75:@483.8]
  wire  _GEN_1075; // @[Bus.scala 409:75:@483.8]
  wire  _GEN_1076; // @[Bus.scala 409:75:@483.8]
  wire  _GEN_1077; // @[Bus.scala 409:75:@483.8]
  wire  _GEN_1078; // @[Bus.scala 409:75:@483.8]
  wire  _GEN_1079; // @[Bus.scala 409:75:@483.8]
  wire [3:0] _GEN_1080; // @[Bus.scala 408:41:@480.6]
  wire [31:0] _GEN_1081; // @[Bus.scala 408:41:@480.6]
  wire [31:0] _GEN_1082; // @[Bus.scala 408:41:@480.6]
  wire [31:0] _GEN_1083; // @[Bus.scala 408:41:@480.6]
  wire [31:0] _GEN_1084; // @[Bus.scala 408:41:@480.6]
  wire [31:0] _GEN_1085; // @[Bus.scala 408:41:@480.6]
  wire [31:0] _GEN_1086; // @[Bus.scala 408:41:@480.6]
  wire [31:0] _GEN_1087; // @[Bus.scala 408:41:@480.6]
  wire  _GEN_1088; // @[Bus.scala 408:41:@480.6]
  wire  _GEN_1089; // @[Bus.scala 408:41:@480.6]
  wire  _GEN_1090; // @[Bus.scala 408:41:@480.6]
  wire  _GEN_1091; // @[Bus.scala 408:41:@480.6]
  wire  _GEN_1092; // @[Bus.scala 408:41:@480.6]
  wire  _GEN_1093; // @[Bus.scala 408:41:@480.6]
  wire  _GEN_1094; // @[Bus.scala 408:41:@480.6]
  wire  _GEN_1095; // @[Bus.scala 408:41:@480.6]
  wire  _GEN_1096; // @[Bus.scala 408:41:@480.6]
  wire  _GEN_1097; // @[Bus.scala 408:41:@480.6]
  wire [3:0] _GEN_1098; // @[Bus.scala 434:57:@510.10]
  wire [31:0] _GEN_1099; // @[Bus.scala 434:57:@510.10]
  wire [31:0] _GEN_1100; // @[Bus.scala 434:57:@510.10]
  wire [31:0] _GEN_1101; // @[Bus.scala 434:57:@510.10]
  wire [31:0] _GEN_1102; // @[Bus.scala 434:57:@510.10]
  wire [31:0] _GEN_1103; // @[Bus.scala 434:57:@510.10]
  wire [31:0] _GEN_1104; // @[Bus.scala 434:57:@510.10]
  wire [31:0] _GEN_1105; // @[Bus.scala 434:57:@510.10]
  wire  _GEN_1106; // @[Bus.scala 434:57:@510.10]
  wire  _GEN_1107; // @[Bus.scala 434:57:@510.10]
  wire  _GEN_1108; // @[Bus.scala 434:57:@510.10]
  wire  _GEN_1109; // @[Bus.scala 434:57:@510.10]
  wire  _GEN_1110; // @[Bus.scala 434:57:@510.10]
  wire  _GEN_1111; // @[Bus.scala 434:57:@510.10]
  wire  _GEN_1112; // @[Bus.scala 434:57:@510.10]
  wire  _GEN_1113; // @[Bus.scala 434:57:@510.10]
  wire  _GEN_1114; // @[Bus.scala 434:57:@510.10]
  wire  _GEN_1115; // @[Bus.scala 434:57:@510.10]
  wire [3:0] _GEN_1116; // @[Bus.scala 433:74:@509.8]
  wire [31:0] _GEN_1117; // @[Bus.scala 433:74:@509.8]
  wire [31:0] _GEN_1118; // @[Bus.scala 433:74:@509.8]
  wire [31:0] _GEN_1119; // @[Bus.scala 433:74:@509.8]
  wire [31:0] _GEN_1120; // @[Bus.scala 433:74:@509.8]
  wire [31:0] _GEN_1121; // @[Bus.scala 433:74:@509.8]
  wire [31:0] _GEN_1122; // @[Bus.scala 433:74:@509.8]
  wire [31:0] _GEN_1123; // @[Bus.scala 433:74:@509.8]
  wire  _GEN_1124; // @[Bus.scala 433:74:@509.8]
  wire  _GEN_1125; // @[Bus.scala 433:74:@509.8]
  wire  _GEN_1126; // @[Bus.scala 433:74:@509.8]
  wire  _GEN_1127; // @[Bus.scala 433:74:@509.8]
  wire  _GEN_1128; // @[Bus.scala 433:74:@509.8]
  wire  _GEN_1129; // @[Bus.scala 433:74:@509.8]
  wire  _GEN_1130; // @[Bus.scala 433:74:@509.8]
  wire  _GEN_1131; // @[Bus.scala 433:74:@509.8]
  wire  _GEN_1132; // @[Bus.scala 433:74:@509.8]
  wire  _GEN_1133; // @[Bus.scala 433:74:@509.8]
  wire [3:0] _GEN_1134; // @[Bus.scala 432:41:@507.6]
  wire [31:0] _GEN_1135; // @[Bus.scala 432:41:@507.6]
  wire [31:0] _GEN_1136; // @[Bus.scala 432:41:@507.6]
  wire [31:0] _GEN_1137; // @[Bus.scala 432:41:@507.6]
  wire [31:0] _GEN_1138; // @[Bus.scala 432:41:@507.6]
  wire [31:0] _GEN_1139; // @[Bus.scala 432:41:@507.6]
  wire [31:0] _GEN_1140; // @[Bus.scala 432:41:@507.6]
  wire [31:0] _GEN_1141; // @[Bus.scala 432:41:@507.6]
  wire  _GEN_1142; // @[Bus.scala 432:41:@507.6]
  wire  _GEN_1143; // @[Bus.scala 432:41:@507.6]
  wire  _GEN_1144; // @[Bus.scala 432:41:@507.6]
  wire  _GEN_1145; // @[Bus.scala 432:41:@507.6]
  wire  _GEN_1146; // @[Bus.scala 432:41:@507.6]
  wire  _GEN_1147; // @[Bus.scala 432:41:@507.6]
  wire  _GEN_1148; // @[Bus.scala 432:41:@507.6]
  wire  _GEN_1149; // @[Bus.scala 432:41:@507.6]
  wire  _GEN_1150; // @[Bus.scala 432:41:@507.6]
  wire  _GEN_1151; // @[Bus.scala 432:41:@507.6]
  wire  _T_429; // @[Bus.scala 456:30:@532.6]
  wire [3:0] _GEN_1152; // @[Bus.scala 457:50:@534.8]
  wire [31:0] _GEN_1153; // @[Bus.scala 457:50:@534.8]
  wire [31:0] _GEN_1154; // @[Bus.scala 457:50:@534.8]
  wire [31:0] _GEN_1155; // @[Bus.scala 457:50:@534.8]
  wire [31:0] _GEN_1156; // @[Bus.scala 457:50:@534.8]
  wire [31:0] _GEN_1157; // @[Bus.scala 457:50:@534.8]
  wire  _GEN_1158; // @[Bus.scala 457:50:@534.8]
  wire  _GEN_1159; // @[Bus.scala 457:50:@534.8]
  wire  _GEN_1160; // @[Bus.scala 457:50:@534.8]
  wire  _GEN_1161; // @[Bus.scala 457:50:@534.8]
  wire  _GEN_1162; // @[Bus.scala 457:50:@534.8]
  wire  _GEN_1163; // @[Bus.scala 457:50:@534.8]
  wire  _GEN_1164; // @[Bus.scala 457:50:@534.8]
  wire  _GEN_1165; // @[Bus.scala 457:50:@534.8]
  wire  _GEN_1166; // @[Bus.scala 457:50:@534.8]
  wire  _GEN_1167; // @[Bus.scala 457:50:@534.8]
  wire [3:0] _GEN_1168; // @[Bus.scala 456:41:@533.6]
  wire [31:0] _GEN_1169; // @[Bus.scala 456:41:@533.6]
  wire [31:0] _GEN_1170; // @[Bus.scala 456:41:@533.6]
  wire [31:0] _GEN_1171; // @[Bus.scala 456:41:@533.6]
  wire [31:0] _GEN_1172; // @[Bus.scala 456:41:@533.6]
  wire [31:0] _GEN_1173; // @[Bus.scala 456:41:@533.6]
  wire  _GEN_1174; // @[Bus.scala 456:41:@533.6]
  wire  _GEN_1175; // @[Bus.scala 456:41:@533.6]
  wire  _GEN_1176; // @[Bus.scala 456:41:@533.6]
  wire  _GEN_1177; // @[Bus.scala 456:41:@533.6]
  wire  _GEN_1178; // @[Bus.scala 456:41:@533.6]
  wire  _GEN_1179; // @[Bus.scala 456:41:@533.6]
  wire  _GEN_1180; // @[Bus.scala 456:41:@533.6]
  wire  _GEN_1181; // @[Bus.scala 456:41:@533.6]
  wire  _GEN_1182; // @[Bus.scala 456:41:@533.6]
  wire  _GEN_1183; // @[Bus.scala 456:41:@533.6]
  wire  _T_440; // @[Bus.scala 476:30:@553.6]
  wire [3:0] _GEN_1184; // @[Bus.scala 477:50:@555.8]
  wire [31:0] _GEN_1185; // @[Bus.scala 477:50:@555.8]
  wire [31:0] _GEN_1186; // @[Bus.scala 477:50:@555.8]
  wire [31:0] _GEN_1187; // @[Bus.scala 477:50:@555.8]
  wire [31:0] _GEN_1188; // @[Bus.scala 477:50:@555.8]
  wire [31:0] _GEN_1189; // @[Bus.scala 477:50:@555.8]
  wire  _GEN_1190; // @[Bus.scala 477:50:@555.8]
  wire  _GEN_1191; // @[Bus.scala 477:50:@555.8]
  wire  _GEN_1192; // @[Bus.scala 477:50:@555.8]
  wire  _GEN_1193; // @[Bus.scala 477:50:@555.8]
  wire  _GEN_1194; // @[Bus.scala 477:50:@555.8]
  wire  _GEN_1195; // @[Bus.scala 477:50:@555.8]
  wire  _GEN_1196; // @[Bus.scala 477:50:@555.8]
  wire  _GEN_1197; // @[Bus.scala 477:50:@555.8]
  wire  _GEN_1198; // @[Bus.scala 477:50:@555.8]
  wire  _GEN_1199; // @[Bus.scala 477:50:@555.8]
  wire [3:0] _GEN_1200; // @[Bus.scala 476:41:@554.6]
  wire [31:0] _GEN_1201; // @[Bus.scala 476:41:@554.6]
  wire [31:0] _GEN_1202; // @[Bus.scala 476:41:@554.6]
  wire [31:0] _GEN_1203; // @[Bus.scala 476:41:@554.6]
  wire [31:0] _GEN_1204; // @[Bus.scala 476:41:@554.6]
  wire [31:0] _GEN_1205; // @[Bus.scala 476:41:@554.6]
  wire  _GEN_1206; // @[Bus.scala 476:41:@554.6]
  wire  _GEN_1207; // @[Bus.scala 476:41:@554.6]
  wire  _GEN_1208; // @[Bus.scala 476:41:@554.6]
  wire  _GEN_1209; // @[Bus.scala 476:41:@554.6]
  wire  _GEN_1210; // @[Bus.scala 476:41:@554.6]
  wire  _GEN_1211; // @[Bus.scala 476:41:@554.6]
  wire  _GEN_1212; // @[Bus.scala 476:41:@554.6]
  wire  _GEN_1213; // @[Bus.scala 476:41:@554.6]
  wire  _GEN_1214; // @[Bus.scala 476:41:@554.6]
  wire  _GEN_1215; // @[Bus.scala 476:41:@554.6]
  wire  _T_451; // @[Bus.scala 496:30:@574.6]
  wire [3:0] _GEN_1216; // @[Bus.scala 498:57:@579.10]
  wire [31:0] _GEN_1217; // @[Bus.scala 498:57:@579.10]
  wire [31:0] _GEN_1218; // @[Bus.scala 498:57:@579.10]
  wire [31:0] _GEN_1219; // @[Bus.scala 498:57:@579.10]
  wire [31:0] _GEN_1220; // @[Bus.scala 498:57:@579.10]
  wire [31:0] _GEN_1221; // @[Bus.scala 498:57:@579.10]
  wire [31:0] _GEN_1222; // @[Bus.scala 498:57:@579.10]
  wire [31:0] _GEN_1223; // @[Bus.scala 498:57:@579.10]
  wire  _GEN_1224; // @[Bus.scala 498:57:@579.10]
  wire  _GEN_1225; // @[Bus.scala 498:57:@579.10]
  wire  _GEN_1226; // @[Bus.scala 498:57:@579.10]
  wire  _GEN_1227; // @[Bus.scala 498:57:@579.10]
  wire  _GEN_1228; // @[Bus.scala 498:57:@579.10]
  wire  _GEN_1229; // @[Bus.scala 498:57:@579.10]
  wire  _GEN_1230; // @[Bus.scala 498:57:@579.10]
  wire  _GEN_1231; // @[Bus.scala 498:57:@579.10]
  wire  _GEN_1232; // @[Bus.scala 498:57:@579.10]
  wire  _GEN_1233; // @[Bus.scala 498:57:@579.10]
  wire [3:0] _GEN_1234; // @[Bus.scala 497:75:@578.8]
  wire [31:0] _GEN_1235; // @[Bus.scala 497:75:@578.8]
  wire [31:0] _GEN_1236; // @[Bus.scala 497:75:@578.8]
  wire [31:0] _GEN_1237; // @[Bus.scala 497:75:@578.8]
  wire [31:0] _GEN_1238; // @[Bus.scala 497:75:@578.8]
  wire [31:0] _GEN_1239; // @[Bus.scala 497:75:@578.8]
  wire [31:0] _GEN_1240; // @[Bus.scala 497:75:@578.8]
  wire [31:0] _GEN_1241; // @[Bus.scala 497:75:@578.8]
  wire  _GEN_1242; // @[Bus.scala 497:75:@578.8]
  wire  _GEN_1243; // @[Bus.scala 497:75:@578.8]
  wire  _GEN_1244; // @[Bus.scala 497:75:@578.8]
  wire  _GEN_1245; // @[Bus.scala 497:75:@578.8]
  wire  _GEN_1246; // @[Bus.scala 497:75:@578.8]
  wire  _GEN_1247; // @[Bus.scala 497:75:@578.8]
  wire  _GEN_1248; // @[Bus.scala 497:75:@578.8]
  wire  _GEN_1249; // @[Bus.scala 497:75:@578.8]
  wire  _GEN_1250; // @[Bus.scala 497:75:@578.8]
  wire  _GEN_1251; // @[Bus.scala 497:75:@578.8]
  wire [3:0] _GEN_1252; // @[Bus.scala 496:41:@575.6]
  wire [31:0] _GEN_1253; // @[Bus.scala 496:41:@575.6]
  wire [31:0] _GEN_1254; // @[Bus.scala 496:41:@575.6]
  wire [31:0] _GEN_1255; // @[Bus.scala 496:41:@575.6]
  wire [31:0] _GEN_1256; // @[Bus.scala 496:41:@575.6]
  wire [31:0] _GEN_1257; // @[Bus.scala 496:41:@575.6]
  wire [31:0] _GEN_1258; // @[Bus.scala 496:41:@575.6]
  wire [31:0] _GEN_1259; // @[Bus.scala 496:41:@575.6]
  wire  _GEN_1260; // @[Bus.scala 496:41:@575.6]
  wire  _GEN_1261; // @[Bus.scala 496:41:@575.6]
  wire  _GEN_1262; // @[Bus.scala 496:41:@575.6]
  wire  _GEN_1263; // @[Bus.scala 496:41:@575.6]
  wire  _GEN_1264; // @[Bus.scala 496:41:@575.6]
  wire  _GEN_1265; // @[Bus.scala 496:41:@575.6]
  wire  _GEN_1266; // @[Bus.scala 496:41:@575.6]
  wire  _GEN_1267; // @[Bus.scala 496:41:@575.6]
  wire  _GEN_1268; // @[Bus.scala 496:41:@575.6]
  wire  _GEN_1269; // @[Bus.scala 496:41:@575.6]
  wire [3:0] _GEN_1270; // @[Bus.scala 522:57:@605.10]
  wire [31:0] _GEN_1271; // @[Bus.scala 522:57:@605.10]
  wire [31:0] _GEN_1272; // @[Bus.scala 522:57:@605.10]
  wire [31:0] _GEN_1273; // @[Bus.scala 522:57:@605.10]
  wire [31:0] _GEN_1274; // @[Bus.scala 522:57:@605.10]
  wire [31:0] _GEN_1275; // @[Bus.scala 522:57:@605.10]
  wire [31:0] _GEN_1276; // @[Bus.scala 522:57:@605.10]
  wire [31:0] _GEN_1277; // @[Bus.scala 522:57:@605.10]
  wire  _GEN_1278; // @[Bus.scala 522:57:@605.10]
  wire  _GEN_1279; // @[Bus.scala 522:57:@605.10]
  wire  _GEN_1280; // @[Bus.scala 522:57:@605.10]
  wire  _GEN_1281; // @[Bus.scala 522:57:@605.10]
  wire  _GEN_1282; // @[Bus.scala 522:57:@605.10]
  wire  _GEN_1283; // @[Bus.scala 522:57:@605.10]
  wire  _GEN_1284; // @[Bus.scala 522:57:@605.10]
  wire  _GEN_1285; // @[Bus.scala 522:57:@605.10]
  wire  _GEN_1286; // @[Bus.scala 522:57:@605.10]
  wire  _GEN_1287; // @[Bus.scala 522:57:@605.10]
  wire [3:0] _GEN_1288; // @[Bus.scala 521:74:@604.8]
  wire [31:0] _GEN_1289; // @[Bus.scala 521:74:@604.8]
  wire [31:0] _GEN_1290; // @[Bus.scala 521:74:@604.8]
  wire [31:0] _GEN_1291; // @[Bus.scala 521:74:@604.8]
  wire [31:0] _GEN_1292; // @[Bus.scala 521:74:@604.8]
  wire [31:0] _GEN_1293; // @[Bus.scala 521:74:@604.8]
  wire [31:0] _GEN_1294; // @[Bus.scala 521:74:@604.8]
  wire [31:0] _GEN_1295; // @[Bus.scala 521:74:@604.8]
  wire  _GEN_1296; // @[Bus.scala 521:74:@604.8]
  wire  _GEN_1297; // @[Bus.scala 521:74:@604.8]
  wire  _GEN_1298; // @[Bus.scala 521:74:@604.8]
  wire  _GEN_1299; // @[Bus.scala 521:74:@604.8]
  wire  _GEN_1300; // @[Bus.scala 521:74:@604.8]
  wire  _GEN_1301; // @[Bus.scala 521:74:@604.8]
  wire  _GEN_1302; // @[Bus.scala 521:74:@604.8]
  wire  _GEN_1303; // @[Bus.scala 521:74:@604.8]
  wire  _GEN_1304; // @[Bus.scala 521:74:@604.8]
  wire  _GEN_1305; // @[Bus.scala 521:74:@604.8]
  wire [3:0] _GEN_1306; // @[Bus.scala 520:41:@602.6]
  wire [31:0] _GEN_1307; // @[Bus.scala 520:41:@602.6]
  wire [31:0] _GEN_1308; // @[Bus.scala 520:41:@602.6]
  wire [31:0] _GEN_1309; // @[Bus.scala 520:41:@602.6]
  wire [31:0] _GEN_1310; // @[Bus.scala 520:41:@602.6]
  wire [31:0] _GEN_1311; // @[Bus.scala 520:41:@602.6]
  wire [31:0] _GEN_1312; // @[Bus.scala 520:41:@602.6]
  wire [31:0] _GEN_1313; // @[Bus.scala 520:41:@602.6]
  wire  _GEN_1314; // @[Bus.scala 520:41:@602.6]
  wire  _GEN_1315; // @[Bus.scala 520:41:@602.6]
  wire  _GEN_1316; // @[Bus.scala 520:41:@602.6]
  wire  _GEN_1317; // @[Bus.scala 520:41:@602.6]
  wire  _GEN_1318; // @[Bus.scala 520:41:@602.6]
  wire  _GEN_1319; // @[Bus.scala 520:41:@602.6]
  wire  _GEN_1320; // @[Bus.scala 520:41:@602.6]
  wire  _GEN_1321; // @[Bus.scala 520:41:@602.6]
  wire  _GEN_1322; // @[Bus.scala 520:41:@602.6]
  wire  _GEN_1323; // @[Bus.scala 520:41:@602.6]
  wire  _T_479; // @[Bus.scala 544:30:@627.6]
  wire [3:0] _GEN_1324; // @[Bus.scala 545:50:@629.8]
  wire [31:0] _GEN_1325; // @[Bus.scala 545:50:@629.8]
  wire [31:0] _GEN_1326; // @[Bus.scala 545:50:@629.8]
  wire [31:0] _GEN_1327; // @[Bus.scala 545:50:@629.8]
  wire [31:0] _GEN_1328; // @[Bus.scala 545:50:@629.8]
  wire [31:0] _GEN_1329; // @[Bus.scala 545:50:@629.8]
  wire  _GEN_1330; // @[Bus.scala 545:50:@629.8]
  wire  _GEN_1331; // @[Bus.scala 545:50:@629.8]
  wire  _GEN_1332; // @[Bus.scala 545:50:@629.8]
  wire  _GEN_1333; // @[Bus.scala 545:50:@629.8]
  wire  _GEN_1334; // @[Bus.scala 545:50:@629.8]
  wire  _GEN_1335; // @[Bus.scala 545:50:@629.8]
  wire  _GEN_1336; // @[Bus.scala 545:50:@629.8]
  wire  _GEN_1337; // @[Bus.scala 545:50:@629.8]
  wire  _GEN_1338; // @[Bus.scala 545:50:@629.8]
  wire  _GEN_1339; // @[Bus.scala 545:50:@629.8]
  wire [3:0] _GEN_1340; // @[Bus.scala 544:41:@628.6]
  wire [31:0] _GEN_1341; // @[Bus.scala 544:41:@628.6]
  wire [31:0] _GEN_1342; // @[Bus.scala 544:41:@628.6]
  wire [31:0] _GEN_1343; // @[Bus.scala 544:41:@628.6]
  wire [31:0] _GEN_1344; // @[Bus.scala 544:41:@628.6]
  wire [31:0] _GEN_1345; // @[Bus.scala 544:41:@628.6]
  wire  _GEN_1346; // @[Bus.scala 544:41:@628.6]
  wire  _GEN_1347; // @[Bus.scala 544:41:@628.6]
  wire  _GEN_1348; // @[Bus.scala 544:41:@628.6]
  wire  _GEN_1349; // @[Bus.scala 544:41:@628.6]
  wire  _GEN_1350; // @[Bus.scala 544:41:@628.6]
  wire  _GEN_1351; // @[Bus.scala 544:41:@628.6]
  wire  _GEN_1352; // @[Bus.scala 544:41:@628.6]
  wire  _GEN_1353; // @[Bus.scala 544:41:@628.6]
  wire  _GEN_1354; // @[Bus.scala 544:41:@628.6]
  wire  _GEN_1355; // @[Bus.scala 544:41:@628.6]
  wire  _T_490; // @[Bus.scala 564:30:@648.6]
  wire [3:0] _GEN_1356; // @[Bus.scala 566:57:@653.10]
  wire [31:0] _GEN_1357; // @[Bus.scala 566:57:@653.10]
  wire [31:0] _GEN_1358; // @[Bus.scala 566:57:@653.10]
  wire [31:0] _GEN_1359; // @[Bus.scala 566:57:@653.10]
  wire [31:0] _GEN_1360; // @[Bus.scala 566:57:@653.10]
  wire [31:0] _GEN_1361; // @[Bus.scala 566:57:@653.10]
  wire [31:0] _GEN_1362; // @[Bus.scala 566:57:@653.10]
  wire [31:0] _GEN_1363; // @[Bus.scala 566:57:@653.10]
  wire  _GEN_1364; // @[Bus.scala 566:57:@653.10]
  wire  _GEN_1365; // @[Bus.scala 566:57:@653.10]
  wire  _GEN_1366; // @[Bus.scala 566:57:@653.10]
  wire  _GEN_1367; // @[Bus.scala 566:57:@653.10]
  wire  _GEN_1368; // @[Bus.scala 566:57:@653.10]
  wire  _GEN_1369; // @[Bus.scala 566:57:@653.10]
  wire  _GEN_1370; // @[Bus.scala 566:57:@653.10]
  wire  _GEN_1371; // @[Bus.scala 566:57:@653.10]
  wire  _GEN_1372; // @[Bus.scala 566:57:@653.10]
  wire  _GEN_1373; // @[Bus.scala 566:57:@653.10]
  wire [3:0] _GEN_1374; // @[Bus.scala 565:75:@652.8]
  wire [31:0] _GEN_1375; // @[Bus.scala 565:75:@652.8]
  wire [31:0] _GEN_1376; // @[Bus.scala 565:75:@652.8]
  wire [31:0] _GEN_1377; // @[Bus.scala 565:75:@652.8]
  wire [31:0] _GEN_1378; // @[Bus.scala 565:75:@652.8]
  wire [31:0] _GEN_1379; // @[Bus.scala 565:75:@652.8]
  wire [31:0] _GEN_1380; // @[Bus.scala 565:75:@652.8]
  wire [31:0] _GEN_1381; // @[Bus.scala 565:75:@652.8]
  wire  _GEN_1382; // @[Bus.scala 565:75:@652.8]
  wire  _GEN_1383; // @[Bus.scala 565:75:@652.8]
  wire  _GEN_1384; // @[Bus.scala 565:75:@652.8]
  wire  _GEN_1385; // @[Bus.scala 565:75:@652.8]
  wire  _GEN_1386; // @[Bus.scala 565:75:@652.8]
  wire  _GEN_1387; // @[Bus.scala 565:75:@652.8]
  wire  _GEN_1388; // @[Bus.scala 565:75:@652.8]
  wire  _GEN_1389; // @[Bus.scala 565:75:@652.8]
  wire  _GEN_1390; // @[Bus.scala 565:75:@652.8]
  wire  _GEN_1391; // @[Bus.scala 565:75:@652.8]
  wire [3:0] _GEN_1392; // @[Bus.scala 564:41:@649.6]
  wire [31:0] _GEN_1393; // @[Bus.scala 564:41:@649.6]
  wire [31:0] _GEN_1394; // @[Bus.scala 564:41:@649.6]
  wire [31:0] _GEN_1395; // @[Bus.scala 564:41:@649.6]
  wire [31:0] _GEN_1396; // @[Bus.scala 564:41:@649.6]
  wire [31:0] _GEN_1397; // @[Bus.scala 564:41:@649.6]
  wire [31:0] _GEN_1398; // @[Bus.scala 564:41:@649.6]
  wire [31:0] _GEN_1399; // @[Bus.scala 564:41:@649.6]
  wire  _GEN_1400; // @[Bus.scala 564:41:@649.6]
  wire  _GEN_1401; // @[Bus.scala 564:41:@649.6]
  wire  _GEN_1402; // @[Bus.scala 564:41:@649.6]
  wire  _GEN_1403; // @[Bus.scala 564:41:@649.6]
  wire  _GEN_1404; // @[Bus.scala 564:41:@649.6]
  wire  _GEN_1405; // @[Bus.scala 564:41:@649.6]
  wire  _GEN_1406; // @[Bus.scala 564:41:@649.6]
  wire  _GEN_1407; // @[Bus.scala 564:41:@649.6]
  wire  _GEN_1408; // @[Bus.scala 564:41:@649.6]
  wire  _GEN_1409; // @[Bus.scala 564:41:@649.6]
  wire [3:0] _GEN_1410; // @[Bus.scala 590:57:@679.10]
  wire [31:0] _GEN_1411; // @[Bus.scala 590:57:@679.10]
  wire [31:0] _GEN_1412; // @[Bus.scala 590:57:@679.10]
  wire [31:0] _GEN_1413; // @[Bus.scala 590:57:@679.10]
  wire [31:0] _GEN_1414; // @[Bus.scala 590:57:@679.10]
  wire [31:0] _GEN_1415; // @[Bus.scala 590:57:@679.10]
  wire [31:0] _GEN_1416; // @[Bus.scala 590:57:@679.10]
  wire [31:0] _GEN_1417; // @[Bus.scala 590:57:@679.10]
  wire  _GEN_1418; // @[Bus.scala 590:57:@679.10]
  wire  _GEN_1419; // @[Bus.scala 590:57:@679.10]
  wire  _GEN_1420; // @[Bus.scala 590:57:@679.10]
  wire  _GEN_1421; // @[Bus.scala 590:57:@679.10]
  wire  _GEN_1422; // @[Bus.scala 590:57:@679.10]
  wire  _GEN_1423; // @[Bus.scala 590:57:@679.10]
  wire  _GEN_1424; // @[Bus.scala 590:57:@679.10]
  wire  _GEN_1425; // @[Bus.scala 590:57:@679.10]
  wire  _GEN_1426; // @[Bus.scala 590:57:@679.10]
  wire  _GEN_1427; // @[Bus.scala 590:57:@679.10]
  wire [3:0] _GEN_1428; // @[Bus.scala 589:74:@678.8]
  wire [31:0] _GEN_1429; // @[Bus.scala 589:74:@678.8]
  wire [31:0] _GEN_1430; // @[Bus.scala 589:74:@678.8]
  wire [31:0] _GEN_1431; // @[Bus.scala 589:74:@678.8]
  wire [31:0] _GEN_1432; // @[Bus.scala 589:74:@678.8]
  wire [31:0] _GEN_1433; // @[Bus.scala 589:74:@678.8]
  wire [31:0] _GEN_1434; // @[Bus.scala 589:74:@678.8]
  wire [31:0] _GEN_1435; // @[Bus.scala 589:74:@678.8]
  wire  _GEN_1436; // @[Bus.scala 589:74:@678.8]
  wire  _GEN_1437; // @[Bus.scala 589:74:@678.8]
  wire  _GEN_1438; // @[Bus.scala 589:74:@678.8]
  wire  _GEN_1439; // @[Bus.scala 589:74:@678.8]
  wire  _GEN_1440; // @[Bus.scala 589:74:@678.8]
  wire  _GEN_1441; // @[Bus.scala 589:74:@678.8]
  wire  _GEN_1442; // @[Bus.scala 589:74:@678.8]
  wire  _GEN_1443; // @[Bus.scala 589:74:@678.8]
  wire  _GEN_1444; // @[Bus.scala 589:74:@678.8]
  wire  _GEN_1445; // @[Bus.scala 589:74:@678.8]
  wire [3:0] _GEN_1446; // @[Bus.scala 588:41:@676.6]
  wire [31:0] _GEN_1447; // @[Bus.scala 588:41:@676.6]
  wire [31:0] _GEN_1448; // @[Bus.scala 588:41:@676.6]
  wire [31:0] _GEN_1449; // @[Bus.scala 588:41:@676.6]
  wire [31:0] _GEN_1450; // @[Bus.scala 588:41:@676.6]
  wire [31:0] _GEN_1451; // @[Bus.scala 588:41:@676.6]
  wire [31:0] _GEN_1452; // @[Bus.scala 588:41:@676.6]
  wire [31:0] _GEN_1453; // @[Bus.scala 588:41:@676.6]
  wire  _GEN_1454; // @[Bus.scala 588:41:@676.6]
  wire  _GEN_1455; // @[Bus.scala 588:41:@676.6]
  wire  _GEN_1456; // @[Bus.scala 588:41:@676.6]
  wire  _GEN_1457; // @[Bus.scala 588:41:@676.6]
  wire  _GEN_1458; // @[Bus.scala 588:41:@676.6]
  wire  _GEN_1459; // @[Bus.scala 588:41:@676.6]
  wire  _GEN_1460; // @[Bus.scala 588:41:@676.6]
  wire  _GEN_1461; // @[Bus.scala 588:41:@676.6]
  wire  _GEN_1462; // @[Bus.scala 588:41:@676.6]
  wire  _GEN_1463; // @[Bus.scala 588:41:@676.6]
  wire  _T_518; // @[Bus.scala 612:30:@701.6]
  wire [3:0] _GEN_1464; // @[Bus.scala 613:50:@703.8]
  wire [31:0] _GEN_1465; // @[Bus.scala 613:50:@703.8]
  wire [31:0] _GEN_1466; // @[Bus.scala 613:50:@703.8]
  wire [31:0] _GEN_1467; // @[Bus.scala 613:50:@703.8]
  wire [31:0] _GEN_1468; // @[Bus.scala 613:50:@703.8]
  wire [31:0] _GEN_1469; // @[Bus.scala 613:50:@703.8]
  wire  _GEN_1470; // @[Bus.scala 613:50:@703.8]
  wire  _GEN_1471; // @[Bus.scala 613:50:@703.8]
  wire  _GEN_1472; // @[Bus.scala 613:50:@703.8]
  wire  _GEN_1473; // @[Bus.scala 613:50:@703.8]
  wire  _GEN_1474; // @[Bus.scala 613:50:@703.8]
  wire  _GEN_1475; // @[Bus.scala 613:50:@703.8]
  wire  _GEN_1476; // @[Bus.scala 613:50:@703.8]
  wire  _GEN_1477; // @[Bus.scala 613:50:@703.8]
  wire  _GEN_1478; // @[Bus.scala 613:50:@703.8]
  wire  _GEN_1479; // @[Bus.scala 613:50:@703.8]
  wire [3:0] _GEN_1480; // @[Bus.scala 612:41:@702.6]
  wire [31:0] _GEN_1481; // @[Bus.scala 612:41:@702.6]
  wire [31:0] _GEN_1482; // @[Bus.scala 612:41:@702.6]
  wire [31:0] _GEN_1483; // @[Bus.scala 612:41:@702.6]
  wire [31:0] _GEN_1484; // @[Bus.scala 612:41:@702.6]
  wire [31:0] _GEN_1485; // @[Bus.scala 612:41:@702.6]
  wire  _GEN_1486; // @[Bus.scala 612:41:@702.6]
  wire  _GEN_1487; // @[Bus.scala 612:41:@702.6]
  wire  _GEN_1488; // @[Bus.scala 612:41:@702.6]
  wire  _GEN_1489; // @[Bus.scala 612:41:@702.6]
  wire  _GEN_1490; // @[Bus.scala 612:41:@702.6]
  wire  _GEN_1491; // @[Bus.scala 612:41:@702.6]
  wire  _GEN_1492; // @[Bus.scala 612:41:@702.6]
  wire  _GEN_1493; // @[Bus.scala 612:41:@702.6]
  wire  _GEN_1494; // @[Bus.scala 612:41:@702.6]
  wire  _GEN_1495; // @[Bus.scala 612:41:@702.6]
  wire  _T_529; // @[Bus.scala 632:30:@722.6]
  wire [3:0] _GEN_1496; // @[Bus.scala 634:57:@727.10]
  wire [31:0] _GEN_1497; // @[Bus.scala 634:57:@727.10]
  wire [31:0] _GEN_1498; // @[Bus.scala 634:57:@727.10]
  wire [31:0] _GEN_1499; // @[Bus.scala 634:57:@727.10]
  wire [31:0] _GEN_1500; // @[Bus.scala 634:57:@727.10]
  wire [31:0] _GEN_1501; // @[Bus.scala 634:57:@727.10]
  wire [31:0] _GEN_1502; // @[Bus.scala 634:57:@727.10]
  wire [31:0] _GEN_1503; // @[Bus.scala 634:57:@727.10]
  wire  _GEN_1504; // @[Bus.scala 634:57:@727.10]
  wire  _GEN_1505; // @[Bus.scala 634:57:@727.10]
  wire  _GEN_1506; // @[Bus.scala 634:57:@727.10]
  wire  _GEN_1507; // @[Bus.scala 634:57:@727.10]
  wire  _GEN_1508; // @[Bus.scala 634:57:@727.10]
  wire  _GEN_1509; // @[Bus.scala 634:57:@727.10]
  wire  _GEN_1510; // @[Bus.scala 634:57:@727.10]
  wire  _GEN_1511; // @[Bus.scala 634:57:@727.10]
  wire  _GEN_1512; // @[Bus.scala 634:57:@727.10]
  wire  _GEN_1513; // @[Bus.scala 634:57:@727.10]
  wire [3:0] _GEN_1514; // @[Bus.scala 633:75:@726.8]
  wire [31:0] _GEN_1515; // @[Bus.scala 633:75:@726.8]
  wire [31:0] _GEN_1516; // @[Bus.scala 633:75:@726.8]
  wire [31:0] _GEN_1517; // @[Bus.scala 633:75:@726.8]
  wire [31:0] _GEN_1518; // @[Bus.scala 633:75:@726.8]
  wire [31:0] _GEN_1519; // @[Bus.scala 633:75:@726.8]
  wire [31:0] _GEN_1520; // @[Bus.scala 633:75:@726.8]
  wire [31:0] _GEN_1521; // @[Bus.scala 633:75:@726.8]
  wire  _GEN_1522; // @[Bus.scala 633:75:@726.8]
  wire  _GEN_1523; // @[Bus.scala 633:75:@726.8]
  wire  _GEN_1524; // @[Bus.scala 633:75:@726.8]
  wire  _GEN_1525; // @[Bus.scala 633:75:@726.8]
  wire  _GEN_1526; // @[Bus.scala 633:75:@726.8]
  wire  _GEN_1527; // @[Bus.scala 633:75:@726.8]
  wire  _GEN_1528; // @[Bus.scala 633:75:@726.8]
  wire  _GEN_1529; // @[Bus.scala 633:75:@726.8]
  wire  _GEN_1530; // @[Bus.scala 633:75:@726.8]
  wire  _GEN_1531; // @[Bus.scala 633:75:@726.8]
  wire [3:0] _GEN_1532; // @[Bus.scala 632:41:@723.6]
  wire [31:0] _GEN_1533; // @[Bus.scala 632:41:@723.6]
  wire [31:0] _GEN_1534; // @[Bus.scala 632:41:@723.6]
  wire [31:0] _GEN_1535; // @[Bus.scala 632:41:@723.6]
  wire [31:0] _GEN_1536; // @[Bus.scala 632:41:@723.6]
  wire [31:0] _GEN_1537; // @[Bus.scala 632:41:@723.6]
  wire [31:0] _GEN_1538; // @[Bus.scala 632:41:@723.6]
  wire [31:0] _GEN_1539; // @[Bus.scala 632:41:@723.6]
  wire  _GEN_1540; // @[Bus.scala 632:41:@723.6]
  wire  _GEN_1541; // @[Bus.scala 632:41:@723.6]
  wire  _GEN_1542; // @[Bus.scala 632:41:@723.6]
  wire  _GEN_1543; // @[Bus.scala 632:41:@723.6]
  wire  _GEN_1544; // @[Bus.scala 632:41:@723.6]
  wire  _GEN_1545; // @[Bus.scala 632:41:@723.6]
  wire  _GEN_1546; // @[Bus.scala 632:41:@723.6]
  wire  _GEN_1547; // @[Bus.scala 632:41:@723.6]
  wire  _GEN_1548; // @[Bus.scala 632:41:@723.6]
  wire  _GEN_1549; // @[Bus.scala 632:41:@723.6]
  wire [3:0] _GEN_1550; // @[Bus.scala 658:57:@753.10]
  wire [31:0] _GEN_1551; // @[Bus.scala 658:57:@753.10]
  wire [31:0] _GEN_1552; // @[Bus.scala 658:57:@753.10]
  wire [31:0] _GEN_1553; // @[Bus.scala 658:57:@753.10]
  wire [31:0] _GEN_1554; // @[Bus.scala 658:57:@753.10]
  wire [31:0] _GEN_1555; // @[Bus.scala 658:57:@753.10]
  wire [31:0] _GEN_1556; // @[Bus.scala 658:57:@753.10]
  wire [31:0] _GEN_1557; // @[Bus.scala 658:57:@753.10]
  wire  _GEN_1558; // @[Bus.scala 658:57:@753.10]
  wire  _GEN_1559; // @[Bus.scala 658:57:@753.10]
  wire  _GEN_1560; // @[Bus.scala 658:57:@753.10]
  wire  _GEN_1561; // @[Bus.scala 658:57:@753.10]
  wire  _GEN_1562; // @[Bus.scala 658:57:@753.10]
  wire  _GEN_1563; // @[Bus.scala 658:57:@753.10]
  wire  _GEN_1564; // @[Bus.scala 658:57:@753.10]
  wire  _GEN_1565; // @[Bus.scala 658:57:@753.10]
  wire  _GEN_1566; // @[Bus.scala 658:57:@753.10]
  wire  _GEN_1567; // @[Bus.scala 658:57:@753.10]
  wire [3:0] _GEN_1568; // @[Bus.scala 657:74:@752.8]
  wire [31:0] _GEN_1569; // @[Bus.scala 657:74:@752.8]
  wire [31:0] _GEN_1570; // @[Bus.scala 657:74:@752.8]
  wire [31:0] _GEN_1571; // @[Bus.scala 657:74:@752.8]
  wire [31:0] _GEN_1572; // @[Bus.scala 657:74:@752.8]
  wire [31:0] _GEN_1573; // @[Bus.scala 657:74:@752.8]
  wire [31:0] _GEN_1574; // @[Bus.scala 657:74:@752.8]
  wire [31:0] _GEN_1575; // @[Bus.scala 657:74:@752.8]
  wire  _GEN_1576; // @[Bus.scala 657:74:@752.8]
  wire  _GEN_1577; // @[Bus.scala 657:74:@752.8]
  wire  _GEN_1578; // @[Bus.scala 657:74:@752.8]
  wire  _GEN_1579; // @[Bus.scala 657:74:@752.8]
  wire  _GEN_1580; // @[Bus.scala 657:74:@752.8]
  wire  _GEN_1581; // @[Bus.scala 657:74:@752.8]
  wire  _GEN_1582; // @[Bus.scala 657:74:@752.8]
  wire  _GEN_1583; // @[Bus.scala 657:74:@752.8]
  wire  _GEN_1584; // @[Bus.scala 657:74:@752.8]
  wire  _GEN_1585; // @[Bus.scala 657:74:@752.8]
  wire [3:0] _GEN_1586; // @[Bus.scala 656:41:@750.6]
  wire [31:0] _GEN_1587; // @[Bus.scala 656:41:@750.6]
  wire [31:0] _GEN_1588; // @[Bus.scala 656:41:@750.6]
  wire [31:0] _GEN_1589; // @[Bus.scala 656:41:@750.6]
  wire [31:0] _GEN_1590; // @[Bus.scala 656:41:@750.6]
  wire [31:0] _GEN_1591; // @[Bus.scala 656:41:@750.6]
  wire [31:0] _GEN_1592; // @[Bus.scala 656:41:@750.6]
  wire [31:0] _GEN_1593; // @[Bus.scala 656:41:@750.6]
  wire  _GEN_1594; // @[Bus.scala 656:41:@750.6]
  wire  _GEN_1595; // @[Bus.scala 656:41:@750.6]
  wire  _GEN_1596; // @[Bus.scala 656:41:@750.6]
  wire  _GEN_1597; // @[Bus.scala 656:41:@750.6]
  wire  _GEN_1598; // @[Bus.scala 656:41:@750.6]
  wire  _GEN_1599; // @[Bus.scala 656:41:@750.6]
  wire  _GEN_1600; // @[Bus.scala 656:41:@750.6]
  wire  _GEN_1601; // @[Bus.scala 656:41:@750.6]
  wire  _GEN_1602; // @[Bus.scala 656:41:@750.6]
  wire  _GEN_1603; // @[Bus.scala 656:41:@750.6]
  assign _T_97 = state_r == 4'h0; // @[Bus.scala 92:30:@46.6]
  assign _T_98 = 32'h0 == io_master_in_trans_type; // @[Bus.scala 93:44:@48.8]
  assign _T_100 = _T_98 == 1'h0; // @[Bus.scala 93:30:@49.8]
  assign _T_102 = $signed(io_master_in_addr) >= $signed(32'sh0); // @[Bus.scala 94:57:@51.10]
  assign _T_104 = $signed(io_master_in_addr) <= $signed(32'sh7); // @[Bus.scala 95:65:@53.12]
  assign _GEN_0 = io_master_in_sync ? 4'h1 : state_r; // @[Bus.scala 96:73:@55.14]
  assign _GEN_1 = io_master_in_sync ? $signed(io_master_in_addr) : $signed(req_signal_r_addr); // @[Bus.scala 96:73:@55.14]
  assign _GEN_2 = io_master_in_sync ? $signed(io_master_in_data) : $signed(req_signal_r_data); // @[Bus.scala 96:73:@55.14]
  assign _GEN_3 = io_master_in_sync ? io_master_in_trans_type : req_signal_r_trans_type; // @[Bus.scala 96:73:@55.14]
  assign _GEN_6 = io_master_in_sync ? $signed(io_master_in_addr) : $signed(slave_out0_r_addr); // @[Bus.scala 96:73:@55.14]
  assign _GEN_7 = io_master_in_sync ? $signed(io_master_in_data) : $signed(slave_out0_r_data); // @[Bus.scala 96:73:@55.14]
  assign _GEN_8 = io_master_in_sync ? io_master_in_trans_type : slave_out0_r_trans_type; // @[Bus.scala 96:73:@55.14]
  assign _GEN_9 = io_master_in_sync ? 1'h0 : master_in_notify_r; // @[Bus.scala 96:73:@55.14]
  assign _GEN_10 = io_master_in_sync ? 1'h0 : master_out_notify_r; // @[Bus.scala 96:73:@55.14]
  assign _GEN_11 = io_master_in_sync ? 1'h0 : slave_in0_notify_r; // @[Bus.scala 96:73:@55.14]
  assign _GEN_12 = io_master_in_sync ? 1'h0 : slave_in1_notify_r; // @[Bus.scala 96:73:@55.14]
  assign _GEN_13 = io_master_in_sync ? 1'h0 : slave_in2_notify_r; // @[Bus.scala 96:73:@55.14]
  assign _GEN_14 = io_master_in_sync ? 1'h0 : slave_in3_notify_r; // @[Bus.scala 96:73:@55.14]
  assign _GEN_15 = io_master_in_sync ? 1'h1 : slave_out0_notify_r; // @[Bus.scala 96:73:@55.14]
  assign _GEN_16 = io_master_in_sync ? 1'h0 : slave_out1_notify_r; // @[Bus.scala 96:73:@55.14]
  assign _GEN_17 = io_master_in_sync ? 1'h0 : slave_out2_notify_r; // @[Bus.scala 96:73:@55.14]
  assign _GEN_18 = io_master_in_sync ? 1'h0 : slave_out3_notify_r; // @[Bus.scala 96:73:@55.14]
  assign _GEN_19 = _T_104 ? _GEN_0 : state_r; // @[Bus.scala 95:80:@54.12]
  assign _GEN_20 = _T_104 ? $signed(_GEN_1) : $signed(req_signal_r_addr); // @[Bus.scala 95:80:@54.12]
  assign _GEN_21 = _T_104 ? $signed(_GEN_2) : $signed(req_signal_r_data); // @[Bus.scala 95:80:@54.12]
  assign _GEN_22 = _T_104 ? _GEN_3 : req_signal_r_trans_type; // @[Bus.scala 95:80:@54.12]
  assign _GEN_25 = _T_104 ? $signed(_GEN_6) : $signed(slave_out0_r_addr); // @[Bus.scala 95:80:@54.12]
  assign _GEN_26 = _T_104 ? $signed(_GEN_7) : $signed(slave_out0_r_data); // @[Bus.scala 95:80:@54.12]
  assign _GEN_27 = _T_104 ? _GEN_8 : slave_out0_r_trans_type; // @[Bus.scala 95:80:@54.12]
  assign _GEN_28 = _T_104 ? _GEN_9 : master_in_notify_r; // @[Bus.scala 95:80:@54.12]
  assign _GEN_29 = _T_104 ? _GEN_10 : master_out_notify_r; // @[Bus.scala 95:80:@54.12]
  assign _GEN_30 = _T_104 ? _GEN_11 : slave_in0_notify_r; // @[Bus.scala 95:80:@54.12]
  assign _GEN_31 = _T_104 ? _GEN_12 : slave_in1_notify_r; // @[Bus.scala 95:80:@54.12]
  assign _GEN_32 = _T_104 ? _GEN_13 : slave_in2_notify_r; // @[Bus.scala 95:80:@54.12]
  assign _GEN_33 = _T_104 ? _GEN_14 : slave_in3_notify_r; // @[Bus.scala 95:80:@54.12]
  assign _GEN_34 = _T_104 ? _GEN_15 : slave_out0_notify_r; // @[Bus.scala 95:80:@54.12]
  assign _GEN_35 = _T_104 ? _GEN_16 : slave_out1_notify_r; // @[Bus.scala 95:80:@54.12]
  assign _GEN_36 = _T_104 ? _GEN_17 : slave_out2_notify_r; // @[Bus.scala 95:80:@54.12]
  assign _GEN_37 = _T_104 ? _GEN_18 : slave_out3_notify_r; // @[Bus.scala 95:80:@54.12]
  assign _GEN_38 = _T_102 ? _GEN_19 : state_r; // @[Bus.scala 94:72:@52.10]
  assign _GEN_39 = _T_102 ? $signed(_GEN_20) : $signed(req_signal_r_addr); // @[Bus.scala 94:72:@52.10]
  assign _GEN_40 = _T_102 ? $signed(_GEN_21) : $signed(req_signal_r_data); // @[Bus.scala 94:72:@52.10]
  assign _GEN_41 = _T_102 ? _GEN_22 : req_signal_r_trans_type; // @[Bus.scala 94:72:@52.10]
  assign _GEN_44 = _T_102 ? $signed(_GEN_25) : $signed(slave_out0_r_addr); // @[Bus.scala 94:72:@52.10]
  assign _GEN_45 = _T_102 ? $signed(_GEN_26) : $signed(slave_out0_r_data); // @[Bus.scala 94:72:@52.10]
  assign _GEN_46 = _T_102 ? _GEN_27 : slave_out0_r_trans_type; // @[Bus.scala 94:72:@52.10]
  assign _GEN_47 = _T_102 ? _GEN_28 : master_in_notify_r; // @[Bus.scala 94:72:@52.10]
  assign _GEN_48 = _T_102 ? _GEN_29 : master_out_notify_r; // @[Bus.scala 94:72:@52.10]
  assign _GEN_49 = _T_102 ? _GEN_30 : slave_in0_notify_r; // @[Bus.scala 94:72:@52.10]
  assign _GEN_50 = _T_102 ? _GEN_31 : slave_in1_notify_r; // @[Bus.scala 94:72:@52.10]
  assign _GEN_51 = _T_102 ? _GEN_32 : slave_in2_notify_r; // @[Bus.scala 94:72:@52.10]
  assign _GEN_52 = _T_102 ? _GEN_33 : slave_in3_notify_r; // @[Bus.scala 94:72:@52.10]
  assign _GEN_53 = _T_102 ? _GEN_34 : slave_out0_notify_r; // @[Bus.scala 94:72:@52.10]
  assign _GEN_54 = _T_102 ? _GEN_35 : slave_out1_notify_r; // @[Bus.scala 94:72:@52.10]
  assign _GEN_55 = _T_102 ? _GEN_36 : slave_out2_notify_r; // @[Bus.scala 94:72:@52.10]
  assign _GEN_56 = _T_102 ? _GEN_37 : slave_out3_notify_r; // @[Bus.scala 94:72:@52.10]
  assign _GEN_57 = _T_100 ? _GEN_38 : state_r; // @[Bus.scala 93:74:@50.8]
  assign _GEN_58 = _T_100 ? $signed(_GEN_39) : $signed(req_signal_r_addr); // @[Bus.scala 93:74:@50.8]
  assign _GEN_59 = _T_100 ? $signed(_GEN_40) : $signed(req_signal_r_data); // @[Bus.scala 93:74:@50.8]
  assign _GEN_60 = _T_100 ? _GEN_41 : req_signal_r_trans_type; // @[Bus.scala 93:74:@50.8]
  assign _GEN_63 = _T_100 ? $signed(_GEN_44) : $signed(slave_out0_r_addr); // @[Bus.scala 93:74:@50.8]
  assign _GEN_64 = _T_100 ? $signed(_GEN_45) : $signed(slave_out0_r_data); // @[Bus.scala 93:74:@50.8]
  assign _GEN_65 = _T_100 ? _GEN_46 : slave_out0_r_trans_type; // @[Bus.scala 93:74:@50.8]
  assign _GEN_66 = _T_100 ? _GEN_47 : master_in_notify_r; // @[Bus.scala 93:74:@50.8]
  assign _GEN_67 = _T_100 ? _GEN_48 : master_out_notify_r; // @[Bus.scala 93:74:@50.8]
  assign _GEN_68 = _T_100 ? _GEN_49 : slave_in0_notify_r; // @[Bus.scala 93:74:@50.8]
  assign _GEN_69 = _T_100 ? _GEN_50 : slave_in1_notify_r; // @[Bus.scala 93:74:@50.8]
  assign _GEN_70 = _T_100 ? _GEN_51 : slave_in2_notify_r; // @[Bus.scala 93:74:@50.8]
  assign _GEN_71 = _T_100 ? _GEN_52 : slave_in3_notify_r; // @[Bus.scala 93:74:@50.8]
  assign _GEN_72 = _T_100 ? _GEN_53 : slave_out0_notify_r; // @[Bus.scala 93:74:@50.8]
  assign _GEN_73 = _T_100 ? _GEN_54 : slave_out1_notify_r; // @[Bus.scala 93:74:@50.8]
  assign _GEN_74 = _T_100 ? _GEN_55 : slave_out2_notify_r; // @[Bus.scala 93:74:@50.8]
  assign _GEN_75 = _T_100 ? _GEN_56 : slave_out3_notify_r; // @[Bus.scala 93:74:@50.8]
  assign _GEN_76 = _T_97 ? _GEN_57 : state_r; // @[Bus.scala 92:41:@47.6]
  assign _GEN_77 = _T_97 ? $signed(_GEN_58) : $signed(req_signal_r_addr); // @[Bus.scala 92:41:@47.6]
  assign _GEN_78 = _T_97 ? $signed(_GEN_59) : $signed(req_signal_r_data); // @[Bus.scala 92:41:@47.6]
  assign _GEN_79 = _T_97 ? _GEN_60 : req_signal_r_trans_type; // @[Bus.scala 92:41:@47.6]
  assign _GEN_82 = _T_97 ? $signed(_GEN_63) : $signed(slave_out0_r_addr); // @[Bus.scala 92:41:@47.6]
  assign _GEN_83 = _T_97 ? $signed(_GEN_64) : $signed(slave_out0_r_data); // @[Bus.scala 92:41:@47.6]
  assign _GEN_84 = _T_97 ? _GEN_65 : slave_out0_r_trans_type; // @[Bus.scala 92:41:@47.6]
  assign _GEN_85 = _T_97 ? _GEN_66 : master_in_notify_r; // @[Bus.scala 92:41:@47.6]
  assign _GEN_86 = _T_97 ? _GEN_67 : master_out_notify_r; // @[Bus.scala 92:41:@47.6]
  assign _GEN_87 = _T_97 ? _GEN_68 : slave_in0_notify_r; // @[Bus.scala 92:41:@47.6]
  assign _GEN_88 = _T_97 ? _GEN_69 : slave_in1_notify_r; // @[Bus.scala 92:41:@47.6]
  assign _GEN_89 = _T_97 ? _GEN_70 : slave_in2_notify_r; // @[Bus.scala 92:41:@47.6]
  assign _GEN_90 = _T_97 ? _GEN_71 : slave_in3_notify_r; // @[Bus.scala 92:41:@47.6]
  assign _GEN_91 = _T_97 ? _GEN_72 : slave_out0_notify_r; // @[Bus.scala 92:41:@47.6]
  assign _GEN_92 = _T_97 ? _GEN_73 : slave_out1_notify_r; // @[Bus.scala 92:41:@47.6]
  assign _GEN_93 = _T_97 ? _GEN_74 : slave_out2_notify_r; // @[Bus.scala 92:41:@47.6]
  assign _GEN_94 = _T_97 ? _GEN_75 : slave_out3_notify_r; // @[Bus.scala 92:41:@47.6]
  assign _GEN_95 = io_master_in_sync ? 4'h1 : _GEN_76; // @[Bus.scala 125:73:@88.14]
  assign _GEN_96 = io_master_in_sync ? $signed(io_master_in_addr) : $signed(_GEN_77); // @[Bus.scala 125:73:@88.14]
  assign _GEN_97 = io_master_in_sync ? $signed(32'sh0) : $signed(_GEN_78); // @[Bus.scala 125:73:@88.14]
  assign _GEN_98 = io_master_in_sync ? io_master_in_trans_type : _GEN_79; // @[Bus.scala 125:73:@88.14]
  assign _GEN_101 = io_master_in_sync ? $signed(io_master_in_addr) : $signed(_GEN_82); // @[Bus.scala 125:73:@88.14]
  assign _GEN_102 = io_master_in_sync ? $signed(32'sh0) : $signed(_GEN_83); // @[Bus.scala 125:73:@88.14]
  assign _GEN_103 = io_master_in_sync ? io_master_in_trans_type : _GEN_84; // @[Bus.scala 125:73:@88.14]
  assign _GEN_104 = io_master_in_sync ? 1'h0 : _GEN_85; // @[Bus.scala 125:73:@88.14]
  assign _GEN_105 = io_master_in_sync ? 1'h0 : _GEN_86; // @[Bus.scala 125:73:@88.14]
  assign _GEN_106 = io_master_in_sync ? 1'h0 : _GEN_87; // @[Bus.scala 125:73:@88.14]
  assign _GEN_107 = io_master_in_sync ? 1'h0 : _GEN_88; // @[Bus.scala 125:73:@88.14]
  assign _GEN_108 = io_master_in_sync ? 1'h0 : _GEN_89; // @[Bus.scala 125:73:@88.14]
  assign _GEN_109 = io_master_in_sync ? 1'h0 : _GEN_90; // @[Bus.scala 125:73:@88.14]
  assign _GEN_110 = io_master_in_sync ? 1'h1 : _GEN_91; // @[Bus.scala 125:73:@88.14]
  assign _GEN_111 = io_master_in_sync ? 1'h0 : _GEN_92; // @[Bus.scala 125:73:@88.14]
  assign _GEN_112 = io_master_in_sync ? 1'h0 : _GEN_93; // @[Bus.scala 125:73:@88.14]
  assign _GEN_113 = io_master_in_sync ? 1'h0 : _GEN_94; // @[Bus.scala 125:73:@88.14]
  assign _GEN_114 = _T_104 ? _GEN_95 : _GEN_76; // @[Bus.scala 124:80:@87.12]
  assign _GEN_115 = _T_104 ? $signed(_GEN_96) : $signed(_GEN_77); // @[Bus.scala 124:80:@87.12]
  assign _GEN_116 = _T_104 ? $signed(_GEN_97) : $signed(_GEN_78); // @[Bus.scala 124:80:@87.12]
  assign _GEN_117 = _T_104 ? _GEN_98 : _GEN_79; // @[Bus.scala 124:80:@87.12]
  assign _GEN_120 = _T_104 ? $signed(_GEN_101) : $signed(_GEN_82); // @[Bus.scala 124:80:@87.12]
  assign _GEN_121 = _T_104 ? $signed(_GEN_102) : $signed(_GEN_83); // @[Bus.scala 124:80:@87.12]
  assign _GEN_122 = _T_104 ? _GEN_103 : _GEN_84; // @[Bus.scala 124:80:@87.12]
  assign _GEN_123 = _T_104 ? _GEN_104 : _GEN_85; // @[Bus.scala 124:80:@87.12]
  assign _GEN_124 = _T_104 ? _GEN_105 : _GEN_86; // @[Bus.scala 124:80:@87.12]
  assign _GEN_125 = _T_104 ? _GEN_106 : _GEN_87; // @[Bus.scala 124:80:@87.12]
  assign _GEN_126 = _T_104 ? _GEN_107 : _GEN_88; // @[Bus.scala 124:80:@87.12]
  assign _GEN_127 = _T_104 ? _GEN_108 : _GEN_89; // @[Bus.scala 124:80:@87.12]
  assign _GEN_128 = _T_104 ? _GEN_109 : _GEN_90; // @[Bus.scala 124:80:@87.12]
  assign _GEN_129 = _T_104 ? _GEN_110 : _GEN_91; // @[Bus.scala 124:80:@87.12]
  assign _GEN_130 = _T_104 ? _GEN_111 : _GEN_92; // @[Bus.scala 124:80:@87.12]
  assign _GEN_131 = _T_104 ? _GEN_112 : _GEN_93; // @[Bus.scala 124:80:@87.12]
  assign _GEN_132 = _T_104 ? _GEN_113 : _GEN_94; // @[Bus.scala 124:80:@87.12]
  assign _GEN_133 = _T_102 ? _GEN_114 : _GEN_76; // @[Bus.scala 123:72:@85.10]
  assign _GEN_134 = _T_102 ? $signed(_GEN_115) : $signed(_GEN_77); // @[Bus.scala 123:72:@85.10]
  assign _GEN_135 = _T_102 ? $signed(_GEN_116) : $signed(_GEN_78); // @[Bus.scala 123:72:@85.10]
  assign _GEN_136 = _T_102 ? _GEN_117 : _GEN_79; // @[Bus.scala 123:72:@85.10]
  assign _GEN_139 = _T_102 ? $signed(_GEN_120) : $signed(_GEN_82); // @[Bus.scala 123:72:@85.10]
  assign _GEN_140 = _T_102 ? $signed(_GEN_121) : $signed(_GEN_83); // @[Bus.scala 123:72:@85.10]
  assign _GEN_141 = _T_102 ? _GEN_122 : _GEN_84; // @[Bus.scala 123:72:@85.10]
  assign _GEN_142 = _T_102 ? _GEN_123 : _GEN_85; // @[Bus.scala 123:72:@85.10]
  assign _GEN_143 = _T_102 ? _GEN_124 : _GEN_86; // @[Bus.scala 123:72:@85.10]
  assign _GEN_144 = _T_102 ? _GEN_125 : _GEN_87; // @[Bus.scala 123:72:@85.10]
  assign _GEN_145 = _T_102 ? _GEN_126 : _GEN_88; // @[Bus.scala 123:72:@85.10]
  assign _GEN_146 = _T_102 ? _GEN_127 : _GEN_89; // @[Bus.scala 123:72:@85.10]
  assign _GEN_147 = _T_102 ? _GEN_128 : _GEN_90; // @[Bus.scala 123:72:@85.10]
  assign _GEN_148 = _T_102 ? _GEN_129 : _GEN_91; // @[Bus.scala 123:72:@85.10]
  assign _GEN_149 = _T_102 ? _GEN_130 : _GEN_92; // @[Bus.scala 123:72:@85.10]
  assign _GEN_150 = _T_102 ? _GEN_131 : _GEN_93; // @[Bus.scala 123:72:@85.10]
  assign _GEN_151 = _T_102 ? _GEN_132 : _GEN_94; // @[Bus.scala 123:72:@85.10]
  assign _GEN_152 = _T_98 ? _GEN_133 : _GEN_76; // @[Bus.scala 122:73:@83.8]
  assign _GEN_153 = _T_98 ? $signed(_GEN_134) : $signed(_GEN_77); // @[Bus.scala 122:73:@83.8]
  assign _GEN_154 = _T_98 ? $signed(_GEN_135) : $signed(_GEN_78); // @[Bus.scala 122:73:@83.8]
  assign _GEN_155 = _T_98 ? _GEN_136 : _GEN_79; // @[Bus.scala 122:73:@83.8]
  assign _GEN_158 = _T_98 ? $signed(_GEN_139) : $signed(_GEN_82); // @[Bus.scala 122:73:@83.8]
  assign _GEN_159 = _T_98 ? $signed(_GEN_140) : $signed(_GEN_83); // @[Bus.scala 122:73:@83.8]
  assign _GEN_160 = _T_98 ? _GEN_141 : _GEN_84; // @[Bus.scala 122:73:@83.8]
  assign _GEN_161 = _T_98 ? _GEN_142 : _GEN_85; // @[Bus.scala 122:73:@83.8]
  assign _GEN_162 = _T_98 ? _GEN_143 : _GEN_86; // @[Bus.scala 122:73:@83.8]
  assign _GEN_163 = _T_98 ? _GEN_144 : _GEN_87; // @[Bus.scala 122:73:@83.8]
  assign _GEN_164 = _T_98 ? _GEN_145 : _GEN_88; // @[Bus.scala 122:73:@83.8]
  assign _GEN_165 = _T_98 ? _GEN_146 : _GEN_89; // @[Bus.scala 122:73:@83.8]
  assign _GEN_166 = _T_98 ? _GEN_147 : _GEN_90; // @[Bus.scala 122:73:@83.8]
  assign _GEN_167 = _T_98 ? _GEN_148 : _GEN_91; // @[Bus.scala 122:73:@83.8]
  assign _GEN_168 = _T_98 ? _GEN_149 : _GEN_92; // @[Bus.scala 122:73:@83.8]
  assign _GEN_169 = _T_98 ? _GEN_150 : _GEN_93; // @[Bus.scala 122:73:@83.8]
  assign _GEN_170 = _T_98 ? _GEN_151 : _GEN_94; // @[Bus.scala 122:73:@83.8]
  assign _GEN_171 = _T_97 ? _GEN_152 : _GEN_76; // @[Bus.scala 121:41:@81.6]
  assign _GEN_172 = _T_97 ? $signed(_GEN_153) : $signed(_GEN_77); // @[Bus.scala 121:41:@81.6]
  assign _GEN_173 = _T_97 ? $signed(_GEN_154) : $signed(_GEN_78); // @[Bus.scala 121:41:@81.6]
  assign _GEN_174 = _T_97 ? _GEN_155 : _GEN_79; // @[Bus.scala 121:41:@81.6]
  assign _GEN_177 = _T_97 ? $signed(_GEN_158) : $signed(_GEN_82); // @[Bus.scala 121:41:@81.6]
  assign _GEN_178 = _T_97 ? $signed(_GEN_159) : $signed(_GEN_83); // @[Bus.scala 121:41:@81.6]
  assign _GEN_179 = _T_97 ? _GEN_160 : _GEN_84; // @[Bus.scala 121:41:@81.6]
  assign _GEN_180 = _T_97 ? _GEN_161 : _GEN_85; // @[Bus.scala 121:41:@81.6]
  assign _GEN_181 = _T_97 ? _GEN_162 : _GEN_86; // @[Bus.scala 121:41:@81.6]
  assign _GEN_182 = _T_97 ? _GEN_163 : _GEN_87; // @[Bus.scala 121:41:@81.6]
  assign _GEN_183 = _T_97 ? _GEN_164 : _GEN_88; // @[Bus.scala 121:41:@81.6]
  assign _GEN_184 = _T_97 ? _GEN_165 : _GEN_89; // @[Bus.scala 121:41:@81.6]
  assign _GEN_185 = _T_97 ? _GEN_166 : _GEN_90; // @[Bus.scala 121:41:@81.6]
  assign _GEN_186 = _T_97 ? _GEN_167 : _GEN_91; // @[Bus.scala 121:41:@81.6]
  assign _GEN_187 = _T_97 ? _GEN_168 : _GEN_92; // @[Bus.scala 121:41:@81.6]
  assign _GEN_188 = _T_97 ? _GEN_169 : _GEN_93; // @[Bus.scala 121:41:@81.6]
  assign _GEN_189 = _T_97 ? _GEN_170 : _GEN_94; // @[Bus.scala 121:41:@81.6]
  assign _T_138 = $signed(32'sh8) <= $signed(io_master_in_addr); // @[Bus.scala 152:88:@118.10]
  assign _T_140 = _T_138 == 1'h0; // @[Bus.scala 152:76:@119.10]
  assign _T_141 = _T_102 & _T_140; // @[Bus.scala 152:73:@120.10]
  assign _T_143 = _T_141 == 1'h0; // @[Bus.scala 152:38:@121.10]
  assign _T_145 = $signed(io_master_in_addr) >= $signed(32'sh8); // @[Bus.scala 153:67:@123.12]
  assign _T_147 = $signed(32'sh10) <= $signed(io_master_in_addr); // @[Bus.scala 153:97:@124.12]
  assign _T_149 = _T_147 == 1'h0; // @[Bus.scala 153:84:@125.12]
  assign _T_150 = _T_145 & _T_149; // @[Bus.scala 153:81:@126.12]
  assign _T_152 = _T_150 == 1'h0; // @[Bus.scala 153:46:@127.12]
  assign _T_154 = $signed(io_master_in_addr) >= $signed(32'sh10); // @[Bus.scala 154:75:@129.14]
  assign _T_156 = $signed(32'sh18) <= $signed(io_master_in_addr); // @[Bus.scala 154:106:@130.14]
  assign _T_158 = _T_156 == 1'h0; // @[Bus.scala 154:93:@131.14]
  assign _T_159 = _T_154 & _T_158; // @[Bus.scala 154:90:@132.14]
  assign _T_161 = _T_159 == 1'h0; // @[Bus.scala 154:54:@133.14]
  assign _T_163 = $signed(io_master_in_addr) >= $signed(32'sh18); // @[Bus.scala 155:83:@135.16]
  assign _T_165 = $signed(32'sh20) <= $signed(io_master_in_addr); // @[Bus.scala 155:114:@136.16]
  assign _T_167 = _T_165 == 1'h0; // @[Bus.scala 155:101:@137.16]
  assign _T_168 = _T_163 & _T_167; // @[Bus.scala 155:98:@138.16]
  assign _T_170 = _T_168 == 1'h0; // @[Bus.scala 155:62:@139.16]
  assign _GEN_190 = io_master_in_sync ? 4'h3 : _GEN_171; // @[Bus.scala 156:89:@141.18]
  assign _GEN_191 = io_master_in_sync ? 32'h0 : master_out_r_ack; // @[Bus.scala 156:89:@141.18]
  assign _GEN_192 = io_master_in_sync ? $signed(32'sh0) : $signed(master_out_r_data); // @[Bus.scala 156:89:@141.18]
  assign _GEN_193 = io_master_in_sync ? $signed(io_master_in_addr) : $signed(_GEN_172); // @[Bus.scala 156:89:@141.18]
  assign _GEN_194 = io_master_in_sync ? $signed(32'sh0) : $signed(_GEN_173); // @[Bus.scala 156:89:@141.18]
  assign _GEN_195 = io_master_in_sync ? io_master_in_trans_type : _GEN_174; // @[Bus.scala 156:89:@141.18]
  assign _GEN_196 = io_master_in_sync ? 32'h0 : resp_signal_r_ack; // @[Bus.scala 156:89:@141.18]
  assign _GEN_197 = io_master_in_sync ? $signed(32'sh0) : $signed(resp_signal_r_data); // @[Bus.scala 156:89:@141.18]
  assign _GEN_198 = io_master_in_sync ? 1'h0 : _GEN_180; // @[Bus.scala 156:89:@141.18]
  assign _GEN_199 = io_master_in_sync ? 1'h1 : _GEN_181; // @[Bus.scala 156:89:@141.18]
  assign _GEN_200 = io_master_in_sync ? 1'h0 : _GEN_182; // @[Bus.scala 156:89:@141.18]
  assign _GEN_201 = io_master_in_sync ? 1'h0 : _GEN_183; // @[Bus.scala 156:89:@141.18]
  assign _GEN_202 = io_master_in_sync ? 1'h0 : _GEN_184; // @[Bus.scala 156:89:@141.18]
  assign _GEN_203 = io_master_in_sync ? 1'h0 : _GEN_185; // @[Bus.scala 156:89:@141.18]
  assign _GEN_204 = io_master_in_sync ? 1'h0 : _GEN_186; // @[Bus.scala 156:89:@141.18]
  assign _GEN_205 = io_master_in_sync ? 1'h0 : _GEN_187; // @[Bus.scala 156:89:@141.18]
  assign _GEN_206 = io_master_in_sync ? 1'h0 : _GEN_188; // @[Bus.scala 156:89:@141.18]
  assign _GEN_207 = io_master_in_sync ? 1'h0 : _GEN_189; // @[Bus.scala 156:89:@141.18]
  assign _GEN_208 = _T_170 ? _GEN_190 : _GEN_171; // @[Bus.scala 155:138:@140.16]
  assign _GEN_209 = _T_170 ? _GEN_191 : master_out_r_ack; // @[Bus.scala 155:138:@140.16]
  assign _GEN_210 = _T_170 ? $signed(_GEN_192) : $signed(master_out_r_data); // @[Bus.scala 155:138:@140.16]
  assign _GEN_211 = _T_170 ? $signed(_GEN_193) : $signed(_GEN_172); // @[Bus.scala 155:138:@140.16]
  assign _GEN_212 = _T_170 ? $signed(_GEN_194) : $signed(_GEN_173); // @[Bus.scala 155:138:@140.16]
  assign _GEN_213 = _T_170 ? _GEN_195 : _GEN_174; // @[Bus.scala 155:138:@140.16]
  assign _GEN_214 = _T_170 ? _GEN_196 : resp_signal_r_ack; // @[Bus.scala 155:138:@140.16]
  assign _GEN_215 = _T_170 ? $signed(_GEN_197) : $signed(resp_signal_r_data); // @[Bus.scala 155:138:@140.16]
  assign _GEN_216 = _T_170 ? _GEN_198 : _GEN_180; // @[Bus.scala 155:138:@140.16]
  assign _GEN_217 = _T_170 ? _GEN_199 : _GEN_181; // @[Bus.scala 155:138:@140.16]
  assign _GEN_218 = _T_170 ? _GEN_200 : _GEN_182; // @[Bus.scala 155:138:@140.16]
  assign _GEN_219 = _T_170 ? _GEN_201 : _GEN_183; // @[Bus.scala 155:138:@140.16]
  assign _GEN_220 = _T_170 ? _GEN_202 : _GEN_184; // @[Bus.scala 155:138:@140.16]
  assign _GEN_221 = _T_170 ? _GEN_203 : _GEN_185; // @[Bus.scala 155:138:@140.16]
  assign _GEN_222 = _T_170 ? _GEN_204 : _GEN_186; // @[Bus.scala 155:138:@140.16]
  assign _GEN_223 = _T_170 ? _GEN_205 : _GEN_187; // @[Bus.scala 155:138:@140.16]
  assign _GEN_224 = _T_170 ? _GEN_206 : _GEN_188; // @[Bus.scala 155:138:@140.16]
  assign _GEN_225 = _T_170 ? _GEN_207 : _GEN_189; // @[Bus.scala 155:138:@140.16]
  assign _GEN_226 = _T_161 ? _GEN_208 : _GEN_171; // @[Bus.scala 154:130:@134.14]
  assign _GEN_227 = _T_161 ? _GEN_209 : master_out_r_ack; // @[Bus.scala 154:130:@134.14]
  assign _GEN_228 = _T_161 ? $signed(_GEN_210) : $signed(master_out_r_data); // @[Bus.scala 154:130:@134.14]
  assign _GEN_229 = _T_161 ? $signed(_GEN_211) : $signed(_GEN_172); // @[Bus.scala 154:130:@134.14]
  assign _GEN_230 = _T_161 ? $signed(_GEN_212) : $signed(_GEN_173); // @[Bus.scala 154:130:@134.14]
  assign _GEN_231 = _T_161 ? _GEN_213 : _GEN_174; // @[Bus.scala 154:130:@134.14]
  assign _GEN_232 = _T_161 ? _GEN_214 : resp_signal_r_ack; // @[Bus.scala 154:130:@134.14]
  assign _GEN_233 = _T_161 ? $signed(_GEN_215) : $signed(resp_signal_r_data); // @[Bus.scala 154:130:@134.14]
  assign _GEN_234 = _T_161 ? _GEN_216 : _GEN_180; // @[Bus.scala 154:130:@134.14]
  assign _GEN_235 = _T_161 ? _GEN_217 : _GEN_181; // @[Bus.scala 154:130:@134.14]
  assign _GEN_236 = _T_161 ? _GEN_218 : _GEN_182; // @[Bus.scala 154:130:@134.14]
  assign _GEN_237 = _T_161 ? _GEN_219 : _GEN_183; // @[Bus.scala 154:130:@134.14]
  assign _GEN_238 = _T_161 ? _GEN_220 : _GEN_184; // @[Bus.scala 154:130:@134.14]
  assign _GEN_239 = _T_161 ? _GEN_221 : _GEN_185; // @[Bus.scala 154:130:@134.14]
  assign _GEN_240 = _T_161 ? _GEN_222 : _GEN_186; // @[Bus.scala 154:130:@134.14]
  assign _GEN_241 = _T_161 ? _GEN_223 : _GEN_187; // @[Bus.scala 154:130:@134.14]
  assign _GEN_242 = _T_161 ? _GEN_224 : _GEN_188; // @[Bus.scala 154:130:@134.14]
  assign _GEN_243 = _T_161 ? _GEN_225 : _GEN_189; // @[Bus.scala 154:130:@134.14]
  assign _GEN_244 = _T_152 ? _GEN_226 : _GEN_171; // @[Bus.scala 153:121:@128.12]
  assign _GEN_245 = _T_152 ? _GEN_227 : master_out_r_ack; // @[Bus.scala 153:121:@128.12]
  assign _GEN_246 = _T_152 ? $signed(_GEN_228) : $signed(master_out_r_data); // @[Bus.scala 153:121:@128.12]
  assign _GEN_247 = _T_152 ? $signed(_GEN_229) : $signed(_GEN_172); // @[Bus.scala 153:121:@128.12]
  assign _GEN_248 = _T_152 ? $signed(_GEN_230) : $signed(_GEN_173); // @[Bus.scala 153:121:@128.12]
  assign _GEN_249 = _T_152 ? _GEN_231 : _GEN_174; // @[Bus.scala 153:121:@128.12]
  assign _GEN_250 = _T_152 ? _GEN_232 : resp_signal_r_ack; // @[Bus.scala 153:121:@128.12]
  assign _GEN_251 = _T_152 ? $signed(_GEN_233) : $signed(resp_signal_r_data); // @[Bus.scala 153:121:@128.12]
  assign _GEN_252 = _T_152 ? _GEN_234 : _GEN_180; // @[Bus.scala 153:121:@128.12]
  assign _GEN_253 = _T_152 ? _GEN_235 : _GEN_181; // @[Bus.scala 153:121:@128.12]
  assign _GEN_254 = _T_152 ? _GEN_236 : _GEN_182; // @[Bus.scala 153:121:@128.12]
  assign _GEN_255 = _T_152 ? _GEN_237 : _GEN_183; // @[Bus.scala 153:121:@128.12]
  assign _GEN_256 = _T_152 ? _GEN_238 : _GEN_184; // @[Bus.scala 153:121:@128.12]
  assign _GEN_257 = _T_152 ? _GEN_239 : _GEN_185; // @[Bus.scala 153:121:@128.12]
  assign _GEN_258 = _T_152 ? _GEN_240 : _GEN_186; // @[Bus.scala 153:121:@128.12]
  assign _GEN_259 = _T_152 ? _GEN_241 : _GEN_187; // @[Bus.scala 153:121:@128.12]
  assign _GEN_260 = _T_152 ? _GEN_242 : _GEN_188; // @[Bus.scala 153:121:@128.12]
  assign _GEN_261 = _T_152 ? _GEN_243 : _GEN_189; // @[Bus.scala 153:121:@128.12]
  assign _GEN_262 = _T_143 ? _GEN_244 : _GEN_171; // @[Bus.scala 152:112:@122.10]
  assign _GEN_263 = _T_143 ? _GEN_245 : master_out_r_ack; // @[Bus.scala 152:112:@122.10]
  assign _GEN_264 = _T_143 ? $signed(_GEN_246) : $signed(master_out_r_data); // @[Bus.scala 152:112:@122.10]
  assign _GEN_265 = _T_143 ? $signed(_GEN_247) : $signed(_GEN_172); // @[Bus.scala 152:112:@122.10]
  assign _GEN_266 = _T_143 ? $signed(_GEN_248) : $signed(_GEN_173); // @[Bus.scala 152:112:@122.10]
  assign _GEN_267 = _T_143 ? _GEN_249 : _GEN_174; // @[Bus.scala 152:112:@122.10]
  assign _GEN_268 = _T_143 ? _GEN_250 : resp_signal_r_ack; // @[Bus.scala 152:112:@122.10]
  assign _GEN_269 = _T_143 ? $signed(_GEN_251) : $signed(resp_signal_r_data); // @[Bus.scala 152:112:@122.10]
  assign _GEN_270 = _T_143 ? _GEN_252 : _GEN_180; // @[Bus.scala 152:112:@122.10]
  assign _GEN_271 = _T_143 ? _GEN_253 : _GEN_181; // @[Bus.scala 152:112:@122.10]
  assign _GEN_272 = _T_143 ? _GEN_254 : _GEN_182; // @[Bus.scala 152:112:@122.10]
  assign _GEN_273 = _T_143 ? _GEN_255 : _GEN_183; // @[Bus.scala 152:112:@122.10]
  assign _GEN_274 = _T_143 ? _GEN_256 : _GEN_184; // @[Bus.scala 152:112:@122.10]
  assign _GEN_275 = _T_143 ? _GEN_257 : _GEN_185; // @[Bus.scala 152:112:@122.10]
  assign _GEN_276 = _T_143 ? _GEN_258 : _GEN_186; // @[Bus.scala 152:112:@122.10]
  assign _GEN_277 = _T_143 ? _GEN_259 : _GEN_187; // @[Bus.scala 152:112:@122.10]
  assign _GEN_278 = _T_143 ? _GEN_260 : _GEN_188; // @[Bus.scala 152:112:@122.10]
  assign _GEN_279 = _T_143 ? _GEN_261 : _GEN_189; // @[Bus.scala 152:112:@122.10]
  assign _GEN_280 = _T_98 ? _GEN_262 : _GEN_171; // @[Bus.scala 151:73:@116.8]
  assign _GEN_281 = _T_98 ? _GEN_263 : master_out_r_ack; // @[Bus.scala 151:73:@116.8]
  assign _GEN_282 = _T_98 ? $signed(_GEN_264) : $signed(master_out_r_data); // @[Bus.scala 151:73:@116.8]
  assign _GEN_283 = _T_98 ? $signed(_GEN_265) : $signed(_GEN_172); // @[Bus.scala 151:73:@116.8]
  assign _GEN_284 = _T_98 ? $signed(_GEN_266) : $signed(_GEN_173); // @[Bus.scala 151:73:@116.8]
  assign _GEN_285 = _T_98 ? _GEN_267 : _GEN_174; // @[Bus.scala 151:73:@116.8]
  assign _GEN_286 = _T_98 ? _GEN_268 : resp_signal_r_ack; // @[Bus.scala 151:73:@116.8]
  assign _GEN_287 = _T_98 ? $signed(_GEN_269) : $signed(resp_signal_r_data); // @[Bus.scala 151:73:@116.8]
  assign _GEN_288 = _T_98 ? _GEN_270 : _GEN_180; // @[Bus.scala 151:73:@116.8]
  assign _GEN_289 = _T_98 ? _GEN_271 : _GEN_181; // @[Bus.scala 151:73:@116.8]
  assign _GEN_290 = _T_98 ? _GEN_272 : _GEN_182; // @[Bus.scala 151:73:@116.8]
  assign _GEN_291 = _T_98 ? _GEN_273 : _GEN_183; // @[Bus.scala 151:73:@116.8]
  assign _GEN_292 = _T_98 ? _GEN_274 : _GEN_184; // @[Bus.scala 151:73:@116.8]
  assign _GEN_293 = _T_98 ? _GEN_275 : _GEN_185; // @[Bus.scala 151:73:@116.8]
  assign _GEN_294 = _T_98 ? _GEN_276 : _GEN_186; // @[Bus.scala 151:73:@116.8]
  assign _GEN_295 = _T_98 ? _GEN_277 : _GEN_187; // @[Bus.scala 151:73:@116.8]
  assign _GEN_296 = _T_98 ? _GEN_278 : _GEN_188; // @[Bus.scala 151:73:@116.8]
  assign _GEN_297 = _T_98 ? _GEN_279 : _GEN_189; // @[Bus.scala 151:73:@116.8]
  assign _GEN_298 = _T_97 ? _GEN_280 : _GEN_171; // @[Bus.scala 150:41:@114.6]
  assign _GEN_299 = _T_97 ? _GEN_281 : master_out_r_ack; // @[Bus.scala 150:41:@114.6]
  assign _GEN_300 = _T_97 ? $signed(_GEN_282) : $signed(master_out_r_data); // @[Bus.scala 150:41:@114.6]
  assign _GEN_301 = _T_97 ? $signed(_GEN_283) : $signed(_GEN_172); // @[Bus.scala 150:41:@114.6]
  assign _GEN_302 = _T_97 ? $signed(_GEN_284) : $signed(_GEN_173); // @[Bus.scala 150:41:@114.6]
  assign _GEN_303 = _T_97 ? _GEN_285 : _GEN_174; // @[Bus.scala 150:41:@114.6]
  assign _GEN_304 = _T_97 ? _GEN_286 : resp_signal_r_ack; // @[Bus.scala 150:41:@114.6]
  assign _GEN_305 = _T_97 ? $signed(_GEN_287) : $signed(resp_signal_r_data); // @[Bus.scala 150:41:@114.6]
  assign _GEN_306 = _T_97 ? _GEN_288 : _GEN_180; // @[Bus.scala 150:41:@114.6]
  assign _GEN_307 = _T_97 ? _GEN_289 : _GEN_181; // @[Bus.scala 150:41:@114.6]
  assign _GEN_308 = _T_97 ? _GEN_290 : _GEN_182; // @[Bus.scala 150:41:@114.6]
  assign _GEN_309 = _T_97 ? _GEN_291 : _GEN_183; // @[Bus.scala 150:41:@114.6]
  assign _GEN_310 = _T_97 ? _GEN_292 : _GEN_184; // @[Bus.scala 150:41:@114.6]
  assign _GEN_311 = _T_97 ? _GEN_293 : _GEN_185; // @[Bus.scala 150:41:@114.6]
  assign _GEN_312 = _T_97 ? _GEN_294 : _GEN_186; // @[Bus.scala 150:41:@114.6]
  assign _GEN_313 = _T_97 ? _GEN_295 : _GEN_187; // @[Bus.scala 150:41:@114.6]
  assign _GEN_314 = _T_97 ? _GEN_296 : _GEN_188; // @[Bus.scala 150:41:@114.6]
  assign _GEN_315 = _T_97 ? _GEN_297 : _GEN_189; // @[Bus.scala 150:41:@114.6]
  assign _T_221 = 32'h1 == io_master_in_trans_type; // @[Bus.scala 187:76:@193.16]
  assign _GEN_316 = io_master_in_sync ? 4'h3 : _GEN_298; // @[Bus.scala 188:89:@195.18]
  assign _GEN_317 = io_master_in_sync ? 32'h0 : _GEN_299; // @[Bus.scala 188:89:@195.18]
  assign _GEN_318 = io_master_in_sync ? $signed(32'sh0) : $signed(_GEN_300); // @[Bus.scala 188:89:@195.18]
  assign _GEN_319 = io_master_in_sync ? $signed(io_master_in_addr) : $signed(_GEN_301); // @[Bus.scala 188:89:@195.18]
  assign _GEN_320 = io_master_in_sync ? $signed(io_master_in_data) : $signed(_GEN_302); // @[Bus.scala 188:89:@195.18]
  assign _GEN_321 = io_master_in_sync ? io_master_in_trans_type : _GEN_303; // @[Bus.scala 188:89:@195.18]
  assign _GEN_322 = io_master_in_sync ? 32'h0 : _GEN_304; // @[Bus.scala 188:89:@195.18]
  assign _GEN_323 = io_master_in_sync ? $signed(32'sh0) : $signed(_GEN_305); // @[Bus.scala 188:89:@195.18]
  assign _GEN_324 = io_master_in_sync ? 1'h0 : _GEN_306; // @[Bus.scala 188:89:@195.18]
  assign _GEN_325 = io_master_in_sync ? 1'h1 : _GEN_307; // @[Bus.scala 188:89:@195.18]
  assign _GEN_326 = io_master_in_sync ? 1'h0 : _GEN_308; // @[Bus.scala 188:89:@195.18]
  assign _GEN_327 = io_master_in_sync ? 1'h0 : _GEN_309; // @[Bus.scala 188:89:@195.18]
  assign _GEN_328 = io_master_in_sync ? 1'h0 : _GEN_310; // @[Bus.scala 188:89:@195.18]
  assign _GEN_329 = io_master_in_sync ? 1'h0 : _GEN_311; // @[Bus.scala 188:89:@195.18]
  assign _GEN_330 = io_master_in_sync ? 1'h0 : _GEN_312; // @[Bus.scala 188:89:@195.18]
  assign _GEN_331 = io_master_in_sync ? 1'h0 : _GEN_313; // @[Bus.scala 188:89:@195.18]
  assign _GEN_332 = io_master_in_sync ? 1'h0 : _GEN_314; // @[Bus.scala 188:89:@195.18]
  assign _GEN_333 = io_master_in_sync ? 1'h0 : _GEN_315; // @[Bus.scala 188:89:@195.18]
  assign _GEN_334 = _T_221 ? _GEN_316 : _GEN_298; // @[Bus.scala 187:106:@194.16]
  assign _GEN_335 = _T_221 ? _GEN_317 : _GEN_299; // @[Bus.scala 187:106:@194.16]
  assign _GEN_336 = _T_221 ? $signed(_GEN_318) : $signed(_GEN_300); // @[Bus.scala 187:106:@194.16]
  assign _GEN_337 = _T_221 ? $signed(_GEN_319) : $signed(_GEN_301); // @[Bus.scala 187:106:@194.16]
  assign _GEN_338 = _T_221 ? $signed(_GEN_320) : $signed(_GEN_302); // @[Bus.scala 187:106:@194.16]
  assign _GEN_339 = _T_221 ? _GEN_321 : _GEN_303; // @[Bus.scala 187:106:@194.16]
  assign _GEN_340 = _T_221 ? _GEN_322 : _GEN_304; // @[Bus.scala 187:106:@194.16]
  assign _GEN_341 = _T_221 ? $signed(_GEN_323) : $signed(_GEN_305); // @[Bus.scala 187:106:@194.16]
  assign _GEN_342 = _T_221 ? _GEN_324 : _GEN_306; // @[Bus.scala 187:106:@194.16]
  assign _GEN_343 = _T_221 ? _GEN_325 : _GEN_307; // @[Bus.scala 187:106:@194.16]
  assign _GEN_344 = _T_221 ? _GEN_326 : _GEN_308; // @[Bus.scala 187:106:@194.16]
  assign _GEN_345 = _T_221 ? _GEN_327 : _GEN_309; // @[Bus.scala 187:106:@194.16]
  assign _GEN_346 = _T_221 ? _GEN_328 : _GEN_310; // @[Bus.scala 187:106:@194.16]
  assign _GEN_347 = _T_221 ? _GEN_329 : _GEN_311; // @[Bus.scala 187:106:@194.16]
  assign _GEN_348 = _T_221 ? _GEN_330 : _GEN_312; // @[Bus.scala 187:106:@194.16]
  assign _GEN_349 = _T_221 ? _GEN_331 : _GEN_313; // @[Bus.scala 187:106:@194.16]
  assign _GEN_350 = _T_221 ? _GEN_332 : _GEN_314; // @[Bus.scala 187:106:@194.16]
  assign _GEN_351 = _T_221 ? _GEN_333 : _GEN_315; // @[Bus.scala 187:106:@194.16]
  assign _GEN_352 = _T_170 ? _GEN_334 : _GEN_298; // @[Bus.scala 186:130:@192.14]
  assign _GEN_353 = _T_170 ? _GEN_335 : _GEN_299; // @[Bus.scala 186:130:@192.14]
  assign _GEN_354 = _T_170 ? $signed(_GEN_336) : $signed(_GEN_300); // @[Bus.scala 186:130:@192.14]
  assign _GEN_355 = _T_170 ? $signed(_GEN_337) : $signed(_GEN_301); // @[Bus.scala 186:130:@192.14]
  assign _GEN_356 = _T_170 ? $signed(_GEN_338) : $signed(_GEN_302); // @[Bus.scala 186:130:@192.14]
  assign _GEN_357 = _T_170 ? _GEN_339 : _GEN_303; // @[Bus.scala 186:130:@192.14]
  assign _GEN_358 = _T_170 ? _GEN_340 : _GEN_304; // @[Bus.scala 186:130:@192.14]
  assign _GEN_359 = _T_170 ? $signed(_GEN_341) : $signed(_GEN_305); // @[Bus.scala 186:130:@192.14]
  assign _GEN_360 = _T_170 ? _GEN_342 : _GEN_306; // @[Bus.scala 186:130:@192.14]
  assign _GEN_361 = _T_170 ? _GEN_343 : _GEN_307; // @[Bus.scala 186:130:@192.14]
  assign _GEN_362 = _T_170 ? _GEN_344 : _GEN_308; // @[Bus.scala 186:130:@192.14]
  assign _GEN_363 = _T_170 ? _GEN_345 : _GEN_309; // @[Bus.scala 186:130:@192.14]
  assign _GEN_364 = _T_170 ? _GEN_346 : _GEN_310; // @[Bus.scala 186:130:@192.14]
  assign _GEN_365 = _T_170 ? _GEN_347 : _GEN_311; // @[Bus.scala 186:130:@192.14]
  assign _GEN_366 = _T_170 ? _GEN_348 : _GEN_312; // @[Bus.scala 186:130:@192.14]
  assign _GEN_367 = _T_170 ? _GEN_349 : _GEN_313; // @[Bus.scala 186:130:@192.14]
  assign _GEN_368 = _T_170 ? _GEN_350 : _GEN_314; // @[Bus.scala 186:130:@192.14]
  assign _GEN_369 = _T_170 ? _GEN_351 : _GEN_315; // @[Bus.scala 186:130:@192.14]
  assign _GEN_370 = _T_161 ? _GEN_352 : _GEN_298; // @[Bus.scala 185:122:@186.12]
  assign _GEN_371 = _T_161 ? _GEN_353 : _GEN_299; // @[Bus.scala 185:122:@186.12]
  assign _GEN_372 = _T_161 ? $signed(_GEN_354) : $signed(_GEN_300); // @[Bus.scala 185:122:@186.12]
  assign _GEN_373 = _T_161 ? $signed(_GEN_355) : $signed(_GEN_301); // @[Bus.scala 185:122:@186.12]
  assign _GEN_374 = _T_161 ? $signed(_GEN_356) : $signed(_GEN_302); // @[Bus.scala 185:122:@186.12]
  assign _GEN_375 = _T_161 ? _GEN_357 : _GEN_303; // @[Bus.scala 185:122:@186.12]
  assign _GEN_376 = _T_161 ? _GEN_358 : _GEN_304; // @[Bus.scala 185:122:@186.12]
  assign _GEN_377 = _T_161 ? $signed(_GEN_359) : $signed(_GEN_305); // @[Bus.scala 185:122:@186.12]
  assign _GEN_378 = _T_161 ? _GEN_360 : _GEN_306; // @[Bus.scala 185:122:@186.12]
  assign _GEN_379 = _T_161 ? _GEN_361 : _GEN_307; // @[Bus.scala 185:122:@186.12]
  assign _GEN_380 = _T_161 ? _GEN_362 : _GEN_308; // @[Bus.scala 185:122:@186.12]
  assign _GEN_381 = _T_161 ? _GEN_363 : _GEN_309; // @[Bus.scala 185:122:@186.12]
  assign _GEN_382 = _T_161 ? _GEN_364 : _GEN_310; // @[Bus.scala 185:122:@186.12]
  assign _GEN_383 = _T_161 ? _GEN_365 : _GEN_311; // @[Bus.scala 185:122:@186.12]
  assign _GEN_384 = _T_161 ? _GEN_366 : _GEN_312; // @[Bus.scala 185:122:@186.12]
  assign _GEN_385 = _T_161 ? _GEN_367 : _GEN_313; // @[Bus.scala 185:122:@186.12]
  assign _GEN_386 = _T_161 ? _GEN_368 : _GEN_314; // @[Bus.scala 185:122:@186.12]
  assign _GEN_387 = _T_161 ? _GEN_369 : _GEN_315; // @[Bus.scala 185:122:@186.12]
  assign _GEN_388 = _T_152 ? _GEN_370 : _GEN_298; // @[Bus.scala 184:113:@180.10]
  assign _GEN_389 = _T_152 ? _GEN_371 : _GEN_299; // @[Bus.scala 184:113:@180.10]
  assign _GEN_390 = _T_152 ? $signed(_GEN_372) : $signed(_GEN_300); // @[Bus.scala 184:113:@180.10]
  assign _GEN_391 = _T_152 ? $signed(_GEN_373) : $signed(_GEN_301); // @[Bus.scala 184:113:@180.10]
  assign _GEN_392 = _T_152 ? $signed(_GEN_374) : $signed(_GEN_302); // @[Bus.scala 184:113:@180.10]
  assign _GEN_393 = _T_152 ? _GEN_375 : _GEN_303; // @[Bus.scala 184:113:@180.10]
  assign _GEN_394 = _T_152 ? _GEN_376 : _GEN_304; // @[Bus.scala 184:113:@180.10]
  assign _GEN_395 = _T_152 ? $signed(_GEN_377) : $signed(_GEN_305); // @[Bus.scala 184:113:@180.10]
  assign _GEN_396 = _T_152 ? _GEN_378 : _GEN_306; // @[Bus.scala 184:113:@180.10]
  assign _GEN_397 = _T_152 ? _GEN_379 : _GEN_307; // @[Bus.scala 184:113:@180.10]
  assign _GEN_398 = _T_152 ? _GEN_380 : _GEN_308; // @[Bus.scala 184:113:@180.10]
  assign _GEN_399 = _T_152 ? _GEN_381 : _GEN_309; // @[Bus.scala 184:113:@180.10]
  assign _GEN_400 = _T_152 ? _GEN_382 : _GEN_310; // @[Bus.scala 184:113:@180.10]
  assign _GEN_401 = _T_152 ? _GEN_383 : _GEN_311; // @[Bus.scala 184:113:@180.10]
  assign _GEN_402 = _T_152 ? _GEN_384 : _GEN_312; // @[Bus.scala 184:113:@180.10]
  assign _GEN_403 = _T_152 ? _GEN_385 : _GEN_313; // @[Bus.scala 184:113:@180.10]
  assign _GEN_404 = _T_152 ? _GEN_386 : _GEN_314; // @[Bus.scala 184:113:@180.10]
  assign _GEN_405 = _T_152 ? _GEN_387 : _GEN_315; // @[Bus.scala 184:113:@180.10]
  assign _GEN_406 = _T_143 ? _GEN_388 : _GEN_298; // @[Bus.scala 183:104:@174.8]
  assign _GEN_407 = _T_143 ? _GEN_389 : _GEN_299; // @[Bus.scala 183:104:@174.8]
  assign _GEN_408 = _T_143 ? $signed(_GEN_390) : $signed(_GEN_300); // @[Bus.scala 183:104:@174.8]
  assign _GEN_409 = _T_143 ? $signed(_GEN_391) : $signed(_GEN_301); // @[Bus.scala 183:104:@174.8]
  assign _GEN_410 = _T_143 ? $signed(_GEN_392) : $signed(_GEN_302); // @[Bus.scala 183:104:@174.8]
  assign _GEN_411 = _T_143 ? _GEN_393 : _GEN_303; // @[Bus.scala 183:104:@174.8]
  assign _GEN_412 = _T_143 ? _GEN_394 : _GEN_304; // @[Bus.scala 183:104:@174.8]
  assign _GEN_413 = _T_143 ? $signed(_GEN_395) : $signed(_GEN_305); // @[Bus.scala 183:104:@174.8]
  assign _GEN_414 = _T_143 ? _GEN_396 : _GEN_306; // @[Bus.scala 183:104:@174.8]
  assign _GEN_415 = _T_143 ? _GEN_397 : _GEN_307; // @[Bus.scala 183:104:@174.8]
  assign _GEN_416 = _T_143 ? _GEN_398 : _GEN_308; // @[Bus.scala 183:104:@174.8]
  assign _GEN_417 = _T_143 ? _GEN_399 : _GEN_309; // @[Bus.scala 183:104:@174.8]
  assign _GEN_418 = _T_143 ? _GEN_400 : _GEN_310; // @[Bus.scala 183:104:@174.8]
  assign _GEN_419 = _T_143 ? _GEN_401 : _GEN_311; // @[Bus.scala 183:104:@174.8]
  assign _GEN_420 = _T_143 ? _GEN_402 : _GEN_312; // @[Bus.scala 183:104:@174.8]
  assign _GEN_421 = _T_143 ? _GEN_403 : _GEN_313; // @[Bus.scala 183:104:@174.8]
  assign _GEN_422 = _T_143 ? _GEN_404 : _GEN_314; // @[Bus.scala 183:104:@174.8]
  assign _GEN_423 = _T_143 ? _GEN_405 : _GEN_315; // @[Bus.scala 183:104:@174.8]
  assign _GEN_424 = _T_97 ? _GEN_406 : _GEN_298; // @[Bus.scala 182:41:@168.6]
  assign _GEN_425 = _T_97 ? _GEN_407 : _GEN_299; // @[Bus.scala 182:41:@168.6]
  assign _GEN_426 = _T_97 ? $signed(_GEN_408) : $signed(_GEN_300); // @[Bus.scala 182:41:@168.6]
  assign _GEN_427 = _T_97 ? $signed(_GEN_409) : $signed(_GEN_301); // @[Bus.scala 182:41:@168.6]
  assign _GEN_428 = _T_97 ? $signed(_GEN_410) : $signed(_GEN_302); // @[Bus.scala 182:41:@168.6]
  assign _GEN_429 = _T_97 ? _GEN_411 : _GEN_303; // @[Bus.scala 182:41:@168.6]
  assign _GEN_430 = _T_97 ? _GEN_412 : _GEN_304; // @[Bus.scala 182:41:@168.6]
  assign _GEN_431 = _T_97 ? $signed(_GEN_413) : $signed(_GEN_305); // @[Bus.scala 182:41:@168.6]
  assign _GEN_432 = _T_97 ? _GEN_414 : _GEN_306; // @[Bus.scala 182:41:@168.6]
  assign _GEN_433 = _T_97 ? _GEN_415 : _GEN_307; // @[Bus.scala 182:41:@168.6]
  assign _GEN_434 = _T_97 ? _GEN_416 : _GEN_308; // @[Bus.scala 182:41:@168.6]
  assign _GEN_435 = _T_97 ? _GEN_417 : _GEN_309; // @[Bus.scala 182:41:@168.6]
  assign _GEN_436 = _T_97 ? _GEN_418 : _GEN_310; // @[Bus.scala 182:41:@168.6]
  assign _GEN_437 = _T_97 ? _GEN_419 : _GEN_311; // @[Bus.scala 182:41:@168.6]
  assign _GEN_438 = _T_97 ? _GEN_420 : _GEN_312; // @[Bus.scala 182:41:@168.6]
  assign _GEN_439 = _T_97 ? _GEN_421 : _GEN_313; // @[Bus.scala 182:41:@168.6]
  assign _GEN_440 = _T_97 ? _GEN_422 : _GEN_314; // @[Bus.scala 182:41:@168.6]
  assign _GEN_441 = _T_97 ? _GEN_423 : _GEN_315; // @[Bus.scala 182:41:@168.6]
  assign _T_241 = $signed(io_master_in_addr) <= $signed(32'shf); // @[Bus.scala 217:65:@228.12]
  assign _T_243 = $signed(-32'sh8) + $signed(io_master_in_addr); // @[Bus.scala 220:92:@232.16]
  assign _T_244 = $signed(-32'sh8) + $signed(io_master_in_addr); // @[Bus.scala 220:92:@233.16]
  assign _T_245 = $signed(_T_244); // @[Bus.scala 220:92:@234.16]
  assign _GEN_442 = io_master_in_sync ? 4'h4 : _GEN_424; // @[Bus.scala 218:73:@230.14]
  assign _GEN_443 = io_master_in_sync ? $signed(_T_245) : $signed(_GEN_427); // @[Bus.scala 218:73:@230.14]
  assign _GEN_444 = io_master_in_sync ? $signed(io_master_in_data) : $signed(_GEN_428); // @[Bus.scala 218:73:@230.14]
  assign _GEN_445 = io_master_in_sync ? io_master_in_trans_type : _GEN_429; // @[Bus.scala 218:73:@230.14]
  assign _GEN_446 = io_master_in_sync ? resp_signal_r_ack : _GEN_430; // @[Bus.scala 218:73:@230.14]
  assign _GEN_447 = io_master_in_sync ? $signed(resp_signal_r_data) : $signed(_GEN_431); // @[Bus.scala 218:73:@230.14]
  assign _GEN_448 = io_master_in_sync ? $signed(_T_245) : $signed(slave_out1_r_addr); // @[Bus.scala 218:73:@230.14]
  assign _GEN_449 = io_master_in_sync ? $signed(io_master_in_data) : $signed(slave_out1_r_data); // @[Bus.scala 218:73:@230.14]
  assign _GEN_450 = io_master_in_sync ? io_master_in_trans_type : slave_out1_r_trans_type; // @[Bus.scala 218:73:@230.14]
  assign _GEN_451 = io_master_in_sync ? 1'h0 : _GEN_432; // @[Bus.scala 218:73:@230.14]
  assign _GEN_452 = io_master_in_sync ? 1'h0 : _GEN_433; // @[Bus.scala 218:73:@230.14]
  assign _GEN_453 = io_master_in_sync ? 1'h0 : _GEN_434; // @[Bus.scala 218:73:@230.14]
  assign _GEN_454 = io_master_in_sync ? 1'h0 : _GEN_435; // @[Bus.scala 218:73:@230.14]
  assign _GEN_455 = io_master_in_sync ? 1'h0 : _GEN_436; // @[Bus.scala 218:73:@230.14]
  assign _GEN_456 = io_master_in_sync ? 1'h0 : _GEN_437; // @[Bus.scala 218:73:@230.14]
  assign _GEN_457 = io_master_in_sync ? 1'h0 : _GEN_438; // @[Bus.scala 218:73:@230.14]
  assign _GEN_458 = io_master_in_sync ? 1'h1 : _GEN_439; // @[Bus.scala 218:73:@230.14]
  assign _GEN_459 = io_master_in_sync ? 1'h0 : _GEN_440; // @[Bus.scala 218:73:@230.14]
  assign _GEN_460 = io_master_in_sync ? 1'h0 : _GEN_441; // @[Bus.scala 218:73:@230.14]
  assign _GEN_461 = _T_241 ? _GEN_442 : _GEN_424; // @[Bus.scala 217:81:@229.12]
  assign _GEN_462 = _T_241 ? $signed(_GEN_443) : $signed(_GEN_427); // @[Bus.scala 217:81:@229.12]
  assign _GEN_463 = _T_241 ? $signed(_GEN_444) : $signed(_GEN_428); // @[Bus.scala 217:81:@229.12]
  assign _GEN_464 = _T_241 ? _GEN_445 : _GEN_429; // @[Bus.scala 217:81:@229.12]
  assign _GEN_465 = _T_241 ? _GEN_446 : _GEN_430; // @[Bus.scala 217:81:@229.12]
  assign _GEN_466 = _T_241 ? $signed(_GEN_447) : $signed(_GEN_431); // @[Bus.scala 217:81:@229.12]
  assign _GEN_467 = _T_241 ? $signed(_GEN_448) : $signed(slave_out1_r_addr); // @[Bus.scala 217:81:@229.12]
  assign _GEN_468 = _T_241 ? $signed(_GEN_449) : $signed(slave_out1_r_data); // @[Bus.scala 217:81:@229.12]
  assign _GEN_469 = _T_241 ? _GEN_450 : slave_out1_r_trans_type; // @[Bus.scala 217:81:@229.12]
  assign _GEN_470 = _T_241 ? _GEN_451 : _GEN_432; // @[Bus.scala 217:81:@229.12]
  assign _GEN_471 = _T_241 ? _GEN_452 : _GEN_433; // @[Bus.scala 217:81:@229.12]
  assign _GEN_472 = _T_241 ? _GEN_453 : _GEN_434; // @[Bus.scala 217:81:@229.12]
  assign _GEN_473 = _T_241 ? _GEN_454 : _GEN_435; // @[Bus.scala 217:81:@229.12]
  assign _GEN_474 = _T_241 ? _GEN_455 : _GEN_436; // @[Bus.scala 217:81:@229.12]
  assign _GEN_475 = _T_241 ? _GEN_456 : _GEN_437; // @[Bus.scala 217:81:@229.12]
  assign _GEN_476 = _T_241 ? _GEN_457 : _GEN_438; // @[Bus.scala 217:81:@229.12]
  assign _GEN_477 = _T_241 ? _GEN_458 : _GEN_439; // @[Bus.scala 217:81:@229.12]
  assign _GEN_478 = _T_241 ? _GEN_459 : _GEN_440; // @[Bus.scala 217:81:@229.12]
  assign _GEN_479 = _T_241 ? _GEN_460 : _GEN_441; // @[Bus.scala 217:81:@229.12]
  assign _GEN_480 = _T_145 ? _GEN_461 : _GEN_424; // @[Bus.scala 216:72:@227.10]
  assign _GEN_481 = _T_145 ? $signed(_GEN_462) : $signed(_GEN_427); // @[Bus.scala 216:72:@227.10]
  assign _GEN_482 = _T_145 ? $signed(_GEN_463) : $signed(_GEN_428); // @[Bus.scala 216:72:@227.10]
  assign _GEN_483 = _T_145 ? _GEN_464 : _GEN_429; // @[Bus.scala 216:72:@227.10]
  assign _GEN_484 = _T_145 ? _GEN_465 : _GEN_430; // @[Bus.scala 216:72:@227.10]
  assign _GEN_485 = _T_145 ? $signed(_GEN_466) : $signed(_GEN_431); // @[Bus.scala 216:72:@227.10]
  assign _GEN_486 = _T_145 ? $signed(_GEN_467) : $signed(slave_out1_r_addr); // @[Bus.scala 216:72:@227.10]
  assign _GEN_487 = _T_145 ? $signed(_GEN_468) : $signed(slave_out1_r_data); // @[Bus.scala 216:72:@227.10]
  assign _GEN_488 = _T_145 ? _GEN_469 : slave_out1_r_trans_type; // @[Bus.scala 216:72:@227.10]
  assign _GEN_489 = _T_145 ? _GEN_470 : _GEN_432; // @[Bus.scala 216:72:@227.10]
  assign _GEN_490 = _T_145 ? _GEN_471 : _GEN_433; // @[Bus.scala 216:72:@227.10]
  assign _GEN_491 = _T_145 ? _GEN_472 : _GEN_434; // @[Bus.scala 216:72:@227.10]
  assign _GEN_492 = _T_145 ? _GEN_473 : _GEN_435; // @[Bus.scala 216:72:@227.10]
  assign _GEN_493 = _T_145 ? _GEN_474 : _GEN_436; // @[Bus.scala 216:72:@227.10]
  assign _GEN_494 = _T_145 ? _GEN_475 : _GEN_437; // @[Bus.scala 216:72:@227.10]
  assign _GEN_495 = _T_145 ? _GEN_476 : _GEN_438; // @[Bus.scala 216:72:@227.10]
  assign _GEN_496 = _T_145 ? _GEN_477 : _GEN_439; // @[Bus.scala 216:72:@227.10]
  assign _GEN_497 = _T_145 ? _GEN_478 : _GEN_440; // @[Bus.scala 216:72:@227.10]
  assign _GEN_498 = _T_145 ? _GEN_479 : _GEN_441; // @[Bus.scala 216:72:@227.10]
  assign _GEN_499 = _T_100 ? _GEN_480 : _GEN_424; // @[Bus.scala 215:74:@225.8]
  assign _GEN_500 = _T_100 ? $signed(_GEN_481) : $signed(_GEN_427); // @[Bus.scala 215:74:@225.8]
  assign _GEN_501 = _T_100 ? $signed(_GEN_482) : $signed(_GEN_428); // @[Bus.scala 215:74:@225.8]
  assign _GEN_502 = _T_100 ? _GEN_483 : _GEN_429; // @[Bus.scala 215:74:@225.8]
  assign _GEN_503 = _T_100 ? _GEN_484 : _GEN_430; // @[Bus.scala 215:74:@225.8]
  assign _GEN_504 = _T_100 ? $signed(_GEN_485) : $signed(_GEN_431); // @[Bus.scala 215:74:@225.8]
  assign _GEN_505 = _T_100 ? $signed(_GEN_486) : $signed(slave_out1_r_addr); // @[Bus.scala 215:74:@225.8]
  assign _GEN_506 = _T_100 ? $signed(_GEN_487) : $signed(slave_out1_r_data); // @[Bus.scala 215:74:@225.8]
  assign _GEN_507 = _T_100 ? _GEN_488 : slave_out1_r_trans_type; // @[Bus.scala 215:74:@225.8]
  assign _GEN_508 = _T_100 ? _GEN_489 : _GEN_432; // @[Bus.scala 215:74:@225.8]
  assign _GEN_509 = _T_100 ? _GEN_490 : _GEN_433; // @[Bus.scala 215:74:@225.8]
  assign _GEN_510 = _T_100 ? _GEN_491 : _GEN_434; // @[Bus.scala 215:74:@225.8]
  assign _GEN_511 = _T_100 ? _GEN_492 : _GEN_435; // @[Bus.scala 215:74:@225.8]
  assign _GEN_512 = _T_100 ? _GEN_493 : _GEN_436; // @[Bus.scala 215:74:@225.8]
  assign _GEN_513 = _T_100 ? _GEN_494 : _GEN_437; // @[Bus.scala 215:74:@225.8]
  assign _GEN_514 = _T_100 ? _GEN_495 : _GEN_438; // @[Bus.scala 215:74:@225.8]
  assign _GEN_515 = _T_100 ? _GEN_496 : _GEN_439; // @[Bus.scala 215:74:@225.8]
  assign _GEN_516 = _T_100 ? _GEN_497 : _GEN_440; // @[Bus.scala 215:74:@225.8]
  assign _GEN_517 = _T_100 ? _GEN_498 : _GEN_441; // @[Bus.scala 215:74:@225.8]
  assign _GEN_518 = _T_97 ? _GEN_499 : _GEN_424; // @[Bus.scala 214:41:@222.6]
  assign _GEN_519 = _T_97 ? $signed(_GEN_500) : $signed(_GEN_427); // @[Bus.scala 214:41:@222.6]
  assign _GEN_520 = _T_97 ? $signed(_GEN_501) : $signed(_GEN_428); // @[Bus.scala 214:41:@222.6]
  assign _GEN_521 = _T_97 ? _GEN_502 : _GEN_429; // @[Bus.scala 214:41:@222.6]
  assign _GEN_522 = _T_97 ? _GEN_503 : _GEN_430; // @[Bus.scala 214:41:@222.6]
  assign _GEN_523 = _T_97 ? $signed(_GEN_504) : $signed(_GEN_431); // @[Bus.scala 214:41:@222.6]
  assign _GEN_524 = _T_97 ? $signed(_GEN_505) : $signed(slave_out1_r_addr); // @[Bus.scala 214:41:@222.6]
  assign _GEN_525 = _T_97 ? $signed(_GEN_506) : $signed(slave_out1_r_data); // @[Bus.scala 214:41:@222.6]
  assign _GEN_526 = _T_97 ? _GEN_507 : slave_out1_r_trans_type; // @[Bus.scala 214:41:@222.6]
  assign _GEN_527 = _T_97 ? _GEN_508 : _GEN_432; // @[Bus.scala 214:41:@222.6]
  assign _GEN_528 = _T_97 ? _GEN_509 : _GEN_433; // @[Bus.scala 214:41:@222.6]
  assign _GEN_529 = _T_97 ? _GEN_510 : _GEN_434; // @[Bus.scala 214:41:@222.6]
  assign _GEN_530 = _T_97 ? _GEN_511 : _GEN_435; // @[Bus.scala 214:41:@222.6]
  assign _GEN_531 = _T_97 ? _GEN_512 : _GEN_436; // @[Bus.scala 214:41:@222.6]
  assign _GEN_532 = _T_97 ? _GEN_513 : _GEN_437; // @[Bus.scala 214:41:@222.6]
  assign _GEN_533 = _T_97 ? _GEN_514 : _GEN_438; // @[Bus.scala 214:41:@222.6]
  assign _GEN_534 = _T_97 ? _GEN_515 : _GEN_439; // @[Bus.scala 214:41:@222.6]
  assign _GEN_535 = _T_97 ? _GEN_516 : _GEN_440; // @[Bus.scala 214:41:@222.6]
  assign _GEN_536 = _T_97 ? _GEN_517 : _GEN_441; // @[Bus.scala 214:41:@222.6]
  assign _GEN_537 = io_master_in_sync ? 4'h4 : _GEN_518; // @[Bus.scala 247:73:@269.14]
  assign _GEN_538 = io_master_in_sync ? $signed(_T_245) : $signed(_GEN_519); // @[Bus.scala 247:73:@269.14]
  assign _GEN_539 = io_master_in_sync ? $signed(32'sh0) : $signed(_GEN_520); // @[Bus.scala 247:73:@269.14]
  assign _GEN_540 = io_master_in_sync ? io_master_in_trans_type : _GEN_521; // @[Bus.scala 247:73:@269.14]
  assign _GEN_541 = io_master_in_sync ? resp_signal_r_ack : _GEN_522; // @[Bus.scala 247:73:@269.14]
  assign _GEN_542 = io_master_in_sync ? $signed(resp_signal_r_data) : $signed(_GEN_523); // @[Bus.scala 247:73:@269.14]
  assign _GEN_543 = io_master_in_sync ? $signed(_T_245) : $signed(_GEN_524); // @[Bus.scala 247:73:@269.14]
  assign _GEN_544 = io_master_in_sync ? $signed(32'sh0) : $signed(_GEN_525); // @[Bus.scala 247:73:@269.14]
  assign _GEN_545 = io_master_in_sync ? io_master_in_trans_type : _GEN_526; // @[Bus.scala 247:73:@269.14]
  assign _GEN_546 = io_master_in_sync ? 1'h0 : _GEN_527; // @[Bus.scala 247:73:@269.14]
  assign _GEN_547 = io_master_in_sync ? 1'h0 : _GEN_528; // @[Bus.scala 247:73:@269.14]
  assign _GEN_548 = io_master_in_sync ? 1'h0 : _GEN_529; // @[Bus.scala 247:73:@269.14]
  assign _GEN_549 = io_master_in_sync ? 1'h0 : _GEN_530; // @[Bus.scala 247:73:@269.14]
  assign _GEN_550 = io_master_in_sync ? 1'h0 : _GEN_531; // @[Bus.scala 247:73:@269.14]
  assign _GEN_551 = io_master_in_sync ? 1'h0 : _GEN_532; // @[Bus.scala 247:73:@269.14]
  assign _GEN_552 = io_master_in_sync ? 1'h0 : _GEN_533; // @[Bus.scala 247:73:@269.14]
  assign _GEN_553 = io_master_in_sync ? 1'h1 : _GEN_534; // @[Bus.scala 247:73:@269.14]
  assign _GEN_554 = io_master_in_sync ? 1'h0 : _GEN_535; // @[Bus.scala 247:73:@269.14]
  assign _GEN_555 = io_master_in_sync ? 1'h0 : _GEN_536; // @[Bus.scala 247:73:@269.14]
  assign _GEN_556 = _T_241 ? _GEN_537 : _GEN_518; // @[Bus.scala 246:81:@268.12]
  assign _GEN_557 = _T_241 ? $signed(_GEN_538) : $signed(_GEN_519); // @[Bus.scala 246:81:@268.12]
  assign _GEN_558 = _T_241 ? $signed(_GEN_539) : $signed(_GEN_520); // @[Bus.scala 246:81:@268.12]
  assign _GEN_559 = _T_241 ? _GEN_540 : _GEN_521; // @[Bus.scala 246:81:@268.12]
  assign _GEN_560 = _T_241 ? _GEN_541 : _GEN_522; // @[Bus.scala 246:81:@268.12]
  assign _GEN_561 = _T_241 ? $signed(_GEN_542) : $signed(_GEN_523); // @[Bus.scala 246:81:@268.12]
  assign _GEN_562 = _T_241 ? $signed(_GEN_543) : $signed(_GEN_524); // @[Bus.scala 246:81:@268.12]
  assign _GEN_563 = _T_241 ? $signed(_GEN_544) : $signed(_GEN_525); // @[Bus.scala 246:81:@268.12]
  assign _GEN_564 = _T_241 ? _GEN_545 : _GEN_526; // @[Bus.scala 246:81:@268.12]
  assign _GEN_565 = _T_241 ? _GEN_546 : _GEN_527; // @[Bus.scala 246:81:@268.12]
  assign _GEN_566 = _T_241 ? _GEN_547 : _GEN_528; // @[Bus.scala 246:81:@268.12]
  assign _GEN_567 = _T_241 ? _GEN_548 : _GEN_529; // @[Bus.scala 246:81:@268.12]
  assign _GEN_568 = _T_241 ? _GEN_549 : _GEN_530; // @[Bus.scala 246:81:@268.12]
  assign _GEN_569 = _T_241 ? _GEN_550 : _GEN_531; // @[Bus.scala 246:81:@268.12]
  assign _GEN_570 = _T_241 ? _GEN_551 : _GEN_532; // @[Bus.scala 246:81:@268.12]
  assign _GEN_571 = _T_241 ? _GEN_552 : _GEN_533; // @[Bus.scala 246:81:@268.12]
  assign _GEN_572 = _T_241 ? _GEN_553 : _GEN_534; // @[Bus.scala 246:81:@268.12]
  assign _GEN_573 = _T_241 ? _GEN_554 : _GEN_535; // @[Bus.scala 246:81:@268.12]
  assign _GEN_574 = _T_241 ? _GEN_555 : _GEN_536; // @[Bus.scala 246:81:@268.12]
  assign _GEN_575 = _T_145 ? _GEN_556 : _GEN_518; // @[Bus.scala 245:72:@266.10]
  assign _GEN_576 = _T_145 ? $signed(_GEN_557) : $signed(_GEN_519); // @[Bus.scala 245:72:@266.10]
  assign _GEN_577 = _T_145 ? $signed(_GEN_558) : $signed(_GEN_520); // @[Bus.scala 245:72:@266.10]
  assign _GEN_578 = _T_145 ? _GEN_559 : _GEN_521; // @[Bus.scala 245:72:@266.10]
  assign _GEN_579 = _T_145 ? _GEN_560 : _GEN_522; // @[Bus.scala 245:72:@266.10]
  assign _GEN_580 = _T_145 ? $signed(_GEN_561) : $signed(_GEN_523); // @[Bus.scala 245:72:@266.10]
  assign _GEN_581 = _T_145 ? $signed(_GEN_562) : $signed(_GEN_524); // @[Bus.scala 245:72:@266.10]
  assign _GEN_582 = _T_145 ? $signed(_GEN_563) : $signed(_GEN_525); // @[Bus.scala 245:72:@266.10]
  assign _GEN_583 = _T_145 ? _GEN_564 : _GEN_526; // @[Bus.scala 245:72:@266.10]
  assign _GEN_584 = _T_145 ? _GEN_565 : _GEN_527; // @[Bus.scala 245:72:@266.10]
  assign _GEN_585 = _T_145 ? _GEN_566 : _GEN_528; // @[Bus.scala 245:72:@266.10]
  assign _GEN_586 = _T_145 ? _GEN_567 : _GEN_529; // @[Bus.scala 245:72:@266.10]
  assign _GEN_587 = _T_145 ? _GEN_568 : _GEN_530; // @[Bus.scala 245:72:@266.10]
  assign _GEN_588 = _T_145 ? _GEN_569 : _GEN_531; // @[Bus.scala 245:72:@266.10]
  assign _GEN_589 = _T_145 ? _GEN_570 : _GEN_532; // @[Bus.scala 245:72:@266.10]
  assign _GEN_590 = _T_145 ? _GEN_571 : _GEN_533; // @[Bus.scala 245:72:@266.10]
  assign _GEN_591 = _T_145 ? _GEN_572 : _GEN_534; // @[Bus.scala 245:72:@266.10]
  assign _GEN_592 = _T_145 ? _GEN_573 : _GEN_535; // @[Bus.scala 245:72:@266.10]
  assign _GEN_593 = _T_145 ? _GEN_574 : _GEN_536; // @[Bus.scala 245:72:@266.10]
  assign _GEN_594 = _T_98 ? _GEN_575 : _GEN_518; // @[Bus.scala 244:73:@264.8]
  assign _GEN_595 = _T_98 ? $signed(_GEN_576) : $signed(_GEN_519); // @[Bus.scala 244:73:@264.8]
  assign _GEN_596 = _T_98 ? $signed(_GEN_577) : $signed(_GEN_520); // @[Bus.scala 244:73:@264.8]
  assign _GEN_597 = _T_98 ? _GEN_578 : _GEN_521; // @[Bus.scala 244:73:@264.8]
  assign _GEN_598 = _T_98 ? _GEN_579 : _GEN_522; // @[Bus.scala 244:73:@264.8]
  assign _GEN_599 = _T_98 ? $signed(_GEN_580) : $signed(_GEN_523); // @[Bus.scala 244:73:@264.8]
  assign _GEN_600 = _T_98 ? $signed(_GEN_581) : $signed(_GEN_524); // @[Bus.scala 244:73:@264.8]
  assign _GEN_601 = _T_98 ? $signed(_GEN_582) : $signed(_GEN_525); // @[Bus.scala 244:73:@264.8]
  assign _GEN_602 = _T_98 ? _GEN_583 : _GEN_526; // @[Bus.scala 244:73:@264.8]
  assign _GEN_603 = _T_98 ? _GEN_584 : _GEN_527; // @[Bus.scala 244:73:@264.8]
  assign _GEN_604 = _T_98 ? _GEN_585 : _GEN_528; // @[Bus.scala 244:73:@264.8]
  assign _GEN_605 = _T_98 ? _GEN_586 : _GEN_529; // @[Bus.scala 244:73:@264.8]
  assign _GEN_606 = _T_98 ? _GEN_587 : _GEN_530; // @[Bus.scala 244:73:@264.8]
  assign _GEN_607 = _T_98 ? _GEN_588 : _GEN_531; // @[Bus.scala 244:73:@264.8]
  assign _GEN_608 = _T_98 ? _GEN_589 : _GEN_532; // @[Bus.scala 244:73:@264.8]
  assign _GEN_609 = _T_98 ? _GEN_590 : _GEN_533; // @[Bus.scala 244:73:@264.8]
  assign _GEN_610 = _T_98 ? _GEN_591 : _GEN_534; // @[Bus.scala 244:73:@264.8]
  assign _GEN_611 = _T_98 ? _GEN_592 : _GEN_535; // @[Bus.scala 244:73:@264.8]
  assign _GEN_612 = _T_98 ? _GEN_593 : _GEN_536; // @[Bus.scala 244:73:@264.8]
  assign _GEN_613 = _T_97 ? _GEN_594 : _GEN_518; // @[Bus.scala 243:41:@262.6]
  assign _GEN_614 = _T_97 ? $signed(_GEN_595) : $signed(_GEN_519); // @[Bus.scala 243:41:@262.6]
  assign _GEN_615 = _T_97 ? $signed(_GEN_596) : $signed(_GEN_520); // @[Bus.scala 243:41:@262.6]
  assign _GEN_616 = _T_97 ? _GEN_597 : _GEN_521; // @[Bus.scala 243:41:@262.6]
  assign _GEN_617 = _T_97 ? _GEN_598 : _GEN_522; // @[Bus.scala 243:41:@262.6]
  assign _GEN_618 = _T_97 ? $signed(_GEN_599) : $signed(_GEN_523); // @[Bus.scala 243:41:@262.6]
  assign _GEN_619 = _T_97 ? $signed(_GEN_600) : $signed(_GEN_524); // @[Bus.scala 243:41:@262.6]
  assign _GEN_620 = _T_97 ? $signed(_GEN_601) : $signed(_GEN_525); // @[Bus.scala 243:41:@262.6]
  assign _GEN_621 = _T_97 ? _GEN_602 : _GEN_526; // @[Bus.scala 243:41:@262.6]
  assign _GEN_622 = _T_97 ? _GEN_603 : _GEN_527; // @[Bus.scala 243:41:@262.6]
  assign _GEN_623 = _T_97 ? _GEN_604 : _GEN_528; // @[Bus.scala 243:41:@262.6]
  assign _GEN_624 = _T_97 ? _GEN_605 : _GEN_529; // @[Bus.scala 243:41:@262.6]
  assign _GEN_625 = _T_97 ? _GEN_606 : _GEN_530; // @[Bus.scala 243:41:@262.6]
  assign _GEN_626 = _T_97 ? _GEN_607 : _GEN_531; // @[Bus.scala 243:41:@262.6]
  assign _GEN_627 = _T_97 ? _GEN_608 : _GEN_532; // @[Bus.scala 243:41:@262.6]
  assign _GEN_628 = _T_97 ? _GEN_609 : _GEN_533; // @[Bus.scala 243:41:@262.6]
  assign _GEN_629 = _T_97 ? _GEN_610 : _GEN_534; // @[Bus.scala 243:41:@262.6]
  assign _GEN_630 = _T_97 ? _GEN_611 : _GEN_535; // @[Bus.scala 243:41:@262.6]
  assign _GEN_631 = _T_97 ? _GEN_612 : _GEN_536; // @[Bus.scala 243:41:@262.6]
  assign _T_293 = $signed(io_master_in_addr) <= $signed(32'sh17); // @[Bus.scala 275:65:@307.12]
  assign _T_295 = $signed(-32'sh10) + $signed(io_master_in_addr); // @[Bus.scala 278:93:@311.16]
  assign _T_296 = $signed(-32'sh10) + $signed(io_master_in_addr); // @[Bus.scala 278:93:@312.16]
  assign _T_297 = $signed(_T_296); // @[Bus.scala 278:93:@313.16]
  assign _GEN_632 = io_master_in_sync ? 4'h6 : _GEN_613; // @[Bus.scala 276:73:@309.14]
  assign _GEN_633 = io_master_in_sync ? $signed(_T_297) : $signed(_GEN_614); // @[Bus.scala 276:73:@309.14]
  assign _GEN_634 = io_master_in_sync ? $signed(io_master_in_data) : $signed(_GEN_615); // @[Bus.scala 276:73:@309.14]
  assign _GEN_635 = io_master_in_sync ? io_master_in_trans_type : _GEN_616; // @[Bus.scala 276:73:@309.14]
  assign _GEN_636 = io_master_in_sync ? resp_signal_r_ack : _GEN_617; // @[Bus.scala 276:73:@309.14]
  assign _GEN_637 = io_master_in_sync ? $signed(resp_signal_r_data) : $signed(_GEN_618); // @[Bus.scala 276:73:@309.14]
  assign _GEN_638 = io_master_in_sync ? $signed(_T_297) : $signed(slave_out2_r_addr); // @[Bus.scala 276:73:@309.14]
  assign _GEN_639 = io_master_in_sync ? $signed(io_master_in_data) : $signed(slave_out2_r_data); // @[Bus.scala 276:73:@309.14]
  assign _GEN_640 = io_master_in_sync ? io_master_in_trans_type : slave_out2_r_trans_type; // @[Bus.scala 276:73:@309.14]
  assign _GEN_641 = io_master_in_sync ? 1'h0 : _GEN_622; // @[Bus.scala 276:73:@309.14]
  assign _GEN_642 = io_master_in_sync ? 1'h0 : _GEN_623; // @[Bus.scala 276:73:@309.14]
  assign _GEN_643 = io_master_in_sync ? 1'h0 : _GEN_624; // @[Bus.scala 276:73:@309.14]
  assign _GEN_644 = io_master_in_sync ? 1'h0 : _GEN_625; // @[Bus.scala 276:73:@309.14]
  assign _GEN_645 = io_master_in_sync ? 1'h0 : _GEN_626; // @[Bus.scala 276:73:@309.14]
  assign _GEN_646 = io_master_in_sync ? 1'h0 : _GEN_627; // @[Bus.scala 276:73:@309.14]
  assign _GEN_647 = io_master_in_sync ? 1'h0 : _GEN_628; // @[Bus.scala 276:73:@309.14]
  assign _GEN_648 = io_master_in_sync ? 1'h0 : _GEN_629; // @[Bus.scala 276:73:@309.14]
  assign _GEN_649 = io_master_in_sync ? 1'h1 : _GEN_630; // @[Bus.scala 276:73:@309.14]
  assign _GEN_650 = io_master_in_sync ? 1'h0 : _GEN_631; // @[Bus.scala 276:73:@309.14]
  assign _GEN_651 = _T_293 ? _GEN_632 : _GEN_613; // @[Bus.scala 275:81:@308.12]
  assign _GEN_652 = _T_293 ? $signed(_GEN_633) : $signed(_GEN_614); // @[Bus.scala 275:81:@308.12]
  assign _GEN_653 = _T_293 ? $signed(_GEN_634) : $signed(_GEN_615); // @[Bus.scala 275:81:@308.12]
  assign _GEN_654 = _T_293 ? _GEN_635 : _GEN_616; // @[Bus.scala 275:81:@308.12]
  assign _GEN_655 = _T_293 ? _GEN_636 : _GEN_617; // @[Bus.scala 275:81:@308.12]
  assign _GEN_656 = _T_293 ? $signed(_GEN_637) : $signed(_GEN_618); // @[Bus.scala 275:81:@308.12]
  assign _GEN_657 = _T_293 ? $signed(_GEN_638) : $signed(slave_out2_r_addr); // @[Bus.scala 275:81:@308.12]
  assign _GEN_658 = _T_293 ? $signed(_GEN_639) : $signed(slave_out2_r_data); // @[Bus.scala 275:81:@308.12]
  assign _GEN_659 = _T_293 ? _GEN_640 : slave_out2_r_trans_type; // @[Bus.scala 275:81:@308.12]
  assign _GEN_660 = _T_293 ? _GEN_641 : _GEN_622; // @[Bus.scala 275:81:@308.12]
  assign _GEN_661 = _T_293 ? _GEN_642 : _GEN_623; // @[Bus.scala 275:81:@308.12]
  assign _GEN_662 = _T_293 ? _GEN_643 : _GEN_624; // @[Bus.scala 275:81:@308.12]
  assign _GEN_663 = _T_293 ? _GEN_644 : _GEN_625; // @[Bus.scala 275:81:@308.12]
  assign _GEN_664 = _T_293 ? _GEN_645 : _GEN_626; // @[Bus.scala 275:81:@308.12]
  assign _GEN_665 = _T_293 ? _GEN_646 : _GEN_627; // @[Bus.scala 275:81:@308.12]
  assign _GEN_666 = _T_293 ? _GEN_647 : _GEN_628; // @[Bus.scala 275:81:@308.12]
  assign _GEN_667 = _T_293 ? _GEN_648 : _GEN_629; // @[Bus.scala 275:81:@308.12]
  assign _GEN_668 = _T_293 ? _GEN_649 : _GEN_630; // @[Bus.scala 275:81:@308.12]
  assign _GEN_669 = _T_293 ? _GEN_650 : _GEN_631; // @[Bus.scala 275:81:@308.12]
  assign _GEN_670 = _T_154 ? _GEN_651 : _GEN_613; // @[Bus.scala 274:73:@306.10]
  assign _GEN_671 = _T_154 ? $signed(_GEN_652) : $signed(_GEN_614); // @[Bus.scala 274:73:@306.10]
  assign _GEN_672 = _T_154 ? $signed(_GEN_653) : $signed(_GEN_615); // @[Bus.scala 274:73:@306.10]
  assign _GEN_673 = _T_154 ? _GEN_654 : _GEN_616; // @[Bus.scala 274:73:@306.10]
  assign _GEN_674 = _T_154 ? _GEN_655 : _GEN_617; // @[Bus.scala 274:73:@306.10]
  assign _GEN_675 = _T_154 ? $signed(_GEN_656) : $signed(_GEN_618); // @[Bus.scala 274:73:@306.10]
  assign _GEN_676 = _T_154 ? $signed(_GEN_657) : $signed(slave_out2_r_addr); // @[Bus.scala 274:73:@306.10]
  assign _GEN_677 = _T_154 ? $signed(_GEN_658) : $signed(slave_out2_r_data); // @[Bus.scala 274:73:@306.10]
  assign _GEN_678 = _T_154 ? _GEN_659 : slave_out2_r_trans_type; // @[Bus.scala 274:73:@306.10]
  assign _GEN_679 = _T_154 ? _GEN_660 : _GEN_622; // @[Bus.scala 274:73:@306.10]
  assign _GEN_680 = _T_154 ? _GEN_661 : _GEN_623; // @[Bus.scala 274:73:@306.10]
  assign _GEN_681 = _T_154 ? _GEN_662 : _GEN_624; // @[Bus.scala 274:73:@306.10]
  assign _GEN_682 = _T_154 ? _GEN_663 : _GEN_625; // @[Bus.scala 274:73:@306.10]
  assign _GEN_683 = _T_154 ? _GEN_664 : _GEN_626; // @[Bus.scala 274:73:@306.10]
  assign _GEN_684 = _T_154 ? _GEN_665 : _GEN_627; // @[Bus.scala 274:73:@306.10]
  assign _GEN_685 = _T_154 ? _GEN_666 : _GEN_628; // @[Bus.scala 274:73:@306.10]
  assign _GEN_686 = _T_154 ? _GEN_667 : _GEN_629; // @[Bus.scala 274:73:@306.10]
  assign _GEN_687 = _T_154 ? _GEN_668 : _GEN_630; // @[Bus.scala 274:73:@306.10]
  assign _GEN_688 = _T_154 ? _GEN_669 : _GEN_631; // @[Bus.scala 274:73:@306.10]
  assign _GEN_689 = _T_100 ? _GEN_670 : _GEN_613; // @[Bus.scala 273:74:@304.8]
  assign _GEN_690 = _T_100 ? $signed(_GEN_671) : $signed(_GEN_614); // @[Bus.scala 273:74:@304.8]
  assign _GEN_691 = _T_100 ? $signed(_GEN_672) : $signed(_GEN_615); // @[Bus.scala 273:74:@304.8]
  assign _GEN_692 = _T_100 ? _GEN_673 : _GEN_616; // @[Bus.scala 273:74:@304.8]
  assign _GEN_693 = _T_100 ? _GEN_674 : _GEN_617; // @[Bus.scala 273:74:@304.8]
  assign _GEN_694 = _T_100 ? $signed(_GEN_675) : $signed(_GEN_618); // @[Bus.scala 273:74:@304.8]
  assign _GEN_695 = _T_100 ? $signed(_GEN_676) : $signed(slave_out2_r_addr); // @[Bus.scala 273:74:@304.8]
  assign _GEN_696 = _T_100 ? $signed(_GEN_677) : $signed(slave_out2_r_data); // @[Bus.scala 273:74:@304.8]
  assign _GEN_697 = _T_100 ? _GEN_678 : slave_out2_r_trans_type; // @[Bus.scala 273:74:@304.8]
  assign _GEN_698 = _T_100 ? _GEN_679 : _GEN_622; // @[Bus.scala 273:74:@304.8]
  assign _GEN_699 = _T_100 ? _GEN_680 : _GEN_623; // @[Bus.scala 273:74:@304.8]
  assign _GEN_700 = _T_100 ? _GEN_681 : _GEN_624; // @[Bus.scala 273:74:@304.8]
  assign _GEN_701 = _T_100 ? _GEN_682 : _GEN_625; // @[Bus.scala 273:74:@304.8]
  assign _GEN_702 = _T_100 ? _GEN_683 : _GEN_626; // @[Bus.scala 273:74:@304.8]
  assign _GEN_703 = _T_100 ? _GEN_684 : _GEN_627; // @[Bus.scala 273:74:@304.8]
  assign _GEN_704 = _T_100 ? _GEN_685 : _GEN_628; // @[Bus.scala 273:74:@304.8]
  assign _GEN_705 = _T_100 ? _GEN_686 : _GEN_629; // @[Bus.scala 273:74:@304.8]
  assign _GEN_706 = _T_100 ? _GEN_687 : _GEN_630; // @[Bus.scala 273:74:@304.8]
  assign _GEN_707 = _T_100 ? _GEN_688 : _GEN_631; // @[Bus.scala 273:74:@304.8]
  assign _GEN_708 = _T_97 ? _GEN_689 : _GEN_613; // @[Bus.scala 272:41:@301.6]
  assign _GEN_709 = _T_97 ? $signed(_GEN_690) : $signed(_GEN_614); // @[Bus.scala 272:41:@301.6]
  assign _GEN_710 = _T_97 ? $signed(_GEN_691) : $signed(_GEN_615); // @[Bus.scala 272:41:@301.6]
  assign _GEN_711 = _T_97 ? _GEN_692 : _GEN_616; // @[Bus.scala 272:41:@301.6]
  assign _GEN_712 = _T_97 ? _GEN_693 : _GEN_617; // @[Bus.scala 272:41:@301.6]
  assign _GEN_713 = _T_97 ? $signed(_GEN_694) : $signed(_GEN_618); // @[Bus.scala 272:41:@301.6]
  assign _GEN_714 = _T_97 ? $signed(_GEN_695) : $signed(slave_out2_r_addr); // @[Bus.scala 272:41:@301.6]
  assign _GEN_715 = _T_97 ? $signed(_GEN_696) : $signed(slave_out2_r_data); // @[Bus.scala 272:41:@301.6]
  assign _GEN_716 = _T_97 ? _GEN_697 : slave_out2_r_trans_type; // @[Bus.scala 272:41:@301.6]
  assign _GEN_717 = _T_97 ? _GEN_698 : _GEN_622; // @[Bus.scala 272:41:@301.6]
  assign _GEN_718 = _T_97 ? _GEN_699 : _GEN_623; // @[Bus.scala 272:41:@301.6]
  assign _GEN_719 = _T_97 ? _GEN_700 : _GEN_624; // @[Bus.scala 272:41:@301.6]
  assign _GEN_720 = _T_97 ? _GEN_701 : _GEN_625; // @[Bus.scala 272:41:@301.6]
  assign _GEN_721 = _T_97 ? _GEN_702 : _GEN_626; // @[Bus.scala 272:41:@301.6]
  assign _GEN_722 = _T_97 ? _GEN_703 : _GEN_627; // @[Bus.scala 272:41:@301.6]
  assign _GEN_723 = _T_97 ? _GEN_704 : _GEN_628; // @[Bus.scala 272:41:@301.6]
  assign _GEN_724 = _T_97 ? _GEN_705 : _GEN_629; // @[Bus.scala 272:41:@301.6]
  assign _GEN_725 = _T_97 ? _GEN_706 : _GEN_630; // @[Bus.scala 272:41:@301.6]
  assign _GEN_726 = _T_97 ? _GEN_707 : _GEN_631; // @[Bus.scala 272:41:@301.6]
  assign _GEN_727 = io_master_in_sync ? 4'h6 : _GEN_708; // @[Bus.scala 305:73:@348.14]
  assign _GEN_728 = io_master_in_sync ? $signed(_T_297) : $signed(_GEN_709); // @[Bus.scala 305:73:@348.14]
  assign _GEN_729 = io_master_in_sync ? $signed(32'sh0) : $signed(_GEN_710); // @[Bus.scala 305:73:@348.14]
  assign _GEN_730 = io_master_in_sync ? io_master_in_trans_type : _GEN_711; // @[Bus.scala 305:73:@348.14]
  assign _GEN_731 = io_master_in_sync ? resp_signal_r_ack : _GEN_712; // @[Bus.scala 305:73:@348.14]
  assign _GEN_732 = io_master_in_sync ? $signed(resp_signal_r_data) : $signed(_GEN_713); // @[Bus.scala 305:73:@348.14]
  assign _GEN_733 = io_master_in_sync ? $signed(_T_297) : $signed(_GEN_714); // @[Bus.scala 305:73:@348.14]
  assign _GEN_734 = io_master_in_sync ? $signed(32'sh0) : $signed(_GEN_715); // @[Bus.scala 305:73:@348.14]
  assign _GEN_735 = io_master_in_sync ? io_master_in_trans_type : _GEN_716; // @[Bus.scala 305:73:@348.14]
  assign _GEN_736 = io_master_in_sync ? 1'h0 : _GEN_717; // @[Bus.scala 305:73:@348.14]
  assign _GEN_737 = io_master_in_sync ? 1'h0 : _GEN_718; // @[Bus.scala 305:73:@348.14]
  assign _GEN_738 = io_master_in_sync ? 1'h0 : _GEN_719; // @[Bus.scala 305:73:@348.14]
  assign _GEN_739 = io_master_in_sync ? 1'h0 : _GEN_720; // @[Bus.scala 305:73:@348.14]
  assign _GEN_740 = io_master_in_sync ? 1'h0 : _GEN_721; // @[Bus.scala 305:73:@348.14]
  assign _GEN_741 = io_master_in_sync ? 1'h0 : _GEN_722; // @[Bus.scala 305:73:@348.14]
  assign _GEN_742 = io_master_in_sync ? 1'h0 : _GEN_723; // @[Bus.scala 305:73:@348.14]
  assign _GEN_743 = io_master_in_sync ? 1'h0 : _GEN_724; // @[Bus.scala 305:73:@348.14]
  assign _GEN_744 = io_master_in_sync ? 1'h1 : _GEN_725; // @[Bus.scala 305:73:@348.14]
  assign _GEN_745 = io_master_in_sync ? 1'h0 : _GEN_726; // @[Bus.scala 305:73:@348.14]
  assign _GEN_746 = _T_293 ? _GEN_727 : _GEN_708; // @[Bus.scala 304:81:@347.12]
  assign _GEN_747 = _T_293 ? $signed(_GEN_728) : $signed(_GEN_709); // @[Bus.scala 304:81:@347.12]
  assign _GEN_748 = _T_293 ? $signed(_GEN_729) : $signed(_GEN_710); // @[Bus.scala 304:81:@347.12]
  assign _GEN_749 = _T_293 ? _GEN_730 : _GEN_711; // @[Bus.scala 304:81:@347.12]
  assign _GEN_750 = _T_293 ? _GEN_731 : _GEN_712; // @[Bus.scala 304:81:@347.12]
  assign _GEN_751 = _T_293 ? $signed(_GEN_732) : $signed(_GEN_713); // @[Bus.scala 304:81:@347.12]
  assign _GEN_752 = _T_293 ? $signed(_GEN_733) : $signed(_GEN_714); // @[Bus.scala 304:81:@347.12]
  assign _GEN_753 = _T_293 ? $signed(_GEN_734) : $signed(_GEN_715); // @[Bus.scala 304:81:@347.12]
  assign _GEN_754 = _T_293 ? _GEN_735 : _GEN_716; // @[Bus.scala 304:81:@347.12]
  assign _GEN_755 = _T_293 ? _GEN_736 : _GEN_717; // @[Bus.scala 304:81:@347.12]
  assign _GEN_756 = _T_293 ? _GEN_737 : _GEN_718; // @[Bus.scala 304:81:@347.12]
  assign _GEN_757 = _T_293 ? _GEN_738 : _GEN_719; // @[Bus.scala 304:81:@347.12]
  assign _GEN_758 = _T_293 ? _GEN_739 : _GEN_720; // @[Bus.scala 304:81:@347.12]
  assign _GEN_759 = _T_293 ? _GEN_740 : _GEN_721; // @[Bus.scala 304:81:@347.12]
  assign _GEN_760 = _T_293 ? _GEN_741 : _GEN_722; // @[Bus.scala 304:81:@347.12]
  assign _GEN_761 = _T_293 ? _GEN_742 : _GEN_723; // @[Bus.scala 304:81:@347.12]
  assign _GEN_762 = _T_293 ? _GEN_743 : _GEN_724; // @[Bus.scala 304:81:@347.12]
  assign _GEN_763 = _T_293 ? _GEN_744 : _GEN_725; // @[Bus.scala 304:81:@347.12]
  assign _GEN_764 = _T_293 ? _GEN_745 : _GEN_726; // @[Bus.scala 304:81:@347.12]
  assign _GEN_765 = _T_154 ? _GEN_746 : _GEN_708; // @[Bus.scala 303:73:@345.10]
  assign _GEN_766 = _T_154 ? $signed(_GEN_747) : $signed(_GEN_709); // @[Bus.scala 303:73:@345.10]
  assign _GEN_767 = _T_154 ? $signed(_GEN_748) : $signed(_GEN_710); // @[Bus.scala 303:73:@345.10]
  assign _GEN_768 = _T_154 ? _GEN_749 : _GEN_711; // @[Bus.scala 303:73:@345.10]
  assign _GEN_769 = _T_154 ? _GEN_750 : _GEN_712; // @[Bus.scala 303:73:@345.10]
  assign _GEN_770 = _T_154 ? $signed(_GEN_751) : $signed(_GEN_713); // @[Bus.scala 303:73:@345.10]
  assign _GEN_771 = _T_154 ? $signed(_GEN_752) : $signed(_GEN_714); // @[Bus.scala 303:73:@345.10]
  assign _GEN_772 = _T_154 ? $signed(_GEN_753) : $signed(_GEN_715); // @[Bus.scala 303:73:@345.10]
  assign _GEN_773 = _T_154 ? _GEN_754 : _GEN_716; // @[Bus.scala 303:73:@345.10]
  assign _GEN_774 = _T_154 ? _GEN_755 : _GEN_717; // @[Bus.scala 303:73:@345.10]
  assign _GEN_775 = _T_154 ? _GEN_756 : _GEN_718; // @[Bus.scala 303:73:@345.10]
  assign _GEN_776 = _T_154 ? _GEN_757 : _GEN_719; // @[Bus.scala 303:73:@345.10]
  assign _GEN_777 = _T_154 ? _GEN_758 : _GEN_720; // @[Bus.scala 303:73:@345.10]
  assign _GEN_778 = _T_154 ? _GEN_759 : _GEN_721; // @[Bus.scala 303:73:@345.10]
  assign _GEN_779 = _T_154 ? _GEN_760 : _GEN_722; // @[Bus.scala 303:73:@345.10]
  assign _GEN_780 = _T_154 ? _GEN_761 : _GEN_723; // @[Bus.scala 303:73:@345.10]
  assign _GEN_781 = _T_154 ? _GEN_762 : _GEN_724; // @[Bus.scala 303:73:@345.10]
  assign _GEN_782 = _T_154 ? _GEN_763 : _GEN_725; // @[Bus.scala 303:73:@345.10]
  assign _GEN_783 = _T_154 ? _GEN_764 : _GEN_726; // @[Bus.scala 303:73:@345.10]
  assign _GEN_784 = _T_98 ? _GEN_765 : _GEN_708; // @[Bus.scala 302:73:@343.8]
  assign _GEN_785 = _T_98 ? $signed(_GEN_766) : $signed(_GEN_709); // @[Bus.scala 302:73:@343.8]
  assign _GEN_786 = _T_98 ? $signed(_GEN_767) : $signed(_GEN_710); // @[Bus.scala 302:73:@343.8]
  assign _GEN_787 = _T_98 ? _GEN_768 : _GEN_711; // @[Bus.scala 302:73:@343.8]
  assign _GEN_788 = _T_98 ? _GEN_769 : _GEN_712; // @[Bus.scala 302:73:@343.8]
  assign _GEN_789 = _T_98 ? $signed(_GEN_770) : $signed(_GEN_713); // @[Bus.scala 302:73:@343.8]
  assign _GEN_790 = _T_98 ? $signed(_GEN_771) : $signed(_GEN_714); // @[Bus.scala 302:73:@343.8]
  assign _GEN_791 = _T_98 ? $signed(_GEN_772) : $signed(_GEN_715); // @[Bus.scala 302:73:@343.8]
  assign _GEN_792 = _T_98 ? _GEN_773 : _GEN_716; // @[Bus.scala 302:73:@343.8]
  assign _GEN_793 = _T_98 ? _GEN_774 : _GEN_717; // @[Bus.scala 302:73:@343.8]
  assign _GEN_794 = _T_98 ? _GEN_775 : _GEN_718; // @[Bus.scala 302:73:@343.8]
  assign _GEN_795 = _T_98 ? _GEN_776 : _GEN_719; // @[Bus.scala 302:73:@343.8]
  assign _GEN_796 = _T_98 ? _GEN_777 : _GEN_720; // @[Bus.scala 302:73:@343.8]
  assign _GEN_797 = _T_98 ? _GEN_778 : _GEN_721; // @[Bus.scala 302:73:@343.8]
  assign _GEN_798 = _T_98 ? _GEN_779 : _GEN_722; // @[Bus.scala 302:73:@343.8]
  assign _GEN_799 = _T_98 ? _GEN_780 : _GEN_723; // @[Bus.scala 302:73:@343.8]
  assign _GEN_800 = _T_98 ? _GEN_781 : _GEN_724; // @[Bus.scala 302:73:@343.8]
  assign _GEN_801 = _T_98 ? _GEN_782 : _GEN_725; // @[Bus.scala 302:73:@343.8]
  assign _GEN_802 = _T_98 ? _GEN_783 : _GEN_726; // @[Bus.scala 302:73:@343.8]
  assign _GEN_803 = _T_97 ? _GEN_784 : _GEN_708; // @[Bus.scala 301:41:@341.6]
  assign _GEN_804 = _T_97 ? $signed(_GEN_785) : $signed(_GEN_709); // @[Bus.scala 301:41:@341.6]
  assign _GEN_805 = _T_97 ? $signed(_GEN_786) : $signed(_GEN_710); // @[Bus.scala 301:41:@341.6]
  assign _GEN_806 = _T_97 ? _GEN_787 : _GEN_711; // @[Bus.scala 301:41:@341.6]
  assign _GEN_807 = _T_97 ? _GEN_788 : _GEN_712; // @[Bus.scala 301:41:@341.6]
  assign _GEN_808 = _T_97 ? $signed(_GEN_789) : $signed(_GEN_713); // @[Bus.scala 301:41:@341.6]
  assign _GEN_809 = _T_97 ? $signed(_GEN_790) : $signed(_GEN_714); // @[Bus.scala 301:41:@341.6]
  assign _GEN_810 = _T_97 ? $signed(_GEN_791) : $signed(_GEN_715); // @[Bus.scala 301:41:@341.6]
  assign _GEN_811 = _T_97 ? _GEN_792 : _GEN_716; // @[Bus.scala 301:41:@341.6]
  assign _GEN_812 = _T_97 ? _GEN_793 : _GEN_717; // @[Bus.scala 301:41:@341.6]
  assign _GEN_813 = _T_97 ? _GEN_794 : _GEN_718; // @[Bus.scala 301:41:@341.6]
  assign _GEN_814 = _T_97 ? _GEN_795 : _GEN_719; // @[Bus.scala 301:41:@341.6]
  assign _GEN_815 = _T_97 ? _GEN_796 : _GEN_720; // @[Bus.scala 301:41:@341.6]
  assign _GEN_816 = _T_97 ? _GEN_797 : _GEN_721; // @[Bus.scala 301:41:@341.6]
  assign _GEN_817 = _T_97 ? _GEN_798 : _GEN_722; // @[Bus.scala 301:41:@341.6]
  assign _GEN_818 = _T_97 ? _GEN_799 : _GEN_723; // @[Bus.scala 301:41:@341.6]
  assign _GEN_819 = _T_97 ? _GEN_800 : _GEN_724; // @[Bus.scala 301:41:@341.6]
  assign _GEN_820 = _T_97 ? _GEN_801 : _GEN_725; // @[Bus.scala 301:41:@341.6]
  assign _GEN_821 = _T_97 ? _GEN_802 : _GEN_726; // @[Bus.scala 301:41:@341.6]
  assign _T_345 = $signed(io_master_in_addr) <= $signed(32'sh1f); // @[Bus.scala 333:65:@386.12]
  assign _T_347 = $signed(-32'sh18) + $signed(io_master_in_addr); // @[Bus.scala 336:93:@390.16]
  assign _T_348 = $signed(-32'sh18) + $signed(io_master_in_addr); // @[Bus.scala 336:93:@391.16]
  assign _T_349 = $signed(_T_348); // @[Bus.scala 336:93:@392.16]
  assign _GEN_822 = io_master_in_sync ? 4'h8 : _GEN_803; // @[Bus.scala 334:73:@388.14]
  assign _GEN_823 = io_master_in_sync ? $signed(_T_349) : $signed(_GEN_804); // @[Bus.scala 334:73:@388.14]
  assign _GEN_824 = io_master_in_sync ? $signed(io_master_in_data) : $signed(_GEN_805); // @[Bus.scala 334:73:@388.14]
  assign _GEN_825 = io_master_in_sync ? io_master_in_trans_type : _GEN_806; // @[Bus.scala 334:73:@388.14]
  assign _GEN_826 = io_master_in_sync ? resp_signal_r_ack : _GEN_807; // @[Bus.scala 334:73:@388.14]
  assign _GEN_827 = io_master_in_sync ? $signed(resp_signal_r_data) : $signed(_GEN_808); // @[Bus.scala 334:73:@388.14]
  assign _GEN_828 = io_master_in_sync ? $signed(_T_349) : $signed(slave_out3_r_addr); // @[Bus.scala 334:73:@388.14]
  assign _GEN_829 = io_master_in_sync ? $signed(io_master_in_data) : $signed(slave_out3_r_data); // @[Bus.scala 334:73:@388.14]
  assign _GEN_830 = io_master_in_sync ? io_master_in_trans_type : slave_out3_r_trans_type; // @[Bus.scala 334:73:@388.14]
  assign _GEN_831 = io_master_in_sync ? 1'h0 : _GEN_812; // @[Bus.scala 334:73:@388.14]
  assign _GEN_832 = io_master_in_sync ? 1'h0 : _GEN_813; // @[Bus.scala 334:73:@388.14]
  assign _GEN_833 = io_master_in_sync ? 1'h0 : _GEN_814; // @[Bus.scala 334:73:@388.14]
  assign _GEN_834 = io_master_in_sync ? 1'h0 : _GEN_815; // @[Bus.scala 334:73:@388.14]
  assign _GEN_835 = io_master_in_sync ? 1'h0 : _GEN_816; // @[Bus.scala 334:73:@388.14]
  assign _GEN_836 = io_master_in_sync ? 1'h0 : _GEN_817; // @[Bus.scala 334:73:@388.14]
  assign _GEN_837 = io_master_in_sync ? 1'h0 : _GEN_818; // @[Bus.scala 334:73:@388.14]
  assign _GEN_838 = io_master_in_sync ? 1'h0 : _GEN_819; // @[Bus.scala 334:73:@388.14]
  assign _GEN_839 = io_master_in_sync ? 1'h0 : _GEN_820; // @[Bus.scala 334:73:@388.14]
  assign _GEN_840 = io_master_in_sync ? 1'h1 : _GEN_821; // @[Bus.scala 334:73:@388.14]
  assign _GEN_841 = _T_345 ? _GEN_822 : _GEN_803; // @[Bus.scala 333:81:@387.12]
  assign _GEN_842 = _T_345 ? $signed(_GEN_823) : $signed(_GEN_804); // @[Bus.scala 333:81:@387.12]
  assign _GEN_843 = _T_345 ? $signed(_GEN_824) : $signed(_GEN_805); // @[Bus.scala 333:81:@387.12]
  assign _GEN_844 = _T_345 ? _GEN_825 : _GEN_806; // @[Bus.scala 333:81:@387.12]
  assign _GEN_845 = _T_345 ? _GEN_826 : _GEN_807; // @[Bus.scala 333:81:@387.12]
  assign _GEN_846 = _T_345 ? $signed(_GEN_827) : $signed(_GEN_808); // @[Bus.scala 333:81:@387.12]
  assign _GEN_847 = _T_345 ? $signed(_GEN_828) : $signed(slave_out3_r_addr); // @[Bus.scala 333:81:@387.12]
  assign _GEN_848 = _T_345 ? $signed(_GEN_829) : $signed(slave_out3_r_data); // @[Bus.scala 333:81:@387.12]
  assign _GEN_849 = _T_345 ? _GEN_830 : slave_out3_r_trans_type; // @[Bus.scala 333:81:@387.12]
  assign _GEN_850 = _T_345 ? _GEN_831 : _GEN_812; // @[Bus.scala 333:81:@387.12]
  assign _GEN_851 = _T_345 ? _GEN_832 : _GEN_813; // @[Bus.scala 333:81:@387.12]
  assign _GEN_852 = _T_345 ? _GEN_833 : _GEN_814; // @[Bus.scala 333:81:@387.12]
  assign _GEN_853 = _T_345 ? _GEN_834 : _GEN_815; // @[Bus.scala 333:81:@387.12]
  assign _GEN_854 = _T_345 ? _GEN_835 : _GEN_816; // @[Bus.scala 333:81:@387.12]
  assign _GEN_855 = _T_345 ? _GEN_836 : _GEN_817; // @[Bus.scala 333:81:@387.12]
  assign _GEN_856 = _T_345 ? _GEN_837 : _GEN_818; // @[Bus.scala 333:81:@387.12]
  assign _GEN_857 = _T_345 ? _GEN_838 : _GEN_819; // @[Bus.scala 333:81:@387.12]
  assign _GEN_858 = _T_345 ? _GEN_839 : _GEN_820; // @[Bus.scala 333:81:@387.12]
  assign _GEN_859 = _T_345 ? _GEN_840 : _GEN_821; // @[Bus.scala 333:81:@387.12]
  assign _GEN_860 = _T_163 ? _GEN_841 : _GEN_803; // @[Bus.scala 332:73:@385.10]
  assign _GEN_861 = _T_163 ? $signed(_GEN_842) : $signed(_GEN_804); // @[Bus.scala 332:73:@385.10]
  assign _GEN_862 = _T_163 ? $signed(_GEN_843) : $signed(_GEN_805); // @[Bus.scala 332:73:@385.10]
  assign _GEN_863 = _T_163 ? _GEN_844 : _GEN_806; // @[Bus.scala 332:73:@385.10]
  assign _GEN_864 = _T_163 ? _GEN_845 : _GEN_807; // @[Bus.scala 332:73:@385.10]
  assign _GEN_865 = _T_163 ? $signed(_GEN_846) : $signed(_GEN_808); // @[Bus.scala 332:73:@385.10]
  assign _GEN_866 = _T_163 ? $signed(_GEN_847) : $signed(slave_out3_r_addr); // @[Bus.scala 332:73:@385.10]
  assign _GEN_867 = _T_163 ? $signed(_GEN_848) : $signed(slave_out3_r_data); // @[Bus.scala 332:73:@385.10]
  assign _GEN_868 = _T_163 ? _GEN_849 : slave_out3_r_trans_type; // @[Bus.scala 332:73:@385.10]
  assign _GEN_869 = _T_163 ? _GEN_850 : _GEN_812; // @[Bus.scala 332:73:@385.10]
  assign _GEN_870 = _T_163 ? _GEN_851 : _GEN_813; // @[Bus.scala 332:73:@385.10]
  assign _GEN_871 = _T_163 ? _GEN_852 : _GEN_814; // @[Bus.scala 332:73:@385.10]
  assign _GEN_872 = _T_163 ? _GEN_853 : _GEN_815; // @[Bus.scala 332:73:@385.10]
  assign _GEN_873 = _T_163 ? _GEN_854 : _GEN_816; // @[Bus.scala 332:73:@385.10]
  assign _GEN_874 = _T_163 ? _GEN_855 : _GEN_817; // @[Bus.scala 332:73:@385.10]
  assign _GEN_875 = _T_163 ? _GEN_856 : _GEN_818; // @[Bus.scala 332:73:@385.10]
  assign _GEN_876 = _T_163 ? _GEN_857 : _GEN_819; // @[Bus.scala 332:73:@385.10]
  assign _GEN_877 = _T_163 ? _GEN_858 : _GEN_820; // @[Bus.scala 332:73:@385.10]
  assign _GEN_878 = _T_163 ? _GEN_859 : _GEN_821; // @[Bus.scala 332:73:@385.10]
  assign _GEN_879 = _T_100 ? _GEN_860 : _GEN_803; // @[Bus.scala 331:74:@383.8]
  assign _GEN_880 = _T_100 ? $signed(_GEN_861) : $signed(_GEN_804); // @[Bus.scala 331:74:@383.8]
  assign _GEN_881 = _T_100 ? $signed(_GEN_862) : $signed(_GEN_805); // @[Bus.scala 331:74:@383.8]
  assign _GEN_882 = _T_100 ? _GEN_863 : _GEN_806; // @[Bus.scala 331:74:@383.8]
  assign _GEN_883 = _T_100 ? _GEN_864 : _GEN_807; // @[Bus.scala 331:74:@383.8]
  assign _GEN_884 = _T_100 ? $signed(_GEN_865) : $signed(_GEN_808); // @[Bus.scala 331:74:@383.8]
  assign _GEN_885 = _T_100 ? $signed(_GEN_866) : $signed(slave_out3_r_addr); // @[Bus.scala 331:74:@383.8]
  assign _GEN_886 = _T_100 ? $signed(_GEN_867) : $signed(slave_out3_r_data); // @[Bus.scala 331:74:@383.8]
  assign _GEN_887 = _T_100 ? _GEN_868 : slave_out3_r_trans_type; // @[Bus.scala 331:74:@383.8]
  assign _GEN_888 = _T_100 ? _GEN_869 : _GEN_812; // @[Bus.scala 331:74:@383.8]
  assign _GEN_889 = _T_100 ? _GEN_870 : _GEN_813; // @[Bus.scala 331:74:@383.8]
  assign _GEN_890 = _T_100 ? _GEN_871 : _GEN_814; // @[Bus.scala 331:74:@383.8]
  assign _GEN_891 = _T_100 ? _GEN_872 : _GEN_815; // @[Bus.scala 331:74:@383.8]
  assign _GEN_892 = _T_100 ? _GEN_873 : _GEN_816; // @[Bus.scala 331:74:@383.8]
  assign _GEN_893 = _T_100 ? _GEN_874 : _GEN_817; // @[Bus.scala 331:74:@383.8]
  assign _GEN_894 = _T_100 ? _GEN_875 : _GEN_818; // @[Bus.scala 331:74:@383.8]
  assign _GEN_895 = _T_100 ? _GEN_876 : _GEN_819; // @[Bus.scala 331:74:@383.8]
  assign _GEN_896 = _T_100 ? _GEN_877 : _GEN_820; // @[Bus.scala 331:74:@383.8]
  assign _GEN_897 = _T_100 ? _GEN_878 : _GEN_821; // @[Bus.scala 331:74:@383.8]
  assign _GEN_898 = _T_97 ? _GEN_879 : _GEN_803; // @[Bus.scala 330:41:@380.6]
  assign _GEN_899 = _T_97 ? $signed(_GEN_880) : $signed(_GEN_804); // @[Bus.scala 330:41:@380.6]
  assign _GEN_900 = _T_97 ? $signed(_GEN_881) : $signed(_GEN_805); // @[Bus.scala 330:41:@380.6]
  assign _GEN_901 = _T_97 ? _GEN_882 : _GEN_806; // @[Bus.scala 330:41:@380.6]
  assign _GEN_902 = _T_97 ? _GEN_883 : _GEN_807; // @[Bus.scala 330:41:@380.6]
  assign _GEN_903 = _T_97 ? $signed(_GEN_884) : $signed(_GEN_808); // @[Bus.scala 330:41:@380.6]
  assign _GEN_904 = _T_97 ? $signed(_GEN_885) : $signed(slave_out3_r_addr); // @[Bus.scala 330:41:@380.6]
  assign _GEN_905 = _T_97 ? $signed(_GEN_886) : $signed(slave_out3_r_data); // @[Bus.scala 330:41:@380.6]
  assign _GEN_906 = _T_97 ? _GEN_887 : slave_out3_r_trans_type; // @[Bus.scala 330:41:@380.6]
  assign _GEN_907 = _T_97 ? _GEN_888 : _GEN_812; // @[Bus.scala 330:41:@380.6]
  assign _GEN_908 = _T_97 ? _GEN_889 : _GEN_813; // @[Bus.scala 330:41:@380.6]
  assign _GEN_909 = _T_97 ? _GEN_890 : _GEN_814; // @[Bus.scala 330:41:@380.6]
  assign _GEN_910 = _T_97 ? _GEN_891 : _GEN_815; // @[Bus.scala 330:41:@380.6]
  assign _GEN_911 = _T_97 ? _GEN_892 : _GEN_816; // @[Bus.scala 330:41:@380.6]
  assign _GEN_912 = _T_97 ? _GEN_893 : _GEN_817; // @[Bus.scala 330:41:@380.6]
  assign _GEN_913 = _T_97 ? _GEN_894 : _GEN_818; // @[Bus.scala 330:41:@380.6]
  assign _GEN_914 = _T_97 ? _GEN_895 : _GEN_819; // @[Bus.scala 330:41:@380.6]
  assign _GEN_915 = _T_97 ? _GEN_896 : _GEN_820; // @[Bus.scala 330:41:@380.6]
  assign _GEN_916 = _T_97 ? _GEN_897 : _GEN_821; // @[Bus.scala 330:41:@380.6]
  assign _GEN_917 = io_master_in_sync ? 4'h8 : _GEN_898; // @[Bus.scala 363:73:@427.14]
  assign _GEN_918 = io_master_in_sync ? $signed(_T_349) : $signed(_GEN_899); // @[Bus.scala 363:73:@427.14]
  assign _GEN_919 = io_master_in_sync ? $signed(32'sh0) : $signed(_GEN_900); // @[Bus.scala 363:73:@427.14]
  assign _GEN_920 = io_master_in_sync ? io_master_in_trans_type : _GEN_901; // @[Bus.scala 363:73:@427.14]
  assign _GEN_921 = io_master_in_sync ? resp_signal_r_ack : _GEN_902; // @[Bus.scala 363:73:@427.14]
  assign _GEN_922 = io_master_in_sync ? $signed(resp_signal_r_data) : $signed(_GEN_903); // @[Bus.scala 363:73:@427.14]
  assign _GEN_923 = io_master_in_sync ? $signed(_T_349) : $signed(_GEN_904); // @[Bus.scala 363:73:@427.14]
  assign _GEN_924 = io_master_in_sync ? $signed(32'sh0) : $signed(_GEN_905); // @[Bus.scala 363:73:@427.14]
  assign _GEN_925 = io_master_in_sync ? io_master_in_trans_type : _GEN_906; // @[Bus.scala 363:73:@427.14]
  assign _GEN_926 = io_master_in_sync ? 1'h0 : _GEN_907; // @[Bus.scala 363:73:@427.14]
  assign _GEN_927 = io_master_in_sync ? 1'h0 : _GEN_908; // @[Bus.scala 363:73:@427.14]
  assign _GEN_928 = io_master_in_sync ? 1'h0 : _GEN_909; // @[Bus.scala 363:73:@427.14]
  assign _GEN_929 = io_master_in_sync ? 1'h0 : _GEN_910; // @[Bus.scala 363:73:@427.14]
  assign _GEN_930 = io_master_in_sync ? 1'h0 : _GEN_911; // @[Bus.scala 363:73:@427.14]
  assign _GEN_931 = io_master_in_sync ? 1'h0 : _GEN_912; // @[Bus.scala 363:73:@427.14]
  assign _GEN_932 = io_master_in_sync ? 1'h0 : _GEN_913; // @[Bus.scala 363:73:@427.14]
  assign _GEN_933 = io_master_in_sync ? 1'h0 : _GEN_914; // @[Bus.scala 363:73:@427.14]
  assign _GEN_934 = io_master_in_sync ? 1'h0 : _GEN_915; // @[Bus.scala 363:73:@427.14]
  assign _GEN_935 = io_master_in_sync ? 1'h1 : _GEN_916; // @[Bus.scala 363:73:@427.14]
  assign _GEN_936 = _T_345 ? _GEN_917 : _GEN_898; // @[Bus.scala 362:81:@426.12]
  assign _GEN_937 = _T_345 ? $signed(_GEN_918) : $signed(_GEN_899); // @[Bus.scala 362:81:@426.12]
  assign _GEN_938 = _T_345 ? $signed(_GEN_919) : $signed(_GEN_900); // @[Bus.scala 362:81:@426.12]
  assign _GEN_939 = _T_345 ? _GEN_920 : _GEN_901; // @[Bus.scala 362:81:@426.12]
  assign _GEN_940 = _T_345 ? _GEN_921 : _GEN_902; // @[Bus.scala 362:81:@426.12]
  assign _GEN_941 = _T_345 ? $signed(_GEN_922) : $signed(_GEN_903); // @[Bus.scala 362:81:@426.12]
  assign _GEN_942 = _T_345 ? $signed(_GEN_923) : $signed(_GEN_904); // @[Bus.scala 362:81:@426.12]
  assign _GEN_943 = _T_345 ? $signed(_GEN_924) : $signed(_GEN_905); // @[Bus.scala 362:81:@426.12]
  assign _GEN_944 = _T_345 ? _GEN_925 : _GEN_906; // @[Bus.scala 362:81:@426.12]
  assign _GEN_945 = _T_345 ? _GEN_926 : _GEN_907; // @[Bus.scala 362:81:@426.12]
  assign _GEN_946 = _T_345 ? _GEN_927 : _GEN_908; // @[Bus.scala 362:81:@426.12]
  assign _GEN_947 = _T_345 ? _GEN_928 : _GEN_909; // @[Bus.scala 362:81:@426.12]
  assign _GEN_948 = _T_345 ? _GEN_929 : _GEN_910; // @[Bus.scala 362:81:@426.12]
  assign _GEN_949 = _T_345 ? _GEN_930 : _GEN_911; // @[Bus.scala 362:81:@426.12]
  assign _GEN_950 = _T_345 ? _GEN_931 : _GEN_912; // @[Bus.scala 362:81:@426.12]
  assign _GEN_951 = _T_345 ? _GEN_932 : _GEN_913; // @[Bus.scala 362:81:@426.12]
  assign _GEN_952 = _T_345 ? _GEN_933 : _GEN_914; // @[Bus.scala 362:81:@426.12]
  assign _GEN_953 = _T_345 ? _GEN_934 : _GEN_915; // @[Bus.scala 362:81:@426.12]
  assign _GEN_954 = _T_345 ? _GEN_935 : _GEN_916; // @[Bus.scala 362:81:@426.12]
  assign _GEN_955 = _T_163 ? _GEN_936 : _GEN_898; // @[Bus.scala 361:73:@424.10]
  assign _GEN_956 = _T_163 ? $signed(_GEN_937) : $signed(_GEN_899); // @[Bus.scala 361:73:@424.10]
  assign _GEN_957 = _T_163 ? $signed(_GEN_938) : $signed(_GEN_900); // @[Bus.scala 361:73:@424.10]
  assign _GEN_958 = _T_163 ? _GEN_939 : _GEN_901; // @[Bus.scala 361:73:@424.10]
  assign _GEN_959 = _T_163 ? _GEN_940 : _GEN_902; // @[Bus.scala 361:73:@424.10]
  assign _GEN_960 = _T_163 ? $signed(_GEN_941) : $signed(_GEN_903); // @[Bus.scala 361:73:@424.10]
  assign _GEN_961 = _T_163 ? $signed(_GEN_942) : $signed(_GEN_904); // @[Bus.scala 361:73:@424.10]
  assign _GEN_962 = _T_163 ? $signed(_GEN_943) : $signed(_GEN_905); // @[Bus.scala 361:73:@424.10]
  assign _GEN_963 = _T_163 ? _GEN_944 : _GEN_906; // @[Bus.scala 361:73:@424.10]
  assign _GEN_964 = _T_163 ? _GEN_945 : _GEN_907; // @[Bus.scala 361:73:@424.10]
  assign _GEN_965 = _T_163 ? _GEN_946 : _GEN_908; // @[Bus.scala 361:73:@424.10]
  assign _GEN_966 = _T_163 ? _GEN_947 : _GEN_909; // @[Bus.scala 361:73:@424.10]
  assign _GEN_967 = _T_163 ? _GEN_948 : _GEN_910; // @[Bus.scala 361:73:@424.10]
  assign _GEN_968 = _T_163 ? _GEN_949 : _GEN_911; // @[Bus.scala 361:73:@424.10]
  assign _GEN_969 = _T_163 ? _GEN_950 : _GEN_912; // @[Bus.scala 361:73:@424.10]
  assign _GEN_970 = _T_163 ? _GEN_951 : _GEN_913; // @[Bus.scala 361:73:@424.10]
  assign _GEN_971 = _T_163 ? _GEN_952 : _GEN_914; // @[Bus.scala 361:73:@424.10]
  assign _GEN_972 = _T_163 ? _GEN_953 : _GEN_915; // @[Bus.scala 361:73:@424.10]
  assign _GEN_973 = _T_163 ? _GEN_954 : _GEN_916; // @[Bus.scala 361:73:@424.10]
  assign _GEN_974 = _T_98 ? _GEN_955 : _GEN_898; // @[Bus.scala 360:73:@422.8]
  assign _GEN_975 = _T_98 ? $signed(_GEN_956) : $signed(_GEN_899); // @[Bus.scala 360:73:@422.8]
  assign _GEN_976 = _T_98 ? $signed(_GEN_957) : $signed(_GEN_900); // @[Bus.scala 360:73:@422.8]
  assign _GEN_977 = _T_98 ? _GEN_958 : _GEN_901; // @[Bus.scala 360:73:@422.8]
  assign _GEN_978 = _T_98 ? _GEN_959 : _GEN_902; // @[Bus.scala 360:73:@422.8]
  assign _GEN_979 = _T_98 ? $signed(_GEN_960) : $signed(_GEN_903); // @[Bus.scala 360:73:@422.8]
  assign _GEN_980 = _T_98 ? $signed(_GEN_961) : $signed(_GEN_904); // @[Bus.scala 360:73:@422.8]
  assign _GEN_981 = _T_98 ? $signed(_GEN_962) : $signed(_GEN_905); // @[Bus.scala 360:73:@422.8]
  assign _GEN_982 = _T_98 ? _GEN_963 : _GEN_906; // @[Bus.scala 360:73:@422.8]
  assign _GEN_983 = _T_98 ? _GEN_964 : _GEN_907; // @[Bus.scala 360:73:@422.8]
  assign _GEN_984 = _T_98 ? _GEN_965 : _GEN_908; // @[Bus.scala 360:73:@422.8]
  assign _GEN_985 = _T_98 ? _GEN_966 : _GEN_909; // @[Bus.scala 360:73:@422.8]
  assign _GEN_986 = _T_98 ? _GEN_967 : _GEN_910; // @[Bus.scala 360:73:@422.8]
  assign _GEN_987 = _T_98 ? _GEN_968 : _GEN_911; // @[Bus.scala 360:73:@422.8]
  assign _GEN_988 = _T_98 ? _GEN_969 : _GEN_912; // @[Bus.scala 360:73:@422.8]
  assign _GEN_989 = _T_98 ? _GEN_970 : _GEN_913; // @[Bus.scala 360:73:@422.8]
  assign _GEN_990 = _T_98 ? _GEN_971 : _GEN_914; // @[Bus.scala 360:73:@422.8]
  assign _GEN_991 = _T_98 ? _GEN_972 : _GEN_915; // @[Bus.scala 360:73:@422.8]
  assign _GEN_992 = _T_98 ? _GEN_973 : _GEN_916; // @[Bus.scala 360:73:@422.8]
  assign _GEN_993 = _T_97 ? _GEN_974 : _GEN_898; // @[Bus.scala 359:41:@420.6]
  assign _GEN_994 = _T_97 ? $signed(_GEN_975) : $signed(_GEN_899); // @[Bus.scala 359:41:@420.6]
  assign _GEN_995 = _T_97 ? $signed(_GEN_976) : $signed(_GEN_900); // @[Bus.scala 359:41:@420.6]
  assign _GEN_996 = _T_97 ? _GEN_977 : _GEN_901; // @[Bus.scala 359:41:@420.6]
  assign _GEN_997 = _T_97 ? _GEN_978 : _GEN_902; // @[Bus.scala 359:41:@420.6]
  assign _GEN_998 = _T_97 ? $signed(_GEN_979) : $signed(_GEN_903); // @[Bus.scala 359:41:@420.6]
  assign _GEN_999 = _T_97 ? $signed(_GEN_980) : $signed(_GEN_904); // @[Bus.scala 359:41:@420.6]
  assign _GEN_1000 = _T_97 ? $signed(_GEN_981) : $signed(_GEN_905); // @[Bus.scala 359:41:@420.6]
  assign _GEN_1001 = _T_97 ? _GEN_982 : _GEN_906; // @[Bus.scala 359:41:@420.6]
  assign _GEN_1002 = _T_97 ? _GEN_983 : _GEN_907; // @[Bus.scala 359:41:@420.6]
  assign _GEN_1003 = _T_97 ? _GEN_984 : _GEN_908; // @[Bus.scala 359:41:@420.6]
  assign _GEN_1004 = _T_97 ? _GEN_985 : _GEN_909; // @[Bus.scala 359:41:@420.6]
  assign _GEN_1005 = _T_97 ? _GEN_986 : _GEN_910; // @[Bus.scala 359:41:@420.6]
  assign _GEN_1006 = _T_97 ? _GEN_987 : _GEN_911; // @[Bus.scala 359:41:@420.6]
  assign _GEN_1007 = _T_97 ? _GEN_988 : _GEN_912; // @[Bus.scala 359:41:@420.6]
  assign _GEN_1008 = _T_97 ? _GEN_989 : _GEN_913; // @[Bus.scala 359:41:@420.6]
  assign _GEN_1009 = _T_97 ? _GEN_990 : _GEN_914; // @[Bus.scala 359:41:@420.6]
  assign _GEN_1010 = _T_97 ? _GEN_991 : _GEN_915; // @[Bus.scala 359:41:@420.6]
  assign _GEN_1011 = _T_97 ? _GEN_992 : _GEN_916; // @[Bus.scala 359:41:@420.6]
  assign _T_390 = state_r == 4'h1; // @[Bus.scala 388:30:@458.6]
  assign _GEN_1012 = io_slave_out0_sync ? 4'h2 : _GEN_993; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1013 = io_slave_out0_sync ? $signed(req_signal_r_addr) : $signed(_GEN_994); // @[Bus.scala 389:50:@460.8]
  assign _GEN_1014 = io_slave_out0_sync ? $signed(req_signal_r_data) : $signed(_GEN_995); // @[Bus.scala 389:50:@460.8]
  assign _GEN_1015 = io_slave_out0_sync ? req_signal_r_trans_type : _GEN_996; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1016 = io_slave_out0_sync ? resp_signal_r_ack : _GEN_997; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1017 = io_slave_out0_sync ? $signed(resp_signal_r_data) : $signed(_GEN_998); // @[Bus.scala 389:50:@460.8]
  assign _GEN_1018 = io_slave_out0_sync ? 1'h0 : _GEN_1002; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1019 = io_slave_out0_sync ? 1'h0 : _GEN_1003; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1020 = io_slave_out0_sync ? 1'h1 : _GEN_1004; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1021 = io_slave_out0_sync ? 1'h0 : _GEN_1005; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1022 = io_slave_out0_sync ? 1'h0 : _GEN_1006; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1023 = io_slave_out0_sync ? 1'h0 : _GEN_1007; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1024 = io_slave_out0_sync ? 1'h0 : _GEN_1008; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1025 = io_slave_out0_sync ? 1'h0 : _GEN_1009; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1026 = io_slave_out0_sync ? 1'h0 : _GEN_1010; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1027 = io_slave_out0_sync ? 1'h0 : _GEN_1011; // @[Bus.scala 389:50:@460.8]
  assign _GEN_1028 = _T_390 ? _GEN_1012 : _GEN_993; // @[Bus.scala 388:41:@459.6]
  assign _GEN_1029 = _T_390 ? $signed(_GEN_1013) : $signed(_GEN_994); // @[Bus.scala 388:41:@459.6]
  assign _GEN_1030 = _T_390 ? $signed(_GEN_1014) : $signed(_GEN_995); // @[Bus.scala 388:41:@459.6]
  assign _GEN_1031 = _T_390 ? _GEN_1015 : _GEN_996; // @[Bus.scala 388:41:@459.6]
  assign _GEN_1032 = _T_390 ? _GEN_1016 : _GEN_997; // @[Bus.scala 388:41:@459.6]
  assign _GEN_1033 = _T_390 ? $signed(_GEN_1017) : $signed(_GEN_998); // @[Bus.scala 388:41:@459.6]
  assign _GEN_1034 = _T_390 ? _GEN_1018 : _GEN_1002; // @[Bus.scala 388:41:@459.6]
  assign _GEN_1035 = _T_390 ? _GEN_1019 : _GEN_1003; // @[Bus.scala 388:41:@459.6]
  assign _GEN_1036 = _T_390 ? _GEN_1020 : _GEN_1004; // @[Bus.scala 388:41:@459.6]
  assign _GEN_1037 = _T_390 ? _GEN_1021 : _GEN_1005; // @[Bus.scala 388:41:@459.6]
  assign _GEN_1038 = _T_390 ? _GEN_1022 : _GEN_1006; // @[Bus.scala 388:41:@459.6]
  assign _GEN_1039 = _T_390 ? _GEN_1023 : _GEN_1007; // @[Bus.scala 388:41:@459.6]
  assign _GEN_1040 = _T_390 ? _GEN_1024 : _GEN_1008; // @[Bus.scala 388:41:@459.6]
  assign _GEN_1041 = _T_390 ? _GEN_1025 : _GEN_1009; // @[Bus.scala 388:41:@459.6]
  assign _GEN_1042 = _T_390 ? _GEN_1026 : _GEN_1010; // @[Bus.scala 388:41:@459.6]
  assign _GEN_1043 = _T_390 ? _GEN_1027 : _GEN_1011; // @[Bus.scala 388:41:@459.6]
  assign _T_401 = state_r == 4'h2; // @[Bus.scala 408:30:@479.6]
  assign _T_402 = 32'h1 == req_signal_r_trans_type; // @[Bus.scala 409:45:@481.8]
  assign _T_404 = _T_402 == 1'h0; // @[Bus.scala 409:30:@482.8]
  assign _GEN_1044 = io_slave_in0_sync ? 4'h3 : _GEN_1028; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1045 = io_slave_in0_sync ? io_slave_in0_ack : _GEN_425; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1046 = io_slave_in0_sync ? $signed(io_slave_in0_data) : $signed(_GEN_426); // @[Bus.scala 410:57:@484.10]
  assign _GEN_1047 = io_slave_in0_sync ? $signed(req_signal_r_addr) : $signed(_GEN_1029); // @[Bus.scala 410:57:@484.10]
  assign _GEN_1048 = io_slave_in0_sync ? $signed(req_signal_r_data) : $signed(_GEN_1030); // @[Bus.scala 410:57:@484.10]
  assign _GEN_1049 = io_slave_in0_sync ? req_signal_r_trans_type : _GEN_1031; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1050 = io_slave_in0_sync ? io_slave_in0_ack : _GEN_1032; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1051 = io_slave_in0_sync ? $signed(io_slave_in0_data) : $signed(_GEN_1033); // @[Bus.scala 410:57:@484.10]
  assign _GEN_1052 = io_slave_in0_sync ? 1'h0 : _GEN_1034; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1053 = io_slave_in0_sync ? 1'h1 : _GEN_1035; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1054 = io_slave_in0_sync ? 1'h0 : _GEN_1036; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1055 = io_slave_in0_sync ? 1'h0 : _GEN_1037; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1056 = io_slave_in0_sync ? 1'h0 : _GEN_1038; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1057 = io_slave_in0_sync ? 1'h0 : _GEN_1039; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1058 = io_slave_in0_sync ? 1'h0 : _GEN_1040; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1059 = io_slave_in0_sync ? 1'h0 : _GEN_1041; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1060 = io_slave_in0_sync ? 1'h0 : _GEN_1042; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1061 = io_slave_in0_sync ? 1'h0 : _GEN_1043; // @[Bus.scala 410:57:@484.10]
  assign _GEN_1062 = _T_404 ? _GEN_1044 : _GEN_1028; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1063 = _T_404 ? _GEN_1045 : _GEN_425; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1064 = _T_404 ? $signed(_GEN_1046) : $signed(_GEN_426); // @[Bus.scala 409:75:@483.8]
  assign _GEN_1065 = _T_404 ? $signed(_GEN_1047) : $signed(_GEN_1029); // @[Bus.scala 409:75:@483.8]
  assign _GEN_1066 = _T_404 ? $signed(_GEN_1048) : $signed(_GEN_1030); // @[Bus.scala 409:75:@483.8]
  assign _GEN_1067 = _T_404 ? _GEN_1049 : _GEN_1031; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1068 = _T_404 ? _GEN_1050 : _GEN_1032; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1069 = _T_404 ? $signed(_GEN_1051) : $signed(_GEN_1033); // @[Bus.scala 409:75:@483.8]
  assign _GEN_1070 = _T_404 ? _GEN_1052 : _GEN_1034; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1071 = _T_404 ? _GEN_1053 : _GEN_1035; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1072 = _T_404 ? _GEN_1054 : _GEN_1036; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1073 = _T_404 ? _GEN_1055 : _GEN_1037; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1074 = _T_404 ? _GEN_1056 : _GEN_1038; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1075 = _T_404 ? _GEN_1057 : _GEN_1039; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1076 = _T_404 ? _GEN_1058 : _GEN_1040; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1077 = _T_404 ? _GEN_1059 : _GEN_1041; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1078 = _T_404 ? _GEN_1060 : _GEN_1042; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1079 = _T_404 ? _GEN_1061 : _GEN_1043; // @[Bus.scala 409:75:@483.8]
  assign _GEN_1080 = _T_401 ? _GEN_1062 : _GEN_1028; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1081 = _T_401 ? _GEN_1063 : _GEN_425; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1082 = _T_401 ? $signed(_GEN_1064) : $signed(_GEN_426); // @[Bus.scala 408:41:@480.6]
  assign _GEN_1083 = _T_401 ? $signed(_GEN_1065) : $signed(_GEN_1029); // @[Bus.scala 408:41:@480.6]
  assign _GEN_1084 = _T_401 ? $signed(_GEN_1066) : $signed(_GEN_1030); // @[Bus.scala 408:41:@480.6]
  assign _GEN_1085 = _T_401 ? _GEN_1067 : _GEN_1031; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1086 = _T_401 ? _GEN_1068 : _GEN_1032; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1087 = _T_401 ? $signed(_GEN_1069) : $signed(_GEN_1033); // @[Bus.scala 408:41:@480.6]
  assign _GEN_1088 = _T_401 ? _GEN_1070 : _GEN_1034; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1089 = _T_401 ? _GEN_1071 : _GEN_1035; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1090 = _T_401 ? _GEN_1072 : _GEN_1036; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1091 = _T_401 ? _GEN_1073 : _GEN_1037; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1092 = _T_401 ? _GEN_1074 : _GEN_1038; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1093 = _T_401 ? _GEN_1075 : _GEN_1039; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1094 = _T_401 ? _GEN_1076 : _GEN_1040; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1095 = _T_401 ? _GEN_1077 : _GEN_1041; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1096 = _T_401 ? _GEN_1078 : _GEN_1042; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1097 = _T_401 ? _GEN_1079 : _GEN_1043; // @[Bus.scala 408:41:@480.6]
  assign _GEN_1098 = io_slave_in0_sync ? 4'h3 : _GEN_1080; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1099 = io_slave_in0_sync ? io_slave_in0_ack : _GEN_1081; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1100 = io_slave_in0_sync ? $signed(32'sh0) : $signed(_GEN_1082); // @[Bus.scala 434:57:@510.10]
  assign _GEN_1101 = io_slave_in0_sync ? $signed(req_signal_r_addr) : $signed(_GEN_1083); // @[Bus.scala 434:57:@510.10]
  assign _GEN_1102 = io_slave_in0_sync ? $signed(req_signal_r_data) : $signed(_GEN_1084); // @[Bus.scala 434:57:@510.10]
  assign _GEN_1103 = io_slave_in0_sync ? req_signal_r_trans_type : _GEN_1085; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1104 = io_slave_in0_sync ? io_slave_in0_ack : _GEN_1086; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1105 = io_slave_in0_sync ? $signed(32'sh0) : $signed(_GEN_1087); // @[Bus.scala 434:57:@510.10]
  assign _GEN_1106 = io_slave_in0_sync ? 1'h0 : _GEN_1088; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1107 = io_slave_in0_sync ? 1'h1 : _GEN_1089; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1108 = io_slave_in0_sync ? 1'h0 : _GEN_1090; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1109 = io_slave_in0_sync ? 1'h0 : _GEN_1091; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1110 = io_slave_in0_sync ? 1'h0 : _GEN_1092; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1111 = io_slave_in0_sync ? 1'h0 : _GEN_1093; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1112 = io_slave_in0_sync ? 1'h0 : _GEN_1094; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1113 = io_slave_in0_sync ? 1'h0 : _GEN_1095; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1114 = io_slave_in0_sync ? 1'h0 : _GEN_1096; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1115 = io_slave_in0_sync ? 1'h0 : _GEN_1097; // @[Bus.scala 434:57:@510.10]
  assign _GEN_1116 = _T_402 ? _GEN_1098 : _GEN_1080; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1117 = _T_402 ? _GEN_1099 : _GEN_1081; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1118 = _T_402 ? $signed(_GEN_1100) : $signed(_GEN_1082); // @[Bus.scala 433:74:@509.8]
  assign _GEN_1119 = _T_402 ? $signed(_GEN_1101) : $signed(_GEN_1083); // @[Bus.scala 433:74:@509.8]
  assign _GEN_1120 = _T_402 ? $signed(_GEN_1102) : $signed(_GEN_1084); // @[Bus.scala 433:74:@509.8]
  assign _GEN_1121 = _T_402 ? _GEN_1103 : _GEN_1085; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1122 = _T_402 ? _GEN_1104 : _GEN_1086; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1123 = _T_402 ? $signed(_GEN_1105) : $signed(_GEN_1087); // @[Bus.scala 433:74:@509.8]
  assign _GEN_1124 = _T_402 ? _GEN_1106 : _GEN_1088; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1125 = _T_402 ? _GEN_1107 : _GEN_1089; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1126 = _T_402 ? _GEN_1108 : _GEN_1090; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1127 = _T_402 ? _GEN_1109 : _GEN_1091; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1128 = _T_402 ? _GEN_1110 : _GEN_1092; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1129 = _T_402 ? _GEN_1111 : _GEN_1093; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1130 = _T_402 ? _GEN_1112 : _GEN_1094; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1131 = _T_402 ? _GEN_1113 : _GEN_1095; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1132 = _T_402 ? _GEN_1114 : _GEN_1096; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1133 = _T_402 ? _GEN_1115 : _GEN_1097; // @[Bus.scala 433:74:@509.8]
  assign _GEN_1134 = _T_401 ? _GEN_1116 : _GEN_1080; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1135 = _T_401 ? _GEN_1117 : _GEN_1081; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1136 = _T_401 ? $signed(_GEN_1118) : $signed(_GEN_1082); // @[Bus.scala 432:41:@507.6]
  assign _GEN_1137 = _T_401 ? $signed(_GEN_1119) : $signed(_GEN_1083); // @[Bus.scala 432:41:@507.6]
  assign _GEN_1138 = _T_401 ? $signed(_GEN_1120) : $signed(_GEN_1084); // @[Bus.scala 432:41:@507.6]
  assign _GEN_1139 = _T_401 ? _GEN_1121 : _GEN_1085; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1140 = _T_401 ? _GEN_1122 : _GEN_1086; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1141 = _T_401 ? $signed(_GEN_1123) : $signed(_GEN_1087); // @[Bus.scala 432:41:@507.6]
  assign _GEN_1142 = _T_401 ? _GEN_1124 : _GEN_1088; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1143 = _T_401 ? _GEN_1125 : _GEN_1089; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1144 = _T_401 ? _GEN_1126 : _GEN_1090; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1145 = _T_401 ? _GEN_1127 : _GEN_1091; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1146 = _T_401 ? _GEN_1128 : _GEN_1092; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1147 = _T_401 ? _GEN_1129 : _GEN_1093; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1148 = _T_401 ? _GEN_1130 : _GEN_1094; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1149 = _T_401 ? _GEN_1131 : _GEN_1095; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1150 = _T_401 ? _GEN_1132 : _GEN_1096; // @[Bus.scala 432:41:@507.6]
  assign _GEN_1151 = _T_401 ? _GEN_1133 : _GEN_1097; // @[Bus.scala 432:41:@507.6]
  assign _T_429 = state_r == 4'h3; // @[Bus.scala 456:30:@532.6]
  assign _GEN_1152 = io_master_out_sync ? 4'h0 : _GEN_1134; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1153 = io_master_out_sync ? $signed(req_signal_r_addr) : $signed(_GEN_1137); // @[Bus.scala 457:50:@534.8]
  assign _GEN_1154 = io_master_out_sync ? $signed(req_signal_r_data) : $signed(_GEN_1138); // @[Bus.scala 457:50:@534.8]
  assign _GEN_1155 = io_master_out_sync ? req_signal_r_trans_type : _GEN_1139; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1156 = io_master_out_sync ? resp_signal_r_ack : _GEN_1140; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1157 = io_master_out_sync ? $signed(resp_signal_r_data) : $signed(_GEN_1141); // @[Bus.scala 457:50:@534.8]
  assign _GEN_1158 = io_master_out_sync ? 1'h1 : _GEN_1142; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1159 = io_master_out_sync ? 1'h0 : _GEN_1143; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1160 = io_master_out_sync ? 1'h0 : _GEN_1144; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1161 = io_master_out_sync ? 1'h0 : _GEN_1145; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1162 = io_master_out_sync ? 1'h0 : _GEN_1146; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1163 = io_master_out_sync ? 1'h0 : _GEN_1147; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1164 = io_master_out_sync ? 1'h0 : _GEN_1148; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1165 = io_master_out_sync ? 1'h0 : _GEN_1149; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1166 = io_master_out_sync ? 1'h0 : _GEN_1150; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1167 = io_master_out_sync ? 1'h0 : _GEN_1151; // @[Bus.scala 457:50:@534.8]
  assign _GEN_1168 = _T_429 ? _GEN_1152 : _GEN_1134; // @[Bus.scala 456:41:@533.6]
  assign _GEN_1169 = _T_429 ? $signed(_GEN_1153) : $signed(_GEN_1137); // @[Bus.scala 456:41:@533.6]
  assign _GEN_1170 = _T_429 ? $signed(_GEN_1154) : $signed(_GEN_1138); // @[Bus.scala 456:41:@533.6]
  assign _GEN_1171 = _T_429 ? _GEN_1155 : _GEN_1139; // @[Bus.scala 456:41:@533.6]
  assign _GEN_1172 = _T_429 ? _GEN_1156 : _GEN_1140; // @[Bus.scala 456:41:@533.6]
  assign _GEN_1173 = _T_429 ? $signed(_GEN_1157) : $signed(_GEN_1141); // @[Bus.scala 456:41:@533.6]
  assign _GEN_1174 = _T_429 ? _GEN_1158 : _GEN_1142; // @[Bus.scala 456:41:@533.6]
  assign _GEN_1175 = _T_429 ? _GEN_1159 : _GEN_1143; // @[Bus.scala 456:41:@533.6]
  assign _GEN_1176 = _T_429 ? _GEN_1160 : _GEN_1144; // @[Bus.scala 456:41:@533.6]
  assign _GEN_1177 = _T_429 ? _GEN_1161 : _GEN_1145; // @[Bus.scala 456:41:@533.6]
  assign _GEN_1178 = _T_429 ? _GEN_1162 : _GEN_1146; // @[Bus.scala 456:41:@533.6]
  assign _GEN_1179 = _T_429 ? _GEN_1163 : _GEN_1147; // @[Bus.scala 456:41:@533.6]
  assign _GEN_1180 = _T_429 ? _GEN_1164 : _GEN_1148; // @[Bus.scala 456:41:@533.6]
  assign _GEN_1181 = _T_429 ? _GEN_1165 : _GEN_1149; // @[Bus.scala 456:41:@533.6]
  assign _GEN_1182 = _T_429 ? _GEN_1166 : _GEN_1150; // @[Bus.scala 456:41:@533.6]
  assign _GEN_1183 = _T_429 ? _GEN_1167 : _GEN_1151; // @[Bus.scala 456:41:@533.6]
  assign _T_440 = state_r == 4'h4; // @[Bus.scala 476:30:@553.6]
  assign _GEN_1184 = io_slave_out1_sync ? 4'h5 : _GEN_1168; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1185 = io_slave_out1_sync ? $signed(req_signal_r_addr) : $signed(_GEN_1169); // @[Bus.scala 477:50:@555.8]
  assign _GEN_1186 = io_slave_out1_sync ? $signed(req_signal_r_data) : $signed(_GEN_1170); // @[Bus.scala 477:50:@555.8]
  assign _GEN_1187 = io_slave_out1_sync ? req_signal_r_trans_type : _GEN_1171; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1188 = io_slave_out1_sync ? resp_signal_r_ack : _GEN_1172; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1189 = io_slave_out1_sync ? $signed(resp_signal_r_data) : $signed(_GEN_1173); // @[Bus.scala 477:50:@555.8]
  assign _GEN_1190 = io_slave_out1_sync ? 1'h0 : _GEN_1174; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1191 = io_slave_out1_sync ? 1'h0 : _GEN_1175; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1192 = io_slave_out1_sync ? 1'h0 : _GEN_1176; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1193 = io_slave_out1_sync ? 1'h1 : _GEN_1177; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1194 = io_slave_out1_sync ? 1'h0 : _GEN_1178; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1195 = io_slave_out1_sync ? 1'h0 : _GEN_1179; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1196 = io_slave_out1_sync ? 1'h0 : _GEN_1180; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1197 = io_slave_out1_sync ? 1'h0 : _GEN_1181; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1198 = io_slave_out1_sync ? 1'h0 : _GEN_1182; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1199 = io_slave_out1_sync ? 1'h0 : _GEN_1183; // @[Bus.scala 477:50:@555.8]
  assign _GEN_1200 = _T_440 ? _GEN_1184 : _GEN_1168; // @[Bus.scala 476:41:@554.6]
  assign _GEN_1201 = _T_440 ? $signed(_GEN_1185) : $signed(_GEN_1169); // @[Bus.scala 476:41:@554.6]
  assign _GEN_1202 = _T_440 ? $signed(_GEN_1186) : $signed(_GEN_1170); // @[Bus.scala 476:41:@554.6]
  assign _GEN_1203 = _T_440 ? _GEN_1187 : _GEN_1171; // @[Bus.scala 476:41:@554.6]
  assign _GEN_1204 = _T_440 ? _GEN_1188 : _GEN_1172; // @[Bus.scala 476:41:@554.6]
  assign _GEN_1205 = _T_440 ? $signed(_GEN_1189) : $signed(_GEN_1173); // @[Bus.scala 476:41:@554.6]
  assign _GEN_1206 = _T_440 ? _GEN_1190 : _GEN_1174; // @[Bus.scala 476:41:@554.6]
  assign _GEN_1207 = _T_440 ? _GEN_1191 : _GEN_1175; // @[Bus.scala 476:41:@554.6]
  assign _GEN_1208 = _T_440 ? _GEN_1192 : _GEN_1176; // @[Bus.scala 476:41:@554.6]
  assign _GEN_1209 = _T_440 ? _GEN_1193 : _GEN_1177; // @[Bus.scala 476:41:@554.6]
  assign _GEN_1210 = _T_440 ? _GEN_1194 : _GEN_1178; // @[Bus.scala 476:41:@554.6]
  assign _GEN_1211 = _T_440 ? _GEN_1195 : _GEN_1179; // @[Bus.scala 476:41:@554.6]
  assign _GEN_1212 = _T_440 ? _GEN_1196 : _GEN_1180; // @[Bus.scala 476:41:@554.6]
  assign _GEN_1213 = _T_440 ? _GEN_1197 : _GEN_1181; // @[Bus.scala 476:41:@554.6]
  assign _GEN_1214 = _T_440 ? _GEN_1198 : _GEN_1182; // @[Bus.scala 476:41:@554.6]
  assign _GEN_1215 = _T_440 ? _GEN_1199 : _GEN_1183; // @[Bus.scala 476:41:@554.6]
  assign _T_451 = state_r == 4'h5; // @[Bus.scala 496:30:@574.6]
  assign _GEN_1216 = io_slave_in1_sync ? 4'h3 : _GEN_1200; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1217 = io_slave_in1_sync ? io_slave_in1_ack : _GEN_1135; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1218 = io_slave_in1_sync ? $signed(io_slave_in1_data) : $signed(_GEN_1136); // @[Bus.scala 498:57:@579.10]
  assign _GEN_1219 = io_slave_in1_sync ? $signed(req_signal_r_addr) : $signed(_GEN_1201); // @[Bus.scala 498:57:@579.10]
  assign _GEN_1220 = io_slave_in1_sync ? $signed(req_signal_r_data) : $signed(_GEN_1202); // @[Bus.scala 498:57:@579.10]
  assign _GEN_1221 = io_slave_in1_sync ? req_signal_r_trans_type : _GEN_1203; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1222 = io_slave_in1_sync ? io_slave_in1_ack : _GEN_1204; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1223 = io_slave_in1_sync ? $signed(io_slave_in1_data) : $signed(_GEN_1205); // @[Bus.scala 498:57:@579.10]
  assign _GEN_1224 = io_slave_in1_sync ? 1'h0 : _GEN_1206; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1225 = io_slave_in1_sync ? 1'h1 : _GEN_1207; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1226 = io_slave_in1_sync ? 1'h0 : _GEN_1208; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1227 = io_slave_in1_sync ? 1'h0 : _GEN_1209; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1228 = io_slave_in1_sync ? 1'h0 : _GEN_1210; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1229 = io_slave_in1_sync ? 1'h0 : _GEN_1211; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1230 = io_slave_in1_sync ? 1'h0 : _GEN_1212; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1231 = io_slave_in1_sync ? 1'h0 : _GEN_1213; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1232 = io_slave_in1_sync ? 1'h0 : _GEN_1214; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1233 = io_slave_in1_sync ? 1'h0 : _GEN_1215; // @[Bus.scala 498:57:@579.10]
  assign _GEN_1234 = _T_404 ? _GEN_1216 : _GEN_1200; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1235 = _T_404 ? _GEN_1217 : _GEN_1135; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1236 = _T_404 ? $signed(_GEN_1218) : $signed(_GEN_1136); // @[Bus.scala 497:75:@578.8]
  assign _GEN_1237 = _T_404 ? $signed(_GEN_1219) : $signed(_GEN_1201); // @[Bus.scala 497:75:@578.8]
  assign _GEN_1238 = _T_404 ? $signed(_GEN_1220) : $signed(_GEN_1202); // @[Bus.scala 497:75:@578.8]
  assign _GEN_1239 = _T_404 ? _GEN_1221 : _GEN_1203; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1240 = _T_404 ? _GEN_1222 : _GEN_1204; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1241 = _T_404 ? $signed(_GEN_1223) : $signed(_GEN_1205); // @[Bus.scala 497:75:@578.8]
  assign _GEN_1242 = _T_404 ? _GEN_1224 : _GEN_1206; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1243 = _T_404 ? _GEN_1225 : _GEN_1207; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1244 = _T_404 ? _GEN_1226 : _GEN_1208; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1245 = _T_404 ? _GEN_1227 : _GEN_1209; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1246 = _T_404 ? _GEN_1228 : _GEN_1210; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1247 = _T_404 ? _GEN_1229 : _GEN_1211; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1248 = _T_404 ? _GEN_1230 : _GEN_1212; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1249 = _T_404 ? _GEN_1231 : _GEN_1213; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1250 = _T_404 ? _GEN_1232 : _GEN_1214; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1251 = _T_404 ? _GEN_1233 : _GEN_1215; // @[Bus.scala 497:75:@578.8]
  assign _GEN_1252 = _T_451 ? _GEN_1234 : _GEN_1200; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1253 = _T_451 ? _GEN_1235 : _GEN_1135; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1254 = _T_451 ? $signed(_GEN_1236) : $signed(_GEN_1136); // @[Bus.scala 496:41:@575.6]
  assign _GEN_1255 = _T_451 ? $signed(_GEN_1237) : $signed(_GEN_1201); // @[Bus.scala 496:41:@575.6]
  assign _GEN_1256 = _T_451 ? $signed(_GEN_1238) : $signed(_GEN_1202); // @[Bus.scala 496:41:@575.6]
  assign _GEN_1257 = _T_451 ? _GEN_1239 : _GEN_1203; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1258 = _T_451 ? _GEN_1240 : _GEN_1204; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1259 = _T_451 ? $signed(_GEN_1241) : $signed(_GEN_1205); // @[Bus.scala 496:41:@575.6]
  assign _GEN_1260 = _T_451 ? _GEN_1242 : _GEN_1206; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1261 = _T_451 ? _GEN_1243 : _GEN_1207; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1262 = _T_451 ? _GEN_1244 : _GEN_1208; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1263 = _T_451 ? _GEN_1245 : _GEN_1209; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1264 = _T_451 ? _GEN_1246 : _GEN_1210; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1265 = _T_451 ? _GEN_1247 : _GEN_1211; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1266 = _T_451 ? _GEN_1248 : _GEN_1212; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1267 = _T_451 ? _GEN_1249 : _GEN_1213; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1268 = _T_451 ? _GEN_1250 : _GEN_1214; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1269 = _T_451 ? _GEN_1251 : _GEN_1215; // @[Bus.scala 496:41:@575.6]
  assign _GEN_1270 = io_slave_in1_sync ? 4'h3 : _GEN_1252; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1271 = io_slave_in1_sync ? io_slave_in1_ack : _GEN_1253; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1272 = io_slave_in1_sync ? $signed(32'sh0) : $signed(_GEN_1254); // @[Bus.scala 522:57:@605.10]
  assign _GEN_1273 = io_slave_in1_sync ? $signed(req_signal_r_addr) : $signed(_GEN_1255); // @[Bus.scala 522:57:@605.10]
  assign _GEN_1274 = io_slave_in1_sync ? $signed(req_signal_r_data) : $signed(_GEN_1256); // @[Bus.scala 522:57:@605.10]
  assign _GEN_1275 = io_slave_in1_sync ? req_signal_r_trans_type : _GEN_1257; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1276 = io_slave_in1_sync ? io_slave_in1_ack : _GEN_1258; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1277 = io_slave_in1_sync ? $signed(32'sh0) : $signed(_GEN_1259); // @[Bus.scala 522:57:@605.10]
  assign _GEN_1278 = io_slave_in1_sync ? 1'h0 : _GEN_1260; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1279 = io_slave_in1_sync ? 1'h1 : _GEN_1261; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1280 = io_slave_in1_sync ? 1'h0 : _GEN_1262; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1281 = io_slave_in1_sync ? 1'h0 : _GEN_1263; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1282 = io_slave_in1_sync ? 1'h0 : _GEN_1264; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1283 = io_slave_in1_sync ? 1'h0 : _GEN_1265; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1284 = io_slave_in1_sync ? 1'h0 : _GEN_1266; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1285 = io_slave_in1_sync ? 1'h0 : _GEN_1267; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1286 = io_slave_in1_sync ? 1'h0 : _GEN_1268; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1287 = io_slave_in1_sync ? 1'h0 : _GEN_1269; // @[Bus.scala 522:57:@605.10]
  assign _GEN_1288 = _T_402 ? _GEN_1270 : _GEN_1252; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1289 = _T_402 ? _GEN_1271 : _GEN_1253; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1290 = _T_402 ? $signed(_GEN_1272) : $signed(_GEN_1254); // @[Bus.scala 521:74:@604.8]
  assign _GEN_1291 = _T_402 ? $signed(_GEN_1273) : $signed(_GEN_1255); // @[Bus.scala 521:74:@604.8]
  assign _GEN_1292 = _T_402 ? $signed(_GEN_1274) : $signed(_GEN_1256); // @[Bus.scala 521:74:@604.8]
  assign _GEN_1293 = _T_402 ? _GEN_1275 : _GEN_1257; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1294 = _T_402 ? _GEN_1276 : _GEN_1258; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1295 = _T_402 ? $signed(_GEN_1277) : $signed(_GEN_1259); // @[Bus.scala 521:74:@604.8]
  assign _GEN_1296 = _T_402 ? _GEN_1278 : _GEN_1260; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1297 = _T_402 ? _GEN_1279 : _GEN_1261; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1298 = _T_402 ? _GEN_1280 : _GEN_1262; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1299 = _T_402 ? _GEN_1281 : _GEN_1263; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1300 = _T_402 ? _GEN_1282 : _GEN_1264; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1301 = _T_402 ? _GEN_1283 : _GEN_1265; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1302 = _T_402 ? _GEN_1284 : _GEN_1266; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1303 = _T_402 ? _GEN_1285 : _GEN_1267; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1304 = _T_402 ? _GEN_1286 : _GEN_1268; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1305 = _T_402 ? _GEN_1287 : _GEN_1269; // @[Bus.scala 521:74:@604.8]
  assign _GEN_1306 = _T_451 ? _GEN_1288 : _GEN_1252; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1307 = _T_451 ? _GEN_1289 : _GEN_1253; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1308 = _T_451 ? $signed(_GEN_1290) : $signed(_GEN_1254); // @[Bus.scala 520:41:@602.6]
  assign _GEN_1309 = _T_451 ? $signed(_GEN_1291) : $signed(_GEN_1255); // @[Bus.scala 520:41:@602.6]
  assign _GEN_1310 = _T_451 ? $signed(_GEN_1292) : $signed(_GEN_1256); // @[Bus.scala 520:41:@602.6]
  assign _GEN_1311 = _T_451 ? _GEN_1293 : _GEN_1257; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1312 = _T_451 ? _GEN_1294 : _GEN_1258; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1313 = _T_451 ? $signed(_GEN_1295) : $signed(_GEN_1259); // @[Bus.scala 520:41:@602.6]
  assign _GEN_1314 = _T_451 ? _GEN_1296 : _GEN_1260; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1315 = _T_451 ? _GEN_1297 : _GEN_1261; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1316 = _T_451 ? _GEN_1298 : _GEN_1262; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1317 = _T_451 ? _GEN_1299 : _GEN_1263; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1318 = _T_451 ? _GEN_1300 : _GEN_1264; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1319 = _T_451 ? _GEN_1301 : _GEN_1265; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1320 = _T_451 ? _GEN_1302 : _GEN_1266; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1321 = _T_451 ? _GEN_1303 : _GEN_1267; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1322 = _T_451 ? _GEN_1304 : _GEN_1268; // @[Bus.scala 520:41:@602.6]
  assign _GEN_1323 = _T_451 ? _GEN_1305 : _GEN_1269; // @[Bus.scala 520:41:@602.6]
  assign _T_479 = state_r == 4'h6; // @[Bus.scala 544:30:@627.6]
  assign _GEN_1324 = io_slave_out2_sync ? 4'h7 : _GEN_1306; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1325 = io_slave_out2_sync ? $signed(req_signal_r_addr) : $signed(_GEN_1309); // @[Bus.scala 545:50:@629.8]
  assign _GEN_1326 = io_slave_out2_sync ? $signed(req_signal_r_data) : $signed(_GEN_1310); // @[Bus.scala 545:50:@629.8]
  assign _GEN_1327 = io_slave_out2_sync ? req_signal_r_trans_type : _GEN_1311; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1328 = io_slave_out2_sync ? resp_signal_r_ack : _GEN_1312; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1329 = io_slave_out2_sync ? $signed(resp_signal_r_data) : $signed(_GEN_1313); // @[Bus.scala 545:50:@629.8]
  assign _GEN_1330 = io_slave_out2_sync ? 1'h0 : _GEN_1314; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1331 = io_slave_out2_sync ? 1'h0 : _GEN_1315; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1332 = io_slave_out2_sync ? 1'h0 : _GEN_1316; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1333 = io_slave_out2_sync ? 1'h0 : _GEN_1317; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1334 = io_slave_out2_sync ? 1'h1 : _GEN_1318; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1335 = io_slave_out2_sync ? 1'h0 : _GEN_1319; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1336 = io_slave_out2_sync ? 1'h0 : _GEN_1320; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1337 = io_slave_out2_sync ? 1'h0 : _GEN_1321; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1338 = io_slave_out2_sync ? 1'h0 : _GEN_1322; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1339 = io_slave_out2_sync ? 1'h0 : _GEN_1323; // @[Bus.scala 545:50:@629.8]
  assign _GEN_1340 = _T_479 ? _GEN_1324 : _GEN_1306; // @[Bus.scala 544:41:@628.6]
  assign _GEN_1341 = _T_479 ? $signed(_GEN_1325) : $signed(_GEN_1309); // @[Bus.scala 544:41:@628.6]
  assign _GEN_1342 = _T_479 ? $signed(_GEN_1326) : $signed(_GEN_1310); // @[Bus.scala 544:41:@628.6]
  assign _GEN_1343 = _T_479 ? _GEN_1327 : _GEN_1311; // @[Bus.scala 544:41:@628.6]
  assign _GEN_1344 = _T_479 ? _GEN_1328 : _GEN_1312; // @[Bus.scala 544:41:@628.6]
  assign _GEN_1345 = _T_479 ? $signed(_GEN_1329) : $signed(_GEN_1313); // @[Bus.scala 544:41:@628.6]
  assign _GEN_1346 = _T_479 ? _GEN_1330 : _GEN_1314; // @[Bus.scala 544:41:@628.6]
  assign _GEN_1347 = _T_479 ? _GEN_1331 : _GEN_1315; // @[Bus.scala 544:41:@628.6]
  assign _GEN_1348 = _T_479 ? _GEN_1332 : _GEN_1316; // @[Bus.scala 544:41:@628.6]
  assign _GEN_1349 = _T_479 ? _GEN_1333 : _GEN_1317; // @[Bus.scala 544:41:@628.6]
  assign _GEN_1350 = _T_479 ? _GEN_1334 : _GEN_1318; // @[Bus.scala 544:41:@628.6]
  assign _GEN_1351 = _T_479 ? _GEN_1335 : _GEN_1319; // @[Bus.scala 544:41:@628.6]
  assign _GEN_1352 = _T_479 ? _GEN_1336 : _GEN_1320; // @[Bus.scala 544:41:@628.6]
  assign _GEN_1353 = _T_479 ? _GEN_1337 : _GEN_1321; // @[Bus.scala 544:41:@628.6]
  assign _GEN_1354 = _T_479 ? _GEN_1338 : _GEN_1322; // @[Bus.scala 544:41:@628.6]
  assign _GEN_1355 = _T_479 ? _GEN_1339 : _GEN_1323; // @[Bus.scala 544:41:@628.6]
  assign _T_490 = state_r == 4'h7; // @[Bus.scala 564:30:@648.6]
  assign _GEN_1356 = io_slave_in2_sync ? 4'h3 : _GEN_1340; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1357 = io_slave_in2_sync ? io_slave_in2_ack : _GEN_1307; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1358 = io_slave_in2_sync ? $signed(io_slave_in2_data) : $signed(_GEN_1308); // @[Bus.scala 566:57:@653.10]
  assign _GEN_1359 = io_slave_in2_sync ? $signed(req_signal_r_addr) : $signed(_GEN_1341); // @[Bus.scala 566:57:@653.10]
  assign _GEN_1360 = io_slave_in2_sync ? $signed(req_signal_r_data) : $signed(_GEN_1342); // @[Bus.scala 566:57:@653.10]
  assign _GEN_1361 = io_slave_in2_sync ? req_signal_r_trans_type : _GEN_1343; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1362 = io_slave_in2_sync ? io_slave_in2_ack : _GEN_1344; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1363 = io_slave_in2_sync ? $signed(io_slave_in2_data) : $signed(_GEN_1345); // @[Bus.scala 566:57:@653.10]
  assign _GEN_1364 = io_slave_in2_sync ? 1'h0 : _GEN_1346; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1365 = io_slave_in2_sync ? 1'h1 : _GEN_1347; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1366 = io_slave_in2_sync ? 1'h0 : _GEN_1348; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1367 = io_slave_in2_sync ? 1'h0 : _GEN_1349; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1368 = io_slave_in2_sync ? 1'h0 : _GEN_1350; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1369 = io_slave_in2_sync ? 1'h0 : _GEN_1351; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1370 = io_slave_in2_sync ? 1'h0 : _GEN_1352; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1371 = io_slave_in2_sync ? 1'h0 : _GEN_1353; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1372 = io_slave_in2_sync ? 1'h0 : _GEN_1354; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1373 = io_slave_in2_sync ? 1'h0 : _GEN_1355; // @[Bus.scala 566:57:@653.10]
  assign _GEN_1374 = _T_404 ? _GEN_1356 : _GEN_1340; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1375 = _T_404 ? _GEN_1357 : _GEN_1307; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1376 = _T_404 ? $signed(_GEN_1358) : $signed(_GEN_1308); // @[Bus.scala 565:75:@652.8]
  assign _GEN_1377 = _T_404 ? $signed(_GEN_1359) : $signed(_GEN_1341); // @[Bus.scala 565:75:@652.8]
  assign _GEN_1378 = _T_404 ? $signed(_GEN_1360) : $signed(_GEN_1342); // @[Bus.scala 565:75:@652.8]
  assign _GEN_1379 = _T_404 ? _GEN_1361 : _GEN_1343; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1380 = _T_404 ? _GEN_1362 : _GEN_1344; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1381 = _T_404 ? $signed(_GEN_1363) : $signed(_GEN_1345); // @[Bus.scala 565:75:@652.8]
  assign _GEN_1382 = _T_404 ? _GEN_1364 : _GEN_1346; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1383 = _T_404 ? _GEN_1365 : _GEN_1347; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1384 = _T_404 ? _GEN_1366 : _GEN_1348; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1385 = _T_404 ? _GEN_1367 : _GEN_1349; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1386 = _T_404 ? _GEN_1368 : _GEN_1350; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1387 = _T_404 ? _GEN_1369 : _GEN_1351; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1388 = _T_404 ? _GEN_1370 : _GEN_1352; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1389 = _T_404 ? _GEN_1371 : _GEN_1353; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1390 = _T_404 ? _GEN_1372 : _GEN_1354; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1391 = _T_404 ? _GEN_1373 : _GEN_1355; // @[Bus.scala 565:75:@652.8]
  assign _GEN_1392 = _T_490 ? _GEN_1374 : _GEN_1340; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1393 = _T_490 ? _GEN_1375 : _GEN_1307; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1394 = _T_490 ? $signed(_GEN_1376) : $signed(_GEN_1308); // @[Bus.scala 564:41:@649.6]
  assign _GEN_1395 = _T_490 ? $signed(_GEN_1377) : $signed(_GEN_1341); // @[Bus.scala 564:41:@649.6]
  assign _GEN_1396 = _T_490 ? $signed(_GEN_1378) : $signed(_GEN_1342); // @[Bus.scala 564:41:@649.6]
  assign _GEN_1397 = _T_490 ? _GEN_1379 : _GEN_1343; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1398 = _T_490 ? _GEN_1380 : _GEN_1344; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1399 = _T_490 ? $signed(_GEN_1381) : $signed(_GEN_1345); // @[Bus.scala 564:41:@649.6]
  assign _GEN_1400 = _T_490 ? _GEN_1382 : _GEN_1346; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1401 = _T_490 ? _GEN_1383 : _GEN_1347; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1402 = _T_490 ? _GEN_1384 : _GEN_1348; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1403 = _T_490 ? _GEN_1385 : _GEN_1349; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1404 = _T_490 ? _GEN_1386 : _GEN_1350; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1405 = _T_490 ? _GEN_1387 : _GEN_1351; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1406 = _T_490 ? _GEN_1388 : _GEN_1352; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1407 = _T_490 ? _GEN_1389 : _GEN_1353; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1408 = _T_490 ? _GEN_1390 : _GEN_1354; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1409 = _T_490 ? _GEN_1391 : _GEN_1355; // @[Bus.scala 564:41:@649.6]
  assign _GEN_1410 = io_slave_in2_sync ? 4'h3 : _GEN_1392; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1411 = io_slave_in2_sync ? io_slave_in2_ack : _GEN_1393; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1412 = io_slave_in2_sync ? $signed(32'sh0) : $signed(_GEN_1394); // @[Bus.scala 590:57:@679.10]
  assign _GEN_1413 = io_slave_in2_sync ? $signed(req_signal_r_addr) : $signed(_GEN_1395); // @[Bus.scala 590:57:@679.10]
  assign _GEN_1414 = io_slave_in2_sync ? $signed(req_signal_r_data) : $signed(_GEN_1396); // @[Bus.scala 590:57:@679.10]
  assign _GEN_1415 = io_slave_in2_sync ? req_signal_r_trans_type : _GEN_1397; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1416 = io_slave_in2_sync ? io_slave_in2_ack : _GEN_1398; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1417 = io_slave_in2_sync ? $signed(32'sh0) : $signed(_GEN_1399); // @[Bus.scala 590:57:@679.10]
  assign _GEN_1418 = io_slave_in2_sync ? 1'h0 : _GEN_1400; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1419 = io_slave_in2_sync ? 1'h1 : _GEN_1401; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1420 = io_slave_in2_sync ? 1'h0 : _GEN_1402; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1421 = io_slave_in2_sync ? 1'h0 : _GEN_1403; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1422 = io_slave_in2_sync ? 1'h0 : _GEN_1404; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1423 = io_slave_in2_sync ? 1'h0 : _GEN_1405; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1424 = io_slave_in2_sync ? 1'h0 : _GEN_1406; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1425 = io_slave_in2_sync ? 1'h0 : _GEN_1407; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1426 = io_slave_in2_sync ? 1'h0 : _GEN_1408; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1427 = io_slave_in2_sync ? 1'h0 : _GEN_1409; // @[Bus.scala 590:57:@679.10]
  assign _GEN_1428 = _T_402 ? _GEN_1410 : _GEN_1392; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1429 = _T_402 ? _GEN_1411 : _GEN_1393; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1430 = _T_402 ? $signed(_GEN_1412) : $signed(_GEN_1394); // @[Bus.scala 589:74:@678.8]
  assign _GEN_1431 = _T_402 ? $signed(_GEN_1413) : $signed(_GEN_1395); // @[Bus.scala 589:74:@678.8]
  assign _GEN_1432 = _T_402 ? $signed(_GEN_1414) : $signed(_GEN_1396); // @[Bus.scala 589:74:@678.8]
  assign _GEN_1433 = _T_402 ? _GEN_1415 : _GEN_1397; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1434 = _T_402 ? _GEN_1416 : _GEN_1398; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1435 = _T_402 ? $signed(_GEN_1417) : $signed(_GEN_1399); // @[Bus.scala 589:74:@678.8]
  assign _GEN_1436 = _T_402 ? _GEN_1418 : _GEN_1400; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1437 = _T_402 ? _GEN_1419 : _GEN_1401; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1438 = _T_402 ? _GEN_1420 : _GEN_1402; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1439 = _T_402 ? _GEN_1421 : _GEN_1403; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1440 = _T_402 ? _GEN_1422 : _GEN_1404; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1441 = _T_402 ? _GEN_1423 : _GEN_1405; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1442 = _T_402 ? _GEN_1424 : _GEN_1406; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1443 = _T_402 ? _GEN_1425 : _GEN_1407; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1444 = _T_402 ? _GEN_1426 : _GEN_1408; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1445 = _T_402 ? _GEN_1427 : _GEN_1409; // @[Bus.scala 589:74:@678.8]
  assign _GEN_1446 = _T_490 ? _GEN_1428 : _GEN_1392; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1447 = _T_490 ? _GEN_1429 : _GEN_1393; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1448 = _T_490 ? $signed(_GEN_1430) : $signed(_GEN_1394); // @[Bus.scala 588:41:@676.6]
  assign _GEN_1449 = _T_490 ? $signed(_GEN_1431) : $signed(_GEN_1395); // @[Bus.scala 588:41:@676.6]
  assign _GEN_1450 = _T_490 ? $signed(_GEN_1432) : $signed(_GEN_1396); // @[Bus.scala 588:41:@676.6]
  assign _GEN_1451 = _T_490 ? _GEN_1433 : _GEN_1397; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1452 = _T_490 ? _GEN_1434 : _GEN_1398; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1453 = _T_490 ? $signed(_GEN_1435) : $signed(_GEN_1399); // @[Bus.scala 588:41:@676.6]
  assign _GEN_1454 = _T_490 ? _GEN_1436 : _GEN_1400; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1455 = _T_490 ? _GEN_1437 : _GEN_1401; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1456 = _T_490 ? _GEN_1438 : _GEN_1402; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1457 = _T_490 ? _GEN_1439 : _GEN_1403; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1458 = _T_490 ? _GEN_1440 : _GEN_1404; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1459 = _T_490 ? _GEN_1441 : _GEN_1405; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1460 = _T_490 ? _GEN_1442 : _GEN_1406; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1461 = _T_490 ? _GEN_1443 : _GEN_1407; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1462 = _T_490 ? _GEN_1444 : _GEN_1408; // @[Bus.scala 588:41:@676.6]
  assign _GEN_1463 = _T_490 ? _GEN_1445 : _GEN_1409; // @[Bus.scala 588:41:@676.6]
  assign _T_518 = state_r == 4'h8; // @[Bus.scala 612:30:@701.6]
  assign _GEN_1464 = io_slave_out3_sync ? 4'h9 : _GEN_1446; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1465 = io_slave_out3_sync ? $signed(req_signal_r_addr) : $signed(_GEN_1449); // @[Bus.scala 613:50:@703.8]
  assign _GEN_1466 = io_slave_out3_sync ? $signed(req_signal_r_data) : $signed(_GEN_1450); // @[Bus.scala 613:50:@703.8]
  assign _GEN_1467 = io_slave_out3_sync ? req_signal_r_trans_type : _GEN_1451; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1468 = io_slave_out3_sync ? resp_signal_r_ack : _GEN_1452; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1469 = io_slave_out3_sync ? $signed(resp_signal_r_data) : $signed(_GEN_1453); // @[Bus.scala 613:50:@703.8]
  assign _GEN_1470 = io_slave_out3_sync ? 1'h0 : _GEN_1454; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1471 = io_slave_out3_sync ? 1'h0 : _GEN_1455; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1472 = io_slave_out3_sync ? 1'h0 : _GEN_1456; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1473 = io_slave_out3_sync ? 1'h0 : _GEN_1457; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1474 = io_slave_out3_sync ? 1'h0 : _GEN_1458; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1475 = io_slave_out3_sync ? 1'h1 : _GEN_1459; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1476 = io_slave_out3_sync ? 1'h0 : _GEN_1460; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1477 = io_slave_out3_sync ? 1'h0 : _GEN_1461; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1478 = io_slave_out3_sync ? 1'h0 : _GEN_1462; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1479 = io_slave_out3_sync ? 1'h0 : _GEN_1463; // @[Bus.scala 613:50:@703.8]
  assign _GEN_1480 = _T_518 ? _GEN_1464 : _GEN_1446; // @[Bus.scala 612:41:@702.6]
  assign _GEN_1481 = _T_518 ? $signed(_GEN_1465) : $signed(_GEN_1449); // @[Bus.scala 612:41:@702.6]
  assign _GEN_1482 = _T_518 ? $signed(_GEN_1466) : $signed(_GEN_1450); // @[Bus.scala 612:41:@702.6]
  assign _GEN_1483 = _T_518 ? _GEN_1467 : _GEN_1451; // @[Bus.scala 612:41:@702.6]
  assign _GEN_1484 = _T_518 ? _GEN_1468 : _GEN_1452; // @[Bus.scala 612:41:@702.6]
  assign _GEN_1485 = _T_518 ? $signed(_GEN_1469) : $signed(_GEN_1453); // @[Bus.scala 612:41:@702.6]
  assign _GEN_1486 = _T_518 ? _GEN_1470 : _GEN_1454; // @[Bus.scala 612:41:@702.6]
  assign _GEN_1487 = _T_518 ? _GEN_1471 : _GEN_1455; // @[Bus.scala 612:41:@702.6]
  assign _GEN_1488 = _T_518 ? _GEN_1472 : _GEN_1456; // @[Bus.scala 612:41:@702.6]
  assign _GEN_1489 = _T_518 ? _GEN_1473 : _GEN_1457; // @[Bus.scala 612:41:@702.6]
  assign _GEN_1490 = _T_518 ? _GEN_1474 : _GEN_1458; // @[Bus.scala 612:41:@702.6]
  assign _GEN_1491 = _T_518 ? _GEN_1475 : _GEN_1459; // @[Bus.scala 612:41:@702.6]
  assign _GEN_1492 = _T_518 ? _GEN_1476 : _GEN_1460; // @[Bus.scala 612:41:@702.6]
  assign _GEN_1493 = _T_518 ? _GEN_1477 : _GEN_1461; // @[Bus.scala 612:41:@702.6]
  assign _GEN_1494 = _T_518 ? _GEN_1478 : _GEN_1462; // @[Bus.scala 612:41:@702.6]
  assign _GEN_1495 = _T_518 ? _GEN_1479 : _GEN_1463; // @[Bus.scala 612:41:@702.6]
  assign _T_529 = state_r == 4'h9; // @[Bus.scala 632:30:@722.6]
  assign _GEN_1496 = io_slave_in3_sync ? 4'h3 : _GEN_1480; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1497 = io_slave_in3_sync ? io_slave_in3_ack : _GEN_1447; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1498 = io_slave_in3_sync ? $signed(io_slave_in3_data) : $signed(_GEN_1448); // @[Bus.scala 634:57:@727.10]
  assign _GEN_1499 = io_slave_in3_sync ? $signed(req_signal_r_addr) : $signed(_GEN_1481); // @[Bus.scala 634:57:@727.10]
  assign _GEN_1500 = io_slave_in3_sync ? $signed(req_signal_r_data) : $signed(_GEN_1482); // @[Bus.scala 634:57:@727.10]
  assign _GEN_1501 = io_slave_in3_sync ? req_signal_r_trans_type : _GEN_1483; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1502 = io_slave_in3_sync ? io_slave_in3_ack : _GEN_1484; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1503 = io_slave_in3_sync ? $signed(io_slave_in3_data) : $signed(_GEN_1485); // @[Bus.scala 634:57:@727.10]
  assign _GEN_1504 = io_slave_in3_sync ? 1'h0 : _GEN_1486; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1505 = io_slave_in3_sync ? 1'h1 : _GEN_1487; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1506 = io_slave_in3_sync ? 1'h0 : _GEN_1488; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1507 = io_slave_in3_sync ? 1'h0 : _GEN_1489; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1508 = io_slave_in3_sync ? 1'h0 : _GEN_1490; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1509 = io_slave_in3_sync ? 1'h0 : _GEN_1491; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1510 = io_slave_in3_sync ? 1'h0 : _GEN_1492; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1511 = io_slave_in3_sync ? 1'h0 : _GEN_1493; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1512 = io_slave_in3_sync ? 1'h0 : _GEN_1494; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1513 = io_slave_in3_sync ? 1'h0 : _GEN_1495; // @[Bus.scala 634:57:@727.10]
  assign _GEN_1514 = _T_404 ? _GEN_1496 : _GEN_1480; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1515 = _T_404 ? _GEN_1497 : _GEN_1447; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1516 = _T_404 ? $signed(_GEN_1498) : $signed(_GEN_1448); // @[Bus.scala 633:75:@726.8]
  assign _GEN_1517 = _T_404 ? $signed(_GEN_1499) : $signed(_GEN_1481); // @[Bus.scala 633:75:@726.8]
  assign _GEN_1518 = _T_404 ? $signed(_GEN_1500) : $signed(_GEN_1482); // @[Bus.scala 633:75:@726.8]
  assign _GEN_1519 = _T_404 ? _GEN_1501 : _GEN_1483; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1520 = _T_404 ? _GEN_1502 : _GEN_1484; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1521 = _T_404 ? $signed(_GEN_1503) : $signed(_GEN_1485); // @[Bus.scala 633:75:@726.8]
  assign _GEN_1522 = _T_404 ? _GEN_1504 : _GEN_1486; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1523 = _T_404 ? _GEN_1505 : _GEN_1487; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1524 = _T_404 ? _GEN_1506 : _GEN_1488; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1525 = _T_404 ? _GEN_1507 : _GEN_1489; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1526 = _T_404 ? _GEN_1508 : _GEN_1490; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1527 = _T_404 ? _GEN_1509 : _GEN_1491; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1528 = _T_404 ? _GEN_1510 : _GEN_1492; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1529 = _T_404 ? _GEN_1511 : _GEN_1493; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1530 = _T_404 ? _GEN_1512 : _GEN_1494; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1531 = _T_404 ? _GEN_1513 : _GEN_1495; // @[Bus.scala 633:75:@726.8]
  assign _GEN_1532 = _T_529 ? _GEN_1514 : _GEN_1480; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1533 = _T_529 ? _GEN_1515 : _GEN_1447; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1534 = _T_529 ? $signed(_GEN_1516) : $signed(_GEN_1448); // @[Bus.scala 632:41:@723.6]
  assign _GEN_1535 = _T_529 ? $signed(_GEN_1517) : $signed(_GEN_1481); // @[Bus.scala 632:41:@723.6]
  assign _GEN_1536 = _T_529 ? $signed(_GEN_1518) : $signed(_GEN_1482); // @[Bus.scala 632:41:@723.6]
  assign _GEN_1537 = _T_529 ? _GEN_1519 : _GEN_1483; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1538 = _T_529 ? _GEN_1520 : _GEN_1484; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1539 = _T_529 ? $signed(_GEN_1521) : $signed(_GEN_1485); // @[Bus.scala 632:41:@723.6]
  assign _GEN_1540 = _T_529 ? _GEN_1522 : _GEN_1486; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1541 = _T_529 ? _GEN_1523 : _GEN_1487; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1542 = _T_529 ? _GEN_1524 : _GEN_1488; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1543 = _T_529 ? _GEN_1525 : _GEN_1489; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1544 = _T_529 ? _GEN_1526 : _GEN_1490; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1545 = _T_529 ? _GEN_1527 : _GEN_1491; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1546 = _T_529 ? _GEN_1528 : _GEN_1492; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1547 = _T_529 ? _GEN_1529 : _GEN_1493; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1548 = _T_529 ? _GEN_1530 : _GEN_1494; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1549 = _T_529 ? _GEN_1531 : _GEN_1495; // @[Bus.scala 632:41:@723.6]
  assign _GEN_1550 = io_slave_in3_sync ? 4'h3 : _GEN_1532; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1551 = io_slave_in3_sync ? io_slave_in3_ack : _GEN_1533; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1552 = io_slave_in3_sync ? $signed(32'sh0) : $signed(_GEN_1534); // @[Bus.scala 658:57:@753.10]
  assign _GEN_1553 = io_slave_in3_sync ? $signed(req_signal_r_addr) : $signed(_GEN_1535); // @[Bus.scala 658:57:@753.10]
  assign _GEN_1554 = io_slave_in3_sync ? $signed(req_signal_r_data) : $signed(_GEN_1536); // @[Bus.scala 658:57:@753.10]
  assign _GEN_1555 = io_slave_in3_sync ? req_signal_r_trans_type : _GEN_1537; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1556 = io_slave_in3_sync ? io_slave_in3_ack : _GEN_1538; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1557 = io_slave_in3_sync ? $signed(32'sh0) : $signed(_GEN_1539); // @[Bus.scala 658:57:@753.10]
  assign _GEN_1558 = io_slave_in3_sync ? 1'h0 : _GEN_1540; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1559 = io_slave_in3_sync ? 1'h1 : _GEN_1541; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1560 = io_slave_in3_sync ? 1'h0 : _GEN_1542; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1561 = io_slave_in3_sync ? 1'h0 : _GEN_1543; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1562 = io_slave_in3_sync ? 1'h0 : _GEN_1544; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1563 = io_slave_in3_sync ? 1'h0 : _GEN_1545; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1564 = io_slave_in3_sync ? 1'h0 : _GEN_1546; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1565 = io_slave_in3_sync ? 1'h0 : _GEN_1547; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1566 = io_slave_in3_sync ? 1'h0 : _GEN_1548; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1567 = io_slave_in3_sync ? 1'h0 : _GEN_1549; // @[Bus.scala 658:57:@753.10]
  assign _GEN_1568 = _T_402 ? _GEN_1550 : _GEN_1532; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1569 = _T_402 ? _GEN_1551 : _GEN_1533; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1570 = _T_402 ? $signed(_GEN_1552) : $signed(_GEN_1534); // @[Bus.scala 657:74:@752.8]
  assign _GEN_1571 = _T_402 ? $signed(_GEN_1553) : $signed(_GEN_1535); // @[Bus.scala 657:74:@752.8]
  assign _GEN_1572 = _T_402 ? $signed(_GEN_1554) : $signed(_GEN_1536); // @[Bus.scala 657:74:@752.8]
  assign _GEN_1573 = _T_402 ? _GEN_1555 : _GEN_1537; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1574 = _T_402 ? _GEN_1556 : _GEN_1538; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1575 = _T_402 ? $signed(_GEN_1557) : $signed(_GEN_1539); // @[Bus.scala 657:74:@752.8]
  assign _GEN_1576 = _T_402 ? _GEN_1558 : _GEN_1540; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1577 = _T_402 ? _GEN_1559 : _GEN_1541; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1578 = _T_402 ? _GEN_1560 : _GEN_1542; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1579 = _T_402 ? _GEN_1561 : _GEN_1543; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1580 = _T_402 ? _GEN_1562 : _GEN_1544; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1581 = _T_402 ? _GEN_1563 : _GEN_1545; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1582 = _T_402 ? _GEN_1564 : _GEN_1546; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1583 = _T_402 ? _GEN_1565 : _GEN_1547; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1584 = _T_402 ? _GEN_1566 : _GEN_1548; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1585 = _T_402 ? _GEN_1567 : _GEN_1549; // @[Bus.scala 657:74:@752.8]
  assign _GEN_1586 = _T_529 ? _GEN_1568 : _GEN_1532; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1587 = _T_529 ? _GEN_1569 : _GEN_1533; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1588 = _T_529 ? $signed(_GEN_1570) : $signed(_GEN_1534); // @[Bus.scala 656:41:@750.6]
  assign _GEN_1589 = _T_529 ? $signed(_GEN_1571) : $signed(_GEN_1535); // @[Bus.scala 656:41:@750.6]
  assign _GEN_1590 = _T_529 ? $signed(_GEN_1572) : $signed(_GEN_1536); // @[Bus.scala 656:41:@750.6]
  assign _GEN_1591 = _T_529 ? _GEN_1573 : _GEN_1537; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1592 = _T_529 ? _GEN_1574 : _GEN_1538; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1593 = _T_529 ? $signed(_GEN_1575) : $signed(_GEN_1539); // @[Bus.scala 656:41:@750.6]
  assign _GEN_1594 = _T_529 ? _GEN_1576 : _GEN_1540; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1595 = _T_529 ? _GEN_1577 : _GEN_1541; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1596 = _T_529 ? _GEN_1578 : _GEN_1542; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1597 = _T_529 ? _GEN_1579 : _GEN_1543; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1598 = _T_529 ? _GEN_1580 : _GEN_1544; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1599 = _T_529 ? _GEN_1581 : _GEN_1545; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1600 = _T_529 ? _GEN_1582 : _GEN_1546; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1601 = _T_529 ? _GEN_1583 : _GEN_1547; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1602 = _T_529 ? _GEN_1584 : _GEN_1548; // @[Bus.scala 656:41:@750.6]
  assign _GEN_1603 = _T_529 ? _GEN_1585 : _GEN_1549; // @[Bus.scala 656:41:@750.6]
  assign io_master_in_notify = master_in_notify_r; // @[Bus.scala 685:29:@776.4]
  assign io_master_out_notify = master_out_notify_r; // @[Bus.scala 686:30:@777.4]
  assign io_slave_in0_notify = slave_in0_notify_r; // @[Bus.scala 687:29:@778.4]
  assign io_slave_in1_notify = slave_in1_notify_r; // @[Bus.scala 688:29:@779.4]
  assign io_slave_in2_notify = slave_in2_notify_r; // @[Bus.scala 689:29:@780.4]
  assign io_slave_in3_notify = slave_in3_notify_r; // @[Bus.scala 690:29:@781.4]
  assign io_slave_out0_notify = slave_out0_notify_r; // @[Bus.scala 691:30:@782.4]
  assign io_slave_out1_notify = slave_out1_notify_r; // @[Bus.scala 692:30:@783.4]
  assign io_slave_out2_notify = slave_out2_notify_r; // @[Bus.scala 693:30:@784.4]
  assign io_slave_out3_notify = slave_out3_notify_r; // @[Bus.scala 694:30:@785.4]
  assign io_master_out_ack = master_out_r_ack; // @[Bus.scala 695:23:@787.4]
  assign io_master_out_data = master_out_r_data; // @[Bus.scala 695:23:@786.4]
  assign io_slave_out0_addr = slave_out0_r_addr; // @[Bus.scala 696:23:@790.4]
  assign io_slave_out0_data = slave_out0_r_data; // @[Bus.scala 696:23:@789.4]
  assign io_slave_out0_trans_type = slave_out0_r_trans_type; // @[Bus.scala 696:23:@788.4]
  assign io_slave_out1_addr = slave_out1_r_addr; // @[Bus.scala 697:23:@793.4]
  assign io_slave_out1_data = slave_out1_r_data; // @[Bus.scala 697:23:@792.4]
  assign io_slave_out1_trans_type = slave_out1_r_trans_type; // @[Bus.scala 697:23:@791.4]
  assign io_slave_out2_addr = slave_out2_r_addr; // @[Bus.scala 698:23:@796.4]
  assign io_slave_out2_data = slave_out2_r_data; // @[Bus.scala 698:23:@795.4]
  assign io_slave_out2_trans_type = slave_out2_r_trans_type; // @[Bus.scala 698:23:@794.4]
  assign io_slave_out3_addr = slave_out3_r_addr; // @[Bus.scala 699:23:@799.4]
  assign io_slave_out3_data = slave_out3_r_data; // @[Bus.scala 699:23:@798.4]
  assign io_slave_out3_trans_type = slave_out3_r_trans_type; // @[Bus.scala 699:23:@797.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  master_in_notify_r = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  master_out_notify_r = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  slave_in0_notify_r = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  slave_in1_notify_r = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  slave_in2_notify_r = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  slave_in3_notify_r = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  slave_out0_notify_r = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  slave_out1_notify_r = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  slave_out2_notify_r = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  slave_out3_notify_r = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  master_out_r_ack = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  master_out_r_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  slave_out0_r_addr = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  slave_out0_r_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  slave_out0_r_trans_type = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  slave_out1_r_addr = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  slave_out1_r_data = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  slave_out1_r_trans_type = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  slave_out2_r_addr = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  slave_out2_r_data = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  slave_out2_r_trans_type = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  slave_out3_r_addr = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  slave_out3_r_data = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  slave_out3_r_trans_type = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  req_signal_r_addr = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  req_signal_r_data = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  req_signal_r_trans_type = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  resp_signal_r_ack = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  resp_signal_r_data = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  state_r = _RAND_29[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      master_in_notify_r <= 1'h1;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            master_in_notify_r <= 1'h0;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  master_in_notify_r <= 1'h0;
                end else begin
                  if (_T_518) begin
                    if (io_slave_out3_sync) begin
                      master_in_notify_r <= 1'h0;
                    end else begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            master_in_notify_r <= 1'h0;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  master_in_notify_r <= 1'h0;
                                end else begin
                                  if (_T_479) begin
                                    if (io_slave_out2_sync) begin
                                      master_in_notify_r <= 1'h0;
                                    end else begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            master_in_notify_r <= 1'h0;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  master_in_notify_r <= 1'h0;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (io_slave_out1_sync) begin
                                                      master_in_notify_r <= 1'h0;
                                                    end else begin
                                                      if (_T_429) begin
                                                        if (io_master_out_sync) begin
                                                          master_in_notify_r <= 1'h1;
                                                        end else begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                master_in_notify_r <= 1'h0;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      master_in_notify_r <= 1'h0;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (io_slave_out0_sync) begin
                                                                          master_in_notify_r <= 1'h0;
                                                                        end else begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    master_in_notify_r <= 1'h0;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              master_in_notify_r <= 1'h0;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        master_in_notify_r <= 1'h0;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  master_in_notify_r <= 1'h0;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            master_in_notify_r <= 1'h0;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      master_in_notify_r <= 1'h0;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    master_in_notify_r <= 1'h0;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  master_in_notify_r <= 1'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            master_in_notify_r <= 1'h0;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      master_in_notify_r <= 1'h0;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    master_in_notify_r <= 1'h0;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  master_in_notify_r <= 1'h0;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                master_in_notify_r <= 1'h0;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    master_in_notify_r <= _GEN_85;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          master_in_notify_r <= 1'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                          master_in_notify_r <= _GEN_85;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        master_in_notify_r <= _GEN_85;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      master_in_notify_r <= _GEN_85;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    master_in_notify_r <= _GEN_85;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  master_in_notify_r <= _GEN_85;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        master_in_notify_r <= 1'h0;
                                                                                                                                                                      end else begin
                                                                                                                                                                        master_in_notify_r <= _GEN_85;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      master_in_notify_r <= _GEN_85;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    master_in_notify_r <= _GEN_85;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  master_in_notify_r <= _GEN_85;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                master_in_notify_r <= _GEN_85;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      master_in_notify_r <= 1'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                      master_in_notify_r <= _GEN_85;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    master_in_notify_r <= _GEN_85;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  master_in_notify_r <= _GEN_85;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                master_in_notify_r <= _GEN_85;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              master_in_notify_r <= _GEN_85;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          master_in_notify_r <= _GEN_180;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        master_in_notify_r <= _GEN_180;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      master_in_notify_r <= _GEN_180;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                master_in_notify_r <= 1'h0;
                                                                                                                                                              end else begin
                                                                                                                                                                master_in_notify_r <= _GEN_180;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              master_in_notify_r <= _GEN_180;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            master_in_notify_r <= _GEN_180;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          master_in_notify_r <= _GEN_180;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        master_in_notify_r <= _GEN_180;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      master_in_notify_r <= _GEN_180;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    master_in_notify_r <= _GEN_180;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              master_in_notify_r <= 1'h0;
                                                                                                                                                            end else begin
                                                                                                                                                              master_in_notify_r <= _GEN_180;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            master_in_notify_r <= _GEN_180;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          master_in_notify_r <= _GEN_180;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        master_in_notify_r <= _GEN_180;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      master_in_notify_r <= _GEN_180;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    master_in_notify_r <= _GEN_180;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  master_in_notify_r <= _GEN_180;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            master_in_notify_r <= 1'h0;
                                                                                                                                                          end else begin
                                                                                                                                                            master_in_notify_r <= _GEN_180;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          master_in_notify_r <= _GEN_180;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        master_in_notify_r <= _GEN_180;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      master_in_notify_r <= _GEN_180;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    master_in_notify_r <= _GEN_180;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  master_in_notify_r <= _GEN_180;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                master_in_notify_r <= _GEN_180;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            master_in_notify_r <= _GEN_306;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          master_in_notify_r <= _GEN_306;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        master_in_notify_r <= _GEN_306;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  master_in_notify_r <= 1'h0;
                                                                                                                                                end else begin
                                                                                                                                                  master_in_notify_r <= _GEN_306;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                master_in_notify_r <= _GEN_306;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              master_in_notify_r <= _GEN_306;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            master_in_notify_r <= _GEN_306;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          master_in_notify_r <= _GEN_306;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        master_in_notify_r <= _GEN_306;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      master_in_notify_r <= _GEN_306;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                master_in_notify_r <= 1'h0;
                                                                                                                                              end else begin
                                                                                                                                                master_in_notify_r <= _GEN_306;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              master_in_notify_r <= _GEN_306;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            master_in_notify_r <= _GEN_306;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          master_in_notify_r <= _GEN_306;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        master_in_notify_r <= _GEN_306;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      master_in_notify_r <= _GEN_306;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    master_in_notify_r <= _GEN_306;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              master_in_notify_r <= 1'h0;
                                                                                                                                            end else begin
                                                                                                                                              master_in_notify_r <= _GEN_306;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            master_in_notify_r <= _GEN_306;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          master_in_notify_r <= _GEN_306;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        master_in_notify_r <= _GEN_306;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      master_in_notify_r <= _GEN_306;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    master_in_notify_r <= _GEN_306;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  master_in_notify_r <= _GEN_306;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              master_in_notify_r <= _GEN_432;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    master_in_notify_r <= 1'h0;
                                                                                                                                  end else begin
                                                                                                                                    master_in_notify_r <= _GEN_432;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  master_in_notify_r <= _GEN_432;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                master_in_notify_r <= _GEN_432;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              master_in_notify_r <= _GEN_432;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            master_in_notify_r <= _GEN_432;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  master_in_notify_r <= 1'h0;
                                                                                                                                end else begin
                                                                                                                                  master_in_notify_r <= _GEN_432;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                master_in_notify_r <= _GEN_432;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              master_in_notify_r <= _GEN_432;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            master_in_notify_r <= _GEN_432;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          master_in_notify_r <= _GEN_432;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                master_in_notify_r <= 1'h0;
                                                                                                                              end else begin
                                                                                                                                master_in_notify_r <= _GEN_432;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              master_in_notify_r <= _GEN_432;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            master_in_notify_r <= _GEN_432;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          master_in_notify_r <= _GEN_432;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        master_in_notify_r <= _GEN_432;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    master_in_notify_r <= _GEN_527;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          master_in_notify_r <= 1'h0;
                                                                                                                        end else begin
                                                                                                                          master_in_notify_r <= _GEN_527;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        master_in_notify_r <= _GEN_527;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      master_in_notify_r <= _GEN_527;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    master_in_notify_r <= _GEN_527;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  master_in_notify_r <= _GEN_527;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        master_in_notify_r <= 1'h0;
                                                                                                                      end else begin
                                                                                                                        master_in_notify_r <= _GEN_527;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      master_in_notify_r <= _GEN_527;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    master_in_notify_r <= _GEN_527;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  master_in_notify_r <= _GEN_527;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                master_in_notify_r <= _GEN_527;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      master_in_notify_r <= 1'h0;
                                                                                                                    end else begin
                                                                                                                      master_in_notify_r <= _GEN_527;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    master_in_notify_r <= _GEN_527;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  master_in_notify_r <= _GEN_527;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                master_in_notify_r <= _GEN_527;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              master_in_notify_r <= _GEN_527;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          master_in_notify_r <= _GEN_622;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                master_in_notify_r <= 1'h0;
                                                                                                              end else begin
                                                                                                                master_in_notify_r <= _GEN_622;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              master_in_notify_r <= _GEN_622;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            master_in_notify_r <= _GEN_622;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          master_in_notify_r <= _GEN_622;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        master_in_notify_r <= _GEN_622;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              master_in_notify_r <= 1'h0;
                                                                                                            end else begin
                                                                                                              master_in_notify_r <= _GEN_622;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            master_in_notify_r <= _GEN_622;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          master_in_notify_r <= _GEN_622;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        master_in_notify_r <= _GEN_622;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      master_in_notify_r <= _GEN_622;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            master_in_notify_r <= 1'h0;
                                                                                                          end else begin
                                                                                                            master_in_notify_r <= _GEN_622;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          master_in_notify_r <= _GEN_622;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        master_in_notify_r <= _GEN_622;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      master_in_notify_r <= _GEN_622;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    master_in_notify_r <= _GEN_622;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                master_in_notify_r <= _GEN_717;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      master_in_notify_r <= 1'h0;
                                                                                                    end else begin
                                                                                                      master_in_notify_r <= _GEN_717;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    master_in_notify_r <= _GEN_717;
                                                                                                  end
                                                                                                end else begin
                                                                                                  master_in_notify_r <= _GEN_717;
                                                                                                end
                                                                                              end else begin
                                                                                                master_in_notify_r <= _GEN_717;
                                                                                              end
                                                                                            end else begin
                                                                                              master_in_notify_r <= _GEN_717;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    master_in_notify_r <= 1'h0;
                                                                                                  end else begin
                                                                                                    master_in_notify_r <= _GEN_717;
                                                                                                  end
                                                                                                end else begin
                                                                                                  master_in_notify_r <= _GEN_717;
                                                                                                end
                                                                                              end else begin
                                                                                                master_in_notify_r <= _GEN_717;
                                                                                              end
                                                                                            end else begin
                                                                                              master_in_notify_r <= _GEN_717;
                                                                                            end
                                                                                          end else begin
                                                                                            master_in_notify_r <= _GEN_717;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  master_in_notify_r <= 1'h0;
                                                                                                end else begin
                                                                                                  master_in_notify_r <= _GEN_717;
                                                                                                end
                                                                                              end else begin
                                                                                                master_in_notify_r <= _GEN_717;
                                                                                              end
                                                                                            end else begin
                                                                                              master_in_notify_r <= _GEN_717;
                                                                                            end
                                                                                          end else begin
                                                                                            master_in_notify_r <= _GEN_717;
                                                                                          end
                                                                                        end else begin
                                                                                          master_in_notify_r <= _GEN_717;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      master_in_notify_r <= _GEN_812;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            master_in_notify_r <= 1'h0;
                                                                                          end else begin
                                                                                            master_in_notify_r <= _GEN_812;
                                                                                          end
                                                                                        end else begin
                                                                                          master_in_notify_r <= _GEN_812;
                                                                                        end
                                                                                      end else begin
                                                                                        master_in_notify_r <= _GEN_812;
                                                                                      end
                                                                                    end else begin
                                                                                      master_in_notify_r <= _GEN_812;
                                                                                    end
                                                                                  end else begin
                                                                                    master_in_notify_r <= _GEN_812;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          master_in_notify_r <= 1'h0;
                                                                                        end else begin
                                                                                          master_in_notify_r <= _GEN_812;
                                                                                        end
                                                                                      end else begin
                                                                                        master_in_notify_r <= _GEN_812;
                                                                                      end
                                                                                    end else begin
                                                                                      master_in_notify_r <= _GEN_812;
                                                                                    end
                                                                                  end else begin
                                                                                    master_in_notify_r <= _GEN_812;
                                                                                  end
                                                                                end else begin
                                                                                  master_in_notify_r <= _GEN_812;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        master_in_notify_r <= 1'h0;
                                                                                      end else begin
                                                                                        master_in_notify_r <= _GEN_812;
                                                                                      end
                                                                                    end else begin
                                                                                      master_in_notify_r <= _GEN_812;
                                                                                    end
                                                                                  end else begin
                                                                                    master_in_notify_r <= _GEN_812;
                                                                                  end
                                                                                end else begin
                                                                                  master_in_notify_r <= _GEN_812;
                                                                                end
                                                                              end else begin
                                                                                master_in_notify_r <= _GEN_812;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            master_in_notify_r <= _GEN_907;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  master_in_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  master_in_notify_r <= _GEN_907;
                                                                                end
                                                                              end else begin
                                                                                master_in_notify_r <= _GEN_907;
                                                                              end
                                                                            end else begin
                                                                              master_in_notify_r <= _GEN_907;
                                                                            end
                                                                          end else begin
                                                                            master_in_notify_r <= _GEN_907;
                                                                          end
                                                                        end else begin
                                                                          master_in_notify_r <= _GEN_907;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        master_in_notify_r <= 1'h0;
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  master_in_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  master_in_notify_r <= _GEN_907;
                                                                                end
                                                                              end else begin
                                                                                master_in_notify_r <= _GEN_907;
                                                                              end
                                                                            end else begin
                                                                              master_in_notify_r <= _GEN_907;
                                                                            end
                                                                          end else begin
                                                                            master_in_notify_r <= _GEN_907;
                                                                          end
                                                                        end else begin
                                                                          master_in_notify_r <= _GEN_907;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                master_in_notify_r <= 1'h0;
                                                                              end else begin
                                                                                master_in_notify_r <= _GEN_907;
                                                                              end
                                                                            end else begin
                                                                              master_in_notify_r <= _GEN_907;
                                                                            end
                                                                          end else begin
                                                                            master_in_notify_r <= _GEN_907;
                                                                          end
                                                                        end else begin
                                                                          master_in_notify_r <= _GEN_907;
                                                                        end
                                                                      end else begin
                                                                        master_in_notify_r <= _GEN_907;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (io_slave_out0_sync) begin
                                                                      master_in_notify_r <= 1'h0;
                                                                    end else begin
                                                                      master_in_notify_r <= _GEN_1002;
                                                                    end
                                                                  end else begin
                                                                    master_in_notify_r <= _GEN_1002;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    master_in_notify_r <= 1'h0;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        master_in_notify_r <= 1'h0;
                                                                      end else begin
                                                                        master_in_notify_r <= _GEN_1002;
                                                                      end
                                                                    end else begin
                                                                      master_in_notify_r <= _GEN_1002;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  master_in_notify_r <= _GEN_1034;
                                                                end
                                                              end else begin
                                                                master_in_notify_r <= _GEN_1034;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  master_in_notify_r <= 1'h0;
                                                                end else begin
                                                                  master_in_notify_r <= _GEN_1034;
                                                                end
                                                              end else begin
                                                                master_in_notify_r <= _GEN_1034;
                                                              end
                                                            end else begin
                                                              master_in_notify_r <= _GEN_1034;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              master_in_notify_r <= 1'h0;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    master_in_notify_r <= 1'h0;
                                                                  end else begin
                                                                    master_in_notify_r <= _GEN_1034;
                                                                  end
                                                                end else begin
                                                                  master_in_notify_r <= _GEN_1034;
                                                                end
                                                              end else begin
                                                                master_in_notify_r <= _GEN_1034;
                                                              end
                                                            end
                                                          end else begin
                                                            master_in_notify_r <= _GEN_1088;
                                                          end
                                                        end else begin
                                                          master_in_notify_r <= _GEN_1088;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        master_in_notify_r <= 1'h1;
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              master_in_notify_r <= 1'h0;
                                                            end else begin
                                                              master_in_notify_r <= _GEN_1088;
                                                            end
                                                          end else begin
                                                            master_in_notify_r <= _GEN_1088;
                                                          end
                                                        end else begin
                                                          master_in_notify_r <= _GEN_1088;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            master_in_notify_r <= 1'h0;
                                                          end else begin
                                                            master_in_notify_r <= _GEN_1088;
                                                          end
                                                        end else begin
                                                          master_in_notify_r <= _GEN_1088;
                                                        end
                                                      end else begin
                                                        master_in_notify_r <= _GEN_1088;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    master_in_notify_r <= 1'h0;
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        master_in_notify_r <= 1'h1;
                                                      end else begin
                                                        master_in_notify_r <= _GEN_1142;
                                                      end
                                                    end else begin
                                                      master_in_notify_r <= _GEN_1142;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (io_master_out_sync) begin
                                                      master_in_notify_r <= 1'h1;
                                                    end else begin
                                                      master_in_notify_r <= _GEN_1142;
                                                    end
                                                  end else begin
                                                    master_in_notify_r <= _GEN_1142;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (io_slave_out1_sync) begin
                                                  master_in_notify_r <= 1'h0;
                                                end else begin
                                                  master_in_notify_r <= _GEN_1174;
                                                end
                                              end else begin
                                                master_in_notify_r <= _GEN_1174;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                master_in_notify_r <= 1'h0;
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    master_in_notify_r <= 1'h0;
                                                  end else begin
                                                    master_in_notify_r <= _GEN_1174;
                                                  end
                                                end else begin
                                                  master_in_notify_r <= _GEN_1174;
                                                end
                                              end
                                            end else begin
                                              master_in_notify_r <= _GEN_1206;
                                            end
                                          end else begin
                                            master_in_notify_r <= _GEN_1206;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              master_in_notify_r <= 1'h0;
                                            end else begin
                                              master_in_notify_r <= _GEN_1206;
                                            end
                                          end else begin
                                            master_in_notify_r <= _GEN_1206;
                                          end
                                        end else begin
                                          master_in_notify_r <= _GEN_1206;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          master_in_notify_r <= 1'h0;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                master_in_notify_r <= 1'h0;
                                              end else begin
                                                master_in_notify_r <= _GEN_1206;
                                              end
                                            end else begin
                                              master_in_notify_r <= _GEN_1206;
                                            end
                                          end else begin
                                            master_in_notify_r <= _GEN_1206;
                                          end
                                        end
                                      end else begin
                                        master_in_notify_r <= _GEN_1260;
                                      end
                                    end else begin
                                      master_in_notify_r <= _GEN_1260;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    master_in_notify_r <= 1'h0;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          master_in_notify_r <= 1'h0;
                                        end else begin
                                          master_in_notify_r <= _GEN_1260;
                                        end
                                      end else begin
                                        master_in_notify_r <= _GEN_1260;
                                      end
                                    end else begin
                                      master_in_notify_r <= _GEN_1260;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        master_in_notify_r <= 1'h0;
                                      end else begin
                                        master_in_notify_r <= _GEN_1260;
                                      end
                                    end else begin
                                      master_in_notify_r <= _GEN_1260;
                                    end
                                  end else begin
                                    master_in_notify_r <= _GEN_1260;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (io_slave_out2_sync) begin
                                  master_in_notify_r <= 1'h0;
                                end else begin
                                  master_in_notify_r <= _GEN_1314;
                                end
                              end else begin
                                master_in_notify_r <= _GEN_1314;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                master_in_notify_r <= 1'h0;
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    master_in_notify_r <= 1'h0;
                                  end else begin
                                    master_in_notify_r <= _GEN_1314;
                                  end
                                end else begin
                                  master_in_notify_r <= _GEN_1314;
                                end
                              end
                            end else begin
                              master_in_notify_r <= _GEN_1346;
                            end
                          end else begin
                            master_in_notify_r <= _GEN_1346;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              master_in_notify_r <= 1'h0;
                            end else begin
                              master_in_notify_r <= _GEN_1346;
                            end
                          end else begin
                            master_in_notify_r <= _GEN_1346;
                          end
                        end else begin
                          master_in_notify_r <= _GEN_1346;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          master_in_notify_r <= 1'h0;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                master_in_notify_r <= 1'h0;
                              end else begin
                                master_in_notify_r <= _GEN_1346;
                              end
                            end else begin
                              master_in_notify_r <= _GEN_1346;
                            end
                          end else begin
                            master_in_notify_r <= _GEN_1346;
                          end
                        end
                      end else begin
                        master_in_notify_r <= _GEN_1400;
                      end
                    end else begin
                      master_in_notify_r <= _GEN_1400;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    master_in_notify_r <= 1'h0;
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          master_in_notify_r <= 1'h0;
                        end else begin
                          master_in_notify_r <= _GEN_1400;
                        end
                      end else begin
                        master_in_notify_r <= _GEN_1400;
                      end
                    end else begin
                      master_in_notify_r <= _GEN_1400;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        master_in_notify_r <= 1'h0;
                      end else begin
                        master_in_notify_r <= _GEN_1400;
                      end
                    end else begin
                      master_in_notify_r <= _GEN_1400;
                    end
                  end else begin
                    master_in_notify_r <= _GEN_1400;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (io_slave_out3_sync) begin
                  master_in_notify_r <= 1'h0;
                end else begin
                  master_in_notify_r <= _GEN_1454;
                end
              end else begin
                master_in_notify_r <= _GEN_1454;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                master_in_notify_r <= 1'h0;
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    master_in_notify_r <= 1'h0;
                  end else begin
                    master_in_notify_r <= _GEN_1454;
                  end
                end else begin
                  master_in_notify_r <= _GEN_1454;
                end
              end
            end else begin
              master_in_notify_r <= _GEN_1486;
            end
          end else begin
            master_in_notify_r <= _GEN_1486;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              master_in_notify_r <= 1'h0;
            end else begin
              master_in_notify_r <= _GEN_1486;
            end
          end else begin
            master_in_notify_r <= _GEN_1486;
          end
        end else begin
          master_in_notify_r <= _GEN_1486;
        end
      end
    end
    if (reset) begin
      master_out_notify_r <= 1'h0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            master_out_notify_r <= 1'h1;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  master_out_notify_r <= 1'h1;
                end else begin
                  if (_T_518) begin
                    if (io_slave_out3_sync) begin
                      master_out_notify_r <= 1'h0;
                    end else begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            master_out_notify_r <= 1'h1;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  master_out_notify_r <= 1'h1;
                                end else begin
                                  if (_T_479) begin
                                    if (io_slave_out2_sync) begin
                                      master_out_notify_r <= 1'h0;
                                    end else begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            master_out_notify_r <= 1'h1;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  master_out_notify_r <= 1'h1;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (io_slave_out1_sync) begin
                                                      master_out_notify_r <= 1'h0;
                                                    end else begin
                                                      if (_T_429) begin
                                                        if (io_master_out_sync) begin
                                                          master_out_notify_r <= 1'h0;
                                                        end else begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                master_out_notify_r <= 1'h1;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      master_out_notify_r <= 1'h1;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (io_slave_out0_sync) begin
                                                                          master_out_notify_r <= 1'h0;
                                                                        end else begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    master_out_notify_r <= 1'h0;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              master_out_notify_r <= 1'h0;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        master_out_notify_r <= 1'h0;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  master_out_notify_r <= 1'h0;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            master_out_notify_r <= 1'h0;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      master_out_notify_r <= 1'h0;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    master_out_notify_r <= 1'h1;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  master_out_notify_r <= 1'h1;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            master_out_notify_r <= 1'h0;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      master_out_notify_r <= 1'h0;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    master_out_notify_r <= 1'h0;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  master_out_notify_r <= 1'h0;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                master_out_notify_r <= 1'h0;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    master_out_notify_r <= _GEN_86;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          master_out_notify_r <= 1'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                          master_out_notify_r <= _GEN_86;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        master_out_notify_r <= _GEN_86;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      master_out_notify_r <= _GEN_86;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    master_out_notify_r <= _GEN_86;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  master_out_notify_r <= _GEN_86;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        master_out_notify_r <= 1'h0;
                                                                                                                                                                      end else begin
                                                                                                                                                                        master_out_notify_r <= _GEN_86;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      master_out_notify_r <= _GEN_86;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    master_out_notify_r <= _GEN_86;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  master_out_notify_r <= _GEN_86;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                master_out_notify_r <= _GEN_86;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      master_out_notify_r <= 1'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                      master_out_notify_r <= _GEN_86;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    master_out_notify_r <= _GEN_86;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  master_out_notify_r <= _GEN_86;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                master_out_notify_r <= _GEN_86;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              master_out_notify_r <= _GEN_86;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          master_out_notify_r <= _GEN_181;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        master_out_notify_r <= _GEN_181;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      master_out_notify_r <= _GEN_181;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                master_out_notify_r <= 1'h1;
                                                                                                                                                              end else begin
                                                                                                                                                                master_out_notify_r <= _GEN_181;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              master_out_notify_r <= _GEN_181;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            master_out_notify_r <= _GEN_181;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          master_out_notify_r <= _GEN_181;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        master_out_notify_r <= _GEN_181;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      master_out_notify_r <= _GEN_181;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    master_out_notify_r <= _GEN_181;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              master_out_notify_r <= 1'h1;
                                                                                                                                                            end else begin
                                                                                                                                                              master_out_notify_r <= _GEN_181;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            master_out_notify_r <= _GEN_181;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          master_out_notify_r <= _GEN_181;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        master_out_notify_r <= _GEN_181;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      master_out_notify_r <= _GEN_181;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    master_out_notify_r <= _GEN_181;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  master_out_notify_r <= _GEN_181;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            master_out_notify_r <= 1'h1;
                                                                                                                                                          end else begin
                                                                                                                                                            master_out_notify_r <= _GEN_181;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          master_out_notify_r <= _GEN_181;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        master_out_notify_r <= _GEN_181;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      master_out_notify_r <= _GEN_181;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    master_out_notify_r <= _GEN_181;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  master_out_notify_r <= _GEN_181;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                master_out_notify_r <= _GEN_181;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            master_out_notify_r <= _GEN_307;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          master_out_notify_r <= _GEN_307;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        master_out_notify_r <= _GEN_307;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  master_out_notify_r <= 1'h1;
                                                                                                                                                end else begin
                                                                                                                                                  master_out_notify_r <= _GEN_307;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                master_out_notify_r <= _GEN_307;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              master_out_notify_r <= _GEN_307;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            master_out_notify_r <= _GEN_307;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          master_out_notify_r <= _GEN_307;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        master_out_notify_r <= _GEN_307;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      master_out_notify_r <= _GEN_307;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                master_out_notify_r <= 1'h1;
                                                                                                                                              end else begin
                                                                                                                                                master_out_notify_r <= _GEN_307;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              master_out_notify_r <= _GEN_307;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            master_out_notify_r <= _GEN_307;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          master_out_notify_r <= _GEN_307;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        master_out_notify_r <= _GEN_307;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      master_out_notify_r <= _GEN_307;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    master_out_notify_r <= _GEN_307;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              master_out_notify_r <= 1'h1;
                                                                                                                                            end else begin
                                                                                                                                              master_out_notify_r <= _GEN_307;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            master_out_notify_r <= _GEN_307;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          master_out_notify_r <= _GEN_307;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        master_out_notify_r <= _GEN_307;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      master_out_notify_r <= _GEN_307;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    master_out_notify_r <= _GEN_307;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  master_out_notify_r <= _GEN_307;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              master_out_notify_r <= _GEN_433;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    master_out_notify_r <= 1'h0;
                                                                                                                                  end else begin
                                                                                                                                    master_out_notify_r <= _GEN_433;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  master_out_notify_r <= _GEN_433;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                master_out_notify_r <= _GEN_433;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              master_out_notify_r <= _GEN_433;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            master_out_notify_r <= _GEN_433;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  master_out_notify_r <= 1'h0;
                                                                                                                                end else begin
                                                                                                                                  master_out_notify_r <= _GEN_433;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                master_out_notify_r <= _GEN_433;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              master_out_notify_r <= _GEN_433;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            master_out_notify_r <= _GEN_433;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          master_out_notify_r <= _GEN_433;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                master_out_notify_r <= 1'h0;
                                                                                                                              end else begin
                                                                                                                                master_out_notify_r <= _GEN_433;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              master_out_notify_r <= _GEN_433;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            master_out_notify_r <= _GEN_433;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          master_out_notify_r <= _GEN_433;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        master_out_notify_r <= _GEN_433;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    master_out_notify_r <= _GEN_528;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          master_out_notify_r <= 1'h0;
                                                                                                                        end else begin
                                                                                                                          master_out_notify_r <= _GEN_528;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        master_out_notify_r <= _GEN_528;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      master_out_notify_r <= _GEN_528;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    master_out_notify_r <= _GEN_528;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  master_out_notify_r <= _GEN_528;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        master_out_notify_r <= 1'h0;
                                                                                                                      end else begin
                                                                                                                        master_out_notify_r <= _GEN_528;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      master_out_notify_r <= _GEN_528;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    master_out_notify_r <= _GEN_528;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  master_out_notify_r <= _GEN_528;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                master_out_notify_r <= _GEN_528;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      master_out_notify_r <= 1'h0;
                                                                                                                    end else begin
                                                                                                                      master_out_notify_r <= _GEN_528;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    master_out_notify_r <= _GEN_528;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  master_out_notify_r <= _GEN_528;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                master_out_notify_r <= _GEN_528;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              master_out_notify_r <= _GEN_528;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          master_out_notify_r <= _GEN_623;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                master_out_notify_r <= 1'h0;
                                                                                                              end else begin
                                                                                                                master_out_notify_r <= _GEN_623;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              master_out_notify_r <= _GEN_623;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            master_out_notify_r <= _GEN_623;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          master_out_notify_r <= _GEN_623;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        master_out_notify_r <= _GEN_623;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              master_out_notify_r <= 1'h0;
                                                                                                            end else begin
                                                                                                              master_out_notify_r <= _GEN_623;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            master_out_notify_r <= _GEN_623;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          master_out_notify_r <= _GEN_623;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        master_out_notify_r <= _GEN_623;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      master_out_notify_r <= _GEN_623;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            master_out_notify_r <= 1'h0;
                                                                                                          end else begin
                                                                                                            master_out_notify_r <= _GEN_623;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          master_out_notify_r <= _GEN_623;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        master_out_notify_r <= _GEN_623;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      master_out_notify_r <= _GEN_623;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    master_out_notify_r <= _GEN_623;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                master_out_notify_r <= _GEN_718;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      master_out_notify_r <= 1'h0;
                                                                                                    end else begin
                                                                                                      master_out_notify_r <= _GEN_718;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    master_out_notify_r <= _GEN_718;
                                                                                                  end
                                                                                                end else begin
                                                                                                  master_out_notify_r <= _GEN_718;
                                                                                                end
                                                                                              end else begin
                                                                                                master_out_notify_r <= _GEN_718;
                                                                                              end
                                                                                            end else begin
                                                                                              master_out_notify_r <= _GEN_718;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    master_out_notify_r <= 1'h0;
                                                                                                  end else begin
                                                                                                    master_out_notify_r <= _GEN_718;
                                                                                                  end
                                                                                                end else begin
                                                                                                  master_out_notify_r <= _GEN_718;
                                                                                                end
                                                                                              end else begin
                                                                                                master_out_notify_r <= _GEN_718;
                                                                                              end
                                                                                            end else begin
                                                                                              master_out_notify_r <= _GEN_718;
                                                                                            end
                                                                                          end else begin
                                                                                            master_out_notify_r <= _GEN_718;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  master_out_notify_r <= 1'h0;
                                                                                                end else begin
                                                                                                  master_out_notify_r <= _GEN_718;
                                                                                                end
                                                                                              end else begin
                                                                                                master_out_notify_r <= _GEN_718;
                                                                                              end
                                                                                            end else begin
                                                                                              master_out_notify_r <= _GEN_718;
                                                                                            end
                                                                                          end else begin
                                                                                            master_out_notify_r <= _GEN_718;
                                                                                          end
                                                                                        end else begin
                                                                                          master_out_notify_r <= _GEN_718;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      master_out_notify_r <= _GEN_813;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            master_out_notify_r <= 1'h0;
                                                                                          end else begin
                                                                                            master_out_notify_r <= _GEN_813;
                                                                                          end
                                                                                        end else begin
                                                                                          master_out_notify_r <= _GEN_813;
                                                                                        end
                                                                                      end else begin
                                                                                        master_out_notify_r <= _GEN_813;
                                                                                      end
                                                                                    end else begin
                                                                                      master_out_notify_r <= _GEN_813;
                                                                                    end
                                                                                  end else begin
                                                                                    master_out_notify_r <= _GEN_813;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          master_out_notify_r <= 1'h0;
                                                                                        end else begin
                                                                                          master_out_notify_r <= _GEN_813;
                                                                                        end
                                                                                      end else begin
                                                                                        master_out_notify_r <= _GEN_813;
                                                                                      end
                                                                                    end else begin
                                                                                      master_out_notify_r <= _GEN_813;
                                                                                    end
                                                                                  end else begin
                                                                                    master_out_notify_r <= _GEN_813;
                                                                                  end
                                                                                end else begin
                                                                                  master_out_notify_r <= _GEN_813;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        master_out_notify_r <= 1'h0;
                                                                                      end else begin
                                                                                        master_out_notify_r <= _GEN_813;
                                                                                      end
                                                                                    end else begin
                                                                                      master_out_notify_r <= _GEN_813;
                                                                                    end
                                                                                  end else begin
                                                                                    master_out_notify_r <= _GEN_813;
                                                                                  end
                                                                                end else begin
                                                                                  master_out_notify_r <= _GEN_813;
                                                                                end
                                                                              end else begin
                                                                                master_out_notify_r <= _GEN_813;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            master_out_notify_r <= _GEN_908;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  master_out_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  master_out_notify_r <= _GEN_908;
                                                                                end
                                                                              end else begin
                                                                                master_out_notify_r <= _GEN_908;
                                                                              end
                                                                            end else begin
                                                                              master_out_notify_r <= _GEN_908;
                                                                            end
                                                                          end else begin
                                                                            master_out_notify_r <= _GEN_908;
                                                                          end
                                                                        end else begin
                                                                          master_out_notify_r <= _GEN_908;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        master_out_notify_r <= 1'h0;
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  master_out_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  master_out_notify_r <= _GEN_908;
                                                                                end
                                                                              end else begin
                                                                                master_out_notify_r <= _GEN_908;
                                                                              end
                                                                            end else begin
                                                                              master_out_notify_r <= _GEN_908;
                                                                            end
                                                                          end else begin
                                                                            master_out_notify_r <= _GEN_908;
                                                                          end
                                                                        end else begin
                                                                          master_out_notify_r <= _GEN_908;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                master_out_notify_r <= 1'h0;
                                                                              end else begin
                                                                                master_out_notify_r <= _GEN_908;
                                                                              end
                                                                            end else begin
                                                                              master_out_notify_r <= _GEN_908;
                                                                            end
                                                                          end else begin
                                                                            master_out_notify_r <= _GEN_908;
                                                                          end
                                                                        end else begin
                                                                          master_out_notify_r <= _GEN_908;
                                                                        end
                                                                      end else begin
                                                                        master_out_notify_r <= _GEN_908;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (io_slave_out0_sync) begin
                                                                      master_out_notify_r <= 1'h0;
                                                                    end else begin
                                                                      master_out_notify_r <= _GEN_1003;
                                                                    end
                                                                  end else begin
                                                                    master_out_notify_r <= _GEN_1003;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    master_out_notify_r <= 1'h1;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        master_out_notify_r <= 1'h0;
                                                                      end else begin
                                                                        master_out_notify_r <= _GEN_1003;
                                                                      end
                                                                    end else begin
                                                                      master_out_notify_r <= _GEN_1003;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  master_out_notify_r <= _GEN_1035;
                                                                end
                                                              end else begin
                                                                master_out_notify_r <= _GEN_1035;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  master_out_notify_r <= 1'h1;
                                                                end else begin
                                                                  master_out_notify_r <= _GEN_1035;
                                                                end
                                                              end else begin
                                                                master_out_notify_r <= _GEN_1035;
                                                              end
                                                            end else begin
                                                              master_out_notify_r <= _GEN_1035;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              master_out_notify_r <= 1'h1;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    master_out_notify_r <= 1'h1;
                                                                  end else begin
                                                                    master_out_notify_r <= _GEN_1035;
                                                                  end
                                                                end else begin
                                                                  master_out_notify_r <= _GEN_1035;
                                                                end
                                                              end else begin
                                                                master_out_notify_r <= _GEN_1035;
                                                              end
                                                            end
                                                          end else begin
                                                            master_out_notify_r <= _GEN_1089;
                                                          end
                                                        end else begin
                                                          master_out_notify_r <= _GEN_1089;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        master_out_notify_r <= 1'h0;
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              master_out_notify_r <= 1'h1;
                                                            end else begin
                                                              master_out_notify_r <= _GEN_1089;
                                                            end
                                                          end else begin
                                                            master_out_notify_r <= _GEN_1089;
                                                          end
                                                        end else begin
                                                          master_out_notify_r <= _GEN_1089;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            master_out_notify_r <= 1'h1;
                                                          end else begin
                                                            master_out_notify_r <= _GEN_1089;
                                                          end
                                                        end else begin
                                                          master_out_notify_r <= _GEN_1089;
                                                        end
                                                      end else begin
                                                        master_out_notify_r <= _GEN_1089;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    master_out_notify_r <= 1'h0;
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        master_out_notify_r <= 1'h0;
                                                      end else begin
                                                        master_out_notify_r <= _GEN_1143;
                                                      end
                                                    end else begin
                                                      master_out_notify_r <= _GEN_1143;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (io_master_out_sync) begin
                                                      master_out_notify_r <= 1'h0;
                                                    end else begin
                                                      master_out_notify_r <= _GEN_1143;
                                                    end
                                                  end else begin
                                                    master_out_notify_r <= _GEN_1143;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (io_slave_out1_sync) begin
                                                  master_out_notify_r <= 1'h0;
                                                end else begin
                                                  master_out_notify_r <= _GEN_1175;
                                                end
                                              end else begin
                                                master_out_notify_r <= _GEN_1175;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                master_out_notify_r <= 1'h1;
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    master_out_notify_r <= 1'h0;
                                                  end else begin
                                                    master_out_notify_r <= _GEN_1175;
                                                  end
                                                end else begin
                                                  master_out_notify_r <= _GEN_1175;
                                                end
                                              end
                                            end else begin
                                              master_out_notify_r <= _GEN_1207;
                                            end
                                          end else begin
                                            master_out_notify_r <= _GEN_1207;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              master_out_notify_r <= 1'h1;
                                            end else begin
                                              master_out_notify_r <= _GEN_1207;
                                            end
                                          end else begin
                                            master_out_notify_r <= _GEN_1207;
                                          end
                                        end else begin
                                          master_out_notify_r <= _GEN_1207;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          master_out_notify_r <= 1'h1;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                master_out_notify_r <= 1'h1;
                                              end else begin
                                                master_out_notify_r <= _GEN_1207;
                                              end
                                            end else begin
                                              master_out_notify_r <= _GEN_1207;
                                            end
                                          end else begin
                                            master_out_notify_r <= _GEN_1207;
                                          end
                                        end
                                      end else begin
                                        master_out_notify_r <= _GEN_1261;
                                      end
                                    end else begin
                                      master_out_notify_r <= _GEN_1261;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    master_out_notify_r <= 1'h0;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          master_out_notify_r <= 1'h1;
                                        end else begin
                                          master_out_notify_r <= _GEN_1261;
                                        end
                                      end else begin
                                        master_out_notify_r <= _GEN_1261;
                                      end
                                    end else begin
                                      master_out_notify_r <= _GEN_1261;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        master_out_notify_r <= 1'h1;
                                      end else begin
                                        master_out_notify_r <= _GEN_1261;
                                      end
                                    end else begin
                                      master_out_notify_r <= _GEN_1261;
                                    end
                                  end else begin
                                    master_out_notify_r <= _GEN_1261;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (io_slave_out2_sync) begin
                                  master_out_notify_r <= 1'h0;
                                end else begin
                                  master_out_notify_r <= _GEN_1315;
                                end
                              end else begin
                                master_out_notify_r <= _GEN_1315;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                master_out_notify_r <= 1'h1;
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    master_out_notify_r <= 1'h0;
                                  end else begin
                                    master_out_notify_r <= _GEN_1315;
                                  end
                                end else begin
                                  master_out_notify_r <= _GEN_1315;
                                end
                              end
                            end else begin
                              master_out_notify_r <= _GEN_1347;
                            end
                          end else begin
                            master_out_notify_r <= _GEN_1347;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              master_out_notify_r <= 1'h1;
                            end else begin
                              master_out_notify_r <= _GEN_1347;
                            end
                          end else begin
                            master_out_notify_r <= _GEN_1347;
                          end
                        end else begin
                          master_out_notify_r <= _GEN_1347;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          master_out_notify_r <= 1'h1;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                master_out_notify_r <= 1'h1;
                              end else begin
                                master_out_notify_r <= _GEN_1347;
                              end
                            end else begin
                              master_out_notify_r <= _GEN_1347;
                            end
                          end else begin
                            master_out_notify_r <= _GEN_1347;
                          end
                        end
                      end else begin
                        master_out_notify_r <= _GEN_1401;
                      end
                    end else begin
                      master_out_notify_r <= _GEN_1401;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    master_out_notify_r <= 1'h0;
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          master_out_notify_r <= 1'h1;
                        end else begin
                          master_out_notify_r <= _GEN_1401;
                        end
                      end else begin
                        master_out_notify_r <= _GEN_1401;
                      end
                    end else begin
                      master_out_notify_r <= _GEN_1401;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        master_out_notify_r <= 1'h1;
                      end else begin
                        master_out_notify_r <= _GEN_1401;
                      end
                    end else begin
                      master_out_notify_r <= _GEN_1401;
                    end
                  end else begin
                    master_out_notify_r <= _GEN_1401;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (io_slave_out3_sync) begin
                  master_out_notify_r <= 1'h0;
                end else begin
                  master_out_notify_r <= _GEN_1455;
                end
              end else begin
                master_out_notify_r <= _GEN_1455;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                master_out_notify_r <= 1'h1;
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    master_out_notify_r <= 1'h0;
                  end else begin
                    master_out_notify_r <= _GEN_1455;
                  end
                end else begin
                  master_out_notify_r <= _GEN_1455;
                end
              end
            end else begin
              master_out_notify_r <= _GEN_1487;
            end
          end else begin
            master_out_notify_r <= _GEN_1487;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              master_out_notify_r <= 1'h1;
            end else begin
              master_out_notify_r <= _GEN_1487;
            end
          end else begin
            master_out_notify_r <= _GEN_1487;
          end
        end else begin
          master_out_notify_r <= _GEN_1487;
        end
      end
    end
    if (reset) begin
      slave_in0_notify_r <= 1'h0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            slave_in0_notify_r <= 1'h0;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  slave_in0_notify_r <= 1'h0;
                end else begin
                  if (_T_518) begin
                    if (io_slave_out3_sync) begin
                      slave_in0_notify_r <= 1'h0;
                    end else begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            slave_in0_notify_r <= 1'h0;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  slave_in0_notify_r <= 1'h0;
                                end else begin
                                  if (_T_479) begin
                                    if (io_slave_out2_sync) begin
                                      slave_in0_notify_r <= 1'h0;
                                    end else begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            slave_in0_notify_r <= 1'h0;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  slave_in0_notify_r <= 1'h0;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (io_slave_out1_sync) begin
                                                      slave_in0_notify_r <= 1'h0;
                                                    end else begin
                                                      if (_T_429) begin
                                                        if (io_master_out_sync) begin
                                                          slave_in0_notify_r <= 1'h0;
                                                        end else begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                slave_in0_notify_r <= 1'h0;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      slave_in0_notify_r <= 1'h0;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (io_slave_out0_sync) begin
                                                                          slave_in0_notify_r <= 1'h1;
                                                                        end else begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    slave_in0_notify_r <= 1'h0;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              slave_in0_notify_r <= 1'h0;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        slave_in0_notify_r <= 1'h0;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  slave_in0_notify_r <= 1'h0;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            slave_in0_notify_r <= 1'h0;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      slave_in0_notify_r <= 1'h0;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    slave_in0_notify_r <= 1'h0;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  slave_in0_notify_r <= 1'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            slave_in0_notify_r <= 1'h0;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      slave_in0_notify_r <= 1'h0;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    slave_in0_notify_r <= 1'h0;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  slave_in0_notify_r <= 1'h0;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                slave_in0_notify_r <= 1'h0;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          slave_in0_notify_r <= 1'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                          slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        slave_in0_notify_r <= 1'h0;
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_in0_notify_r <= _GEN_87;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      slave_in0_notify_r <= 1'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_in0_notify_r <= _GEN_87;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_in0_notify_r <= _GEN_87;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_in0_notify_r <= _GEN_87;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in0_notify_r <= _GEN_182;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in0_notify_r <= _GEN_182;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in0_notify_r <= _GEN_182;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                slave_in0_notify_r <= 1'h0;
                                                                                                                                                              end else begin
                                                                                                                                                                slave_in0_notify_r <= _GEN_182;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_in0_notify_r <= _GEN_182;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_in0_notify_r <= _GEN_182;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in0_notify_r <= _GEN_182;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in0_notify_r <= _GEN_182;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in0_notify_r <= _GEN_182;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_in0_notify_r <= _GEN_182;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              slave_in0_notify_r <= 1'h0;
                                                                                                                                                            end else begin
                                                                                                                                                              slave_in0_notify_r <= _GEN_182;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_in0_notify_r <= _GEN_182;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in0_notify_r <= _GEN_182;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in0_notify_r <= _GEN_182;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in0_notify_r <= _GEN_182;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_in0_notify_r <= _GEN_182;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_in0_notify_r <= _GEN_182;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            slave_in0_notify_r <= 1'h0;
                                                                                                                                                          end else begin
                                                                                                                                                            slave_in0_notify_r <= _GEN_182;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in0_notify_r <= _GEN_182;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in0_notify_r <= _GEN_182;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in0_notify_r <= _GEN_182;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_in0_notify_r <= _GEN_182;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_in0_notify_r <= _GEN_182;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_in0_notify_r <= _GEN_182;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in0_notify_r <= _GEN_308;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in0_notify_r <= _GEN_308;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in0_notify_r <= _GEN_308;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  slave_in0_notify_r <= 1'h0;
                                                                                                                                                end else begin
                                                                                                                                                  slave_in0_notify_r <= _GEN_308;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_in0_notify_r <= _GEN_308;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_in0_notify_r <= _GEN_308;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in0_notify_r <= _GEN_308;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in0_notify_r <= _GEN_308;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in0_notify_r <= _GEN_308;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_in0_notify_r <= _GEN_308;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                slave_in0_notify_r <= 1'h0;
                                                                                                                                              end else begin
                                                                                                                                                slave_in0_notify_r <= _GEN_308;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_in0_notify_r <= _GEN_308;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in0_notify_r <= _GEN_308;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in0_notify_r <= _GEN_308;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in0_notify_r <= _GEN_308;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_in0_notify_r <= _GEN_308;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_in0_notify_r <= _GEN_308;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              slave_in0_notify_r <= 1'h0;
                                                                                                                                            end else begin
                                                                                                                                              slave_in0_notify_r <= _GEN_308;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in0_notify_r <= _GEN_308;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in0_notify_r <= _GEN_308;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in0_notify_r <= _GEN_308;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_in0_notify_r <= _GEN_308;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_in0_notify_r <= _GEN_308;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_in0_notify_r <= _GEN_308;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in0_notify_r <= _GEN_434;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    slave_in0_notify_r <= 1'h0;
                                                                                                                                  end else begin
                                                                                                                                    slave_in0_notify_r <= _GEN_434;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_in0_notify_r <= _GEN_434;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_in0_notify_r <= _GEN_434;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in0_notify_r <= _GEN_434;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_in0_notify_r <= _GEN_434;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  slave_in0_notify_r <= 1'h0;
                                                                                                                                end else begin
                                                                                                                                  slave_in0_notify_r <= _GEN_434;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_in0_notify_r <= _GEN_434;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in0_notify_r <= _GEN_434;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_in0_notify_r <= _GEN_434;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_in0_notify_r <= _GEN_434;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                slave_in0_notify_r <= 1'h0;
                                                                                                                              end else begin
                                                                                                                                slave_in0_notify_r <= _GEN_434;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in0_notify_r <= _GEN_434;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_in0_notify_r <= _GEN_434;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_in0_notify_r <= _GEN_434;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_in0_notify_r <= _GEN_434;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in0_notify_r <= _GEN_529;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          slave_in0_notify_r <= 1'h0;
                                                                                                                        end else begin
                                                                                                                          slave_in0_notify_r <= _GEN_529;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_in0_notify_r <= _GEN_529;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_in0_notify_r <= _GEN_529;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in0_notify_r <= _GEN_529;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_in0_notify_r <= _GEN_529;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        slave_in0_notify_r <= 1'h0;
                                                                                                                      end else begin
                                                                                                                        slave_in0_notify_r <= _GEN_529;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_in0_notify_r <= _GEN_529;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in0_notify_r <= _GEN_529;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_in0_notify_r <= _GEN_529;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_in0_notify_r <= _GEN_529;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      slave_in0_notify_r <= 1'h0;
                                                                                                                    end else begin
                                                                                                                      slave_in0_notify_r <= _GEN_529;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in0_notify_r <= _GEN_529;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_in0_notify_r <= _GEN_529;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_in0_notify_r <= _GEN_529;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_in0_notify_r <= _GEN_529;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in0_notify_r <= _GEN_624;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                slave_in0_notify_r <= 1'h0;
                                                                                                              end else begin
                                                                                                                slave_in0_notify_r <= _GEN_624;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_in0_notify_r <= _GEN_624;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_in0_notify_r <= _GEN_624;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in0_notify_r <= _GEN_624;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_in0_notify_r <= _GEN_624;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              slave_in0_notify_r <= 1'h0;
                                                                                                            end else begin
                                                                                                              slave_in0_notify_r <= _GEN_624;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_in0_notify_r <= _GEN_624;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in0_notify_r <= _GEN_624;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_in0_notify_r <= _GEN_624;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_in0_notify_r <= _GEN_624;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            slave_in0_notify_r <= 1'h0;
                                                                                                          end else begin
                                                                                                            slave_in0_notify_r <= _GEN_624;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in0_notify_r <= _GEN_624;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_in0_notify_r <= _GEN_624;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_in0_notify_r <= _GEN_624;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_in0_notify_r <= _GEN_624;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in0_notify_r <= _GEN_719;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      slave_in0_notify_r <= 1'h0;
                                                                                                    end else begin
                                                                                                      slave_in0_notify_r <= _GEN_719;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_in0_notify_r <= _GEN_719;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_in0_notify_r <= _GEN_719;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in0_notify_r <= _GEN_719;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_in0_notify_r <= _GEN_719;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    slave_in0_notify_r <= 1'h0;
                                                                                                  end else begin
                                                                                                    slave_in0_notify_r <= _GEN_719;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_in0_notify_r <= _GEN_719;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in0_notify_r <= _GEN_719;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_in0_notify_r <= _GEN_719;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_in0_notify_r <= _GEN_719;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  slave_in0_notify_r <= 1'h0;
                                                                                                end else begin
                                                                                                  slave_in0_notify_r <= _GEN_719;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in0_notify_r <= _GEN_719;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_in0_notify_r <= _GEN_719;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_in0_notify_r <= _GEN_719;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_in0_notify_r <= _GEN_719;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in0_notify_r <= _GEN_814;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            slave_in0_notify_r <= 1'h0;
                                                                                          end else begin
                                                                                            slave_in0_notify_r <= _GEN_814;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_in0_notify_r <= _GEN_814;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_in0_notify_r <= _GEN_814;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in0_notify_r <= _GEN_814;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_in0_notify_r <= _GEN_814;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          slave_in0_notify_r <= 1'h0;
                                                                                        end else begin
                                                                                          slave_in0_notify_r <= _GEN_814;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_in0_notify_r <= _GEN_814;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in0_notify_r <= _GEN_814;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_in0_notify_r <= _GEN_814;
                                                                                  end
                                                                                end else begin
                                                                                  slave_in0_notify_r <= _GEN_814;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        slave_in0_notify_r <= 1'h0;
                                                                                      end else begin
                                                                                        slave_in0_notify_r <= _GEN_814;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in0_notify_r <= _GEN_814;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_in0_notify_r <= _GEN_814;
                                                                                  end
                                                                                end else begin
                                                                                  slave_in0_notify_r <= _GEN_814;
                                                                                end
                                                                              end else begin
                                                                                slave_in0_notify_r <= _GEN_814;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            slave_in0_notify_r <= _GEN_909;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_in0_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_in0_notify_r <= _GEN_909;
                                                                                end
                                                                              end else begin
                                                                                slave_in0_notify_r <= _GEN_909;
                                                                              end
                                                                            end else begin
                                                                              slave_in0_notify_r <= _GEN_909;
                                                                            end
                                                                          end else begin
                                                                            slave_in0_notify_r <= _GEN_909;
                                                                          end
                                                                        end else begin
                                                                          slave_in0_notify_r <= _GEN_909;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_in0_notify_r <= 1'h1;
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_in0_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_in0_notify_r <= _GEN_909;
                                                                                end
                                                                              end else begin
                                                                                slave_in0_notify_r <= _GEN_909;
                                                                              end
                                                                            end else begin
                                                                              slave_in0_notify_r <= _GEN_909;
                                                                            end
                                                                          end else begin
                                                                            slave_in0_notify_r <= _GEN_909;
                                                                          end
                                                                        end else begin
                                                                          slave_in0_notify_r <= _GEN_909;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                slave_in0_notify_r <= 1'h0;
                                                                              end else begin
                                                                                slave_in0_notify_r <= _GEN_909;
                                                                              end
                                                                            end else begin
                                                                              slave_in0_notify_r <= _GEN_909;
                                                                            end
                                                                          end else begin
                                                                            slave_in0_notify_r <= _GEN_909;
                                                                          end
                                                                        end else begin
                                                                          slave_in0_notify_r <= _GEN_909;
                                                                        end
                                                                      end else begin
                                                                        slave_in0_notify_r <= _GEN_909;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (io_slave_out0_sync) begin
                                                                      slave_in0_notify_r <= 1'h1;
                                                                    end else begin
                                                                      slave_in0_notify_r <= _GEN_1004;
                                                                    end
                                                                  end else begin
                                                                    slave_in0_notify_r <= _GEN_1004;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_in0_notify_r <= 1'h0;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_in0_notify_r <= 1'h1;
                                                                      end else begin
                                                                        slave_in0_notify_r <= _GEN_1004;
                                                                      end
                                                                    end else begin
                                                                      slave_in0_notify_r <= _GEN_1004;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  slave_in0_notify_r <= _GEN_1036;
                                                                end
                                                              end else begin
                                                                slave_in0_notify_r <= _GEN_1036;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  slave_in0_notify_r <= 1'h0;
                                                                end else begin
                                                                  slave_in0_notify_r <= _GEN_1036;
                                                                end
                                                              end else begin
                                                                slave_in0_notify_r <= _GEN_1036;
                                                              end
                                                            end else begin
                                                              slave_in0_notify_r <= _GEN_1036;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_in0_notify_r <= 1'h0;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_in0_notify_r <= 1'h0;
                                                                  end else begin
                                                                    slave_in0_notify_r <= _GEN_1036;
                                                                  end
                                                                end else begin
                                                                  slave_in0_notify_r <= _GEN_1036;
                                                                end
                                                              end else begin
                                                                slave_in0_notify_r <= _GEN_1036;
                                                              end
                                                            end
                                                          end else begin
                                                            slave_in0_notify_r <= _GEN_1090;
                                                          end
                                                        end else begin
                                                          slave_in0_notify_r <= _GEN_1090;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_in0_notify_r <= 1'h0;
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_in0_notify_r <= 1'h0;
                                                            end else begin
                                                              slave_in0_notify_r <= _GEN_1090;
                                                            end
                                                          end else begin
                                                            slave_in0_notify_r <= _GEN_1090;
                                                          end
                                                        end else begin
                                                          slave_in0_notify_r <= _GEN_1090;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            slave_in0_notify_r <= 1'h0;
                                                          end else begin
                                                            slave_in0_notify_r <= _GEN_1090;
                                                          end
                                                        end else begin
                                                          slave_in0_notify_r <= _GEN_1090;
                                                        end
                                                      end else begin
                                                        slave_in0_notify_r <= _GEN_1090;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_in0_notify_r <= 1'h0;
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_in0_notify_r <= 1'h0;
                                                      end else begin
                                                        slave_in0_notify_r <= _GEN_1144;
                                                      end
                                                    end else begin
                                                      slave_in0_notify_r <= _GEN_1144;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (io_master_out_sync) begin
                                                      slave_in0_notify_r <= 1'h0;
                                                    end else begin
                                                      slave_in0_notify_r <= _GEN_1144;
                                                    end
                                                  end else begin
                                                    slave_in0_notify_r <= _GEN_1144;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (io_slave_out1_sync) begin
                                                  slave_in0_notify_r <= 1'h0;
                                                end else begin
                                                  slave_in0_notify_r <= _GEN_1176;
                                                end
                                              end else begin
                                                slave_in0_notify_r <= _GEN_1176;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_in0_notify_r <= 1'h0;
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_in0_notify_r <= 1'h0;
                                                  end else begin
                                                    slave_in0_notify_r <= _GEN_1176;
                                                  end
                                                end else begin
                                                  slave_in0_notify_r <= _GEN_1176;
                                                end
                                              end
                                            end else begin
                                              slave_in0_notify_r <= _GEN_1208;
                                            end
                                          end else begin
                                            slave_in0_notify_r <= _GEN_1208;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              slave_in0_notify_r <= 1'h0;
                                            end else begin
                                              slave_in0_notify_r <= _GEN_1208;
                                            end
                                          end else begin
                                            slave_in0_notify_r <= _GEN_1208;
                                          end
                                        end else begin
                                          slave_in0_notify_r <= _GEN_1208;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_in0_notify_r <= 1'h0;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_in0_notify_r <= 1'h0;
                                              end else begin
                                                slave_in0_notify_r <= _GEN_1208;
                                              end
                                            end else begin
                                              slave_in0_notify_r <= _GEN_1208;
                                            end
                                          end else begin
                                            slave_in0_notify_r <= _GEN_1208;
                                          end
                                        end
                                      end else begin
                                        slave_in0_notify_r <= _GEN_1262;
                                      end
                                    end else begin
                                      slave_in0_notify_r <= _GEN_1262;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_in0_notify_r <= 1'h0;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_in0_notify_r <= 1'h0;
                                        end else begin
                                          slave_in0_notify_r <= _GEN_1262;
                                        end
                                      end else begin
                                        slave_in0_notify_r <= _GEN_1262;
                                      end
                                    end else begin
                                      slave_in0_notify_r <= _GEN_1262;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        slave_in0_notify_r <= 1'h0;
                                      end else begin
                                        slave_in0_notify_r <= _GEN_1262;
                                      end
                                    end else begin
                                      slave_in0_notify_r <= _GEN_1262;
                                    end
                                  end else begin
                                    slave_in0_notify_r <= _GEN_1262;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (io_slave_out2_sync) begin
                                  slave_in0_notify_r <= 1'h0;
                                end else begin
                                  slave_in0_notify_r <= _GEN_1316;
                                end
                              end else begin
                                slave_in0_notify_r <= _GEN_1316;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_in0_notify_r <= 1'h0;
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_in0_notify_r <= 1'h0;
                                  end else begin
                                    slave_in0_notify_r <= _GEN_1316;
                                  end
                                end else begin
                                  slave_in0_notify_r <= _GEN_1316;
                                end
                              end
                            end else begin
                              slave_in0_notify_r <= _GEN_1348;
                            end
                          end else begin
                            slave_in0_notify_r <= _GEN_1348;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              slave_in0_notify_r <= 1'h0;
                            end else begin
                              slave_in0_notify_r <= _GEN_1348;
                            end
                          end else begin
                            slave_in0_notify_r <= _GEN_1348;
                          end
                        end else begin
                          slave_in0_notify_r <= _GEN_1348;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_in0_notify_r <= 1'h0;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_in0_notify_r <= 1'h0;
                              end else begin
                                slave_in0_notify_r <= _GEN_1348;
                              end
                            end else begin
                              slave_in0_notify_r <= _GEN_1348;
                            end
                          end else begin
                            slave_in0_notify_r <= _GEN_1348;
                          end
                        end
                      end else begin
                        slave_in0_notify_r <= _GEN_1402;
                      end
                    end else begin
                      slave_in0_notify_r <= _GEN_1402;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_in0_notify_r <= 1'h0;
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_in0_notify_r <= 1'h0;
                        end else begin
                          slave_in0_notify_r <= _GEN_1402;
                        end
                      end else begin
                        slave_in0_notify_r <= _GEN_1402;
                      end
                    end else begin
                      slave_in0_notify_r <= _GEN_1402;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        slave_in0_notify_r <= 1'h0;
                      end else begin
                        slave_in0_notify_r <= _GEN_1402;
                      end
                    end else begin
                      slave_in0_notify_r <= _GEN_1402;
                    end
                  end else begin
                    slave_in0_notify_r <= _GEN_1402;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (io_slave_out3_sync) begin
                  slave_in0_notify_r <= 1'h0;
                end else begin
                  slave_in0_notify_r <= _GEN_1456;
                end
              end else begin
                slave_in0_notify_r <= _GEN_1456;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                slave_in0_notify_r <= 1'h0;
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_in0_notify_r <= 1'h0;
                  end else begin
                    slave_in0_notify_r <= _GEN_1456;
                  end
                end else begin
                  slave_in0_notify_r <= _GEN_1456;
                end
              end
            end else begin
              slave_in0_notify_r <= _GEN_1488;
            end
          end else begin
            slave_in0_notify_r <= _GEN_1488;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              slave_in0_notify_r <= 1'h0;
            end else begin
              slave_in0_notify_r <= _GEN_1488;
            end
          end else begin
            slave_in0_notify_r <= _GEN_1488;
          end
        end else begin
          slave_in0_notify_r <= _GEN_1488;
        end
      end
    end
    if (reset) begin
      slave_in1_notify_r <= 1'h0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            slave_in1_notify_r <= 1'h0;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  slave_in1_notify_r <= 1'h0;
                end else begin
                  if (_T_518) begin
                    if (io_slave_out3_sync) begin
                      slave_in1_notify_r <= 1'h0;
                    end else begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            slave_in1_notify_r <= 1'h0;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  slave_in1_notify_r <= 1'h0;
                                end else begin
                                  if (_T_479) begin
                                    if (io_slave_out2_sync) begin
                                      slave_in1_notify_r <= 1'h0;
                                    end else begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            slave_in1_notify_r <= 1'h0;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  slave_in1_notify_r <= 1'h0;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (io_slave_out1_sync) begin
                                                      slave_in1_notify_r <= 1'h1;
                                                    end else begin
                                                      if (_T_429) begin
                                                        if (io_master_out_sync) begin
                                                          slave_in1_notify_r <= 1'h0;
                                                        end else begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                slave_in1_notify_r <= 1'h0;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      slave_in1_notify_r <= 1'h0;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (io_slave_out0_sync) begin
                                                                          slave_in1_notify_r <= 1'h0;
                                                                        end else begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    slave_in1_notify_r <= 1'h0;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              slave_in1_notify_r <= 1'h0;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        slave_in1_notify_r <= 1'h0;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  slave_in1_notify_r <= 1'h0;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            slave_in1_notify_r <= 1'h0;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      slave_in1_notify_r <= 1'h0;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    slave_in1_notify_r <= 1'h0;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  slave_in1_notify_r <= 1'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            slave_in1_notify_r <= 1'h0;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      slave_in1_notify_r <= 1'h0;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    slave_in1_notify_r <= 1'h0;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  slave_in1_notify_r <= 1'h0;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                slave_in1_notify_r <= 1'h0;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          slave_in1_notify_r <= 1'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                          slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        slave_in1_notify_r <= 1'h0;
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_in1_notify_r <= _GEN_88;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      slave_in1_notify_r <= 1'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_in1_notify_r <= _GEN_88;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_in1_notify_r <= _GEN_88;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_in1_notify_r <= _GEN_88;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in1_notify_r <= _GEN_183;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in1_notify_r <= _GEN_183;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in1_notify_r <= _GEN_183;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                slave_in1_notify_r <= 1'h0;
                                                                                                                                                              end else begin
                                                                                                                                                                slave_in1_notify_r <= _GEN_183;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_in1_notify_r <= _GEN_183;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_in1_notify_r <= _GEN_183;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in1_notify_r <= _GEN_183;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in1_notify_r <= _GEN_183;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in1_notify_r <= _GEN_183;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_in1_notify_r <= _GEN_183;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              slave_in1_notify_r <= 1'h0;
                                                                                                                                                            end else begin
                                                                                                                                                              slave_in1_notify_r <= _GEN_183;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_in1_notify_r <= _GEN_183;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in1_notify_r <= _GEN_183;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in1_notify_r <= _GEN_183;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in1_notify_r <= _GEN_183;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_in1_notify_r <= _GEN_183;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_in1_notify_r <= _GEN_183;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            slave_in1_notify_r <= 1'h0;
                                                                                                                                                          end else begin
                                                                                                                                                            slave_in1_notify_r <= _GEN_183;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in1_notify_r <= _GEN_183;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in1_notify_r <= _GEN_183;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in1_notify_r <= _GEN_183;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_in1_notify_r <= _GEN_183;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_in1_notify_r <= _GEN_183;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_in1_notify_r <= _GEN_183;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in1_notify_r <= _GEN_309;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in1_notify_r <= _GEN_309;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in1_notify_r <= _GEN_309;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  slave_in1_notify_r <= 1'h0;
                                                                                                                                                end else begin
                                                                                                                                                  slave_in1_notify_r <= _GEN_309;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_in1_notify_r <= _GEN_309;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_in1_notify_r <= _GEN_309;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in1_notify_r <= _GEN_309;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in1_notify_r <= _GEN_309;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in1_notify_r <= _GEN_309;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_in1_notify_r <= _GEN_309;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                slave_in1_notify_r <= 1'h0;
                                                                                                                                              end else begin
                                                                                                                                                slave_in1_notify_r <= _GEN_309;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_in1_notify_r <= _GEN_309;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in1_notify_r <= _GEN_309;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in1_notify_r <= _GEN_309;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in1_notify_r <= _GEN_309;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_in1_notify_r <= _GEN_309;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_in1_notify_r <= _GEN_309;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              slave_in1_notify_r <= 1'h0;
                                                                                                                                            end else begin
                                                                                                                                              slave_in1_notify_r <= _GEN_309;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in1_notify_r <= _GEN_309;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in1_notify_r <= _GEN_309;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in1_notify_r <= _GEN_309;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_in1_notify_r <= _GEN_309;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_in1_notify_r <= _GEN_309;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_in1_notify_r <= _GEN_309;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in1_notify_r <= _GEN_435;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    slave_in1_notify_r <= 1'h0;
                                                                                                                                  end else begin
                                                                                                                                    slave_in1_notify_r <= _GEN_435;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_in1_notify_r <= _GEN_435;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_in1_notify_r <= _GEN_435;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in1_notify_r <= _GEN_435;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_in1_notify_r <= _GEN_435;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  slave_in1_notify_r <= 1'h0;
                                                                                                                                end else begin
                                                                                                                                  slave_in1_notify_r <= _GEN_435;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_in1_notify_r <= _GEN_435;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in1_notify_r <= _GEN_435;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_in1_notify_r <= _GEN_435;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_in1_notify_r <= _GEN_435;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                slave_in1_notify_r <= 1'h0;
                                                                                                                              end else begin
                                                                                                                                slave_in1_notify_r <= _GEN_435;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in1_notify_r <= _GEN_435;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_in1_notify_r <= _GEN_435;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_in1_notify_r <= _GEN_435;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_in1_notify_r <= _GEN_435;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in1_notify_r <= _GEN_530;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          slave_in1_notify_r <= 1'h0;
                                                                                                                        end else begin
                                                                                                                          slave_in1_notify_r <= _GEN_530;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_in1_notify_r <= _GEN_530;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_in1_notify_r <= _GEN_530;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in1_notify_r <= _GEN_530;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_in1_notify_r <= _GEN_530;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        slave_in1_notify_r <= 1'h0;
                                                                                                                      end else begin
                                                                                                                        slave_in1_notify_r <= _GEN_530;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_in1_notify_r <= _GEN_530;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in1_notify_r <= _GEN_530;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_in1_notify_r <= _GEN_530;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_in1_notify_r <= _GEN_530;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      slave_in1_notify_r <= 1'h0;
                                                                                                                    end else begin
                                                                                                                      slave_in1_notify_r <= _GEN_530;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in1_notify_r <= _GEN_530;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_in1_notify_r <= _GEN_530;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_in1_notify_r <= _GEN_530;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_in1_notify_r <= _GEN_530;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in1_notify_r <= _GEN_625;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                slave_in1_notify_r <= 1'h0;
                                                                                                              end else begin
                                                                                                                slave_in1_notify_r <= _GEN_625;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_in1_notify_r <= _GEN_625;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_in1_notify_r <= _GEN_625;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in1_notify_r <= _GEN_625;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_in1_notify_r <= _GEN_625;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              slave_in1_notify_r <= 1'h0;
                                                                                                            end else begin
                                                                                                              slave_in1_notify_r <= _GEN_625;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_in1_notify_r <= _GEN_625;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in1_notify_r <= _GEN_625;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_in1_notify_r <= _GEN_625;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_in1_notify_r <= _GEN_625;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            slave_in1_notify_r <= 1'h0;
                                                                                                          end else begin
                                                                                                            slave_in1_notify_r <= _GEN_625;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in1_notify_r <= _GEN_625;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_in1_notify_r <= _GEN_625;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_in1_notify_r <= _GEN_625;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_in1_notify_r <= _GEN_625;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in1_notify_r <= _GEN_720;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      slave_in1_notify_r <= 1'h0;
                                                                                                    end else begin
                                                                                                      slave_in1_notify_r <= _GEN_720;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_in1_notify_r <= _GEN_720;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_in1_notify_r <= _GEN_720;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in1_notify_r <= _GEN_720;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_in1_notify_r <= _GEN_720;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    slave_in1_notify_r <= 1'h0;
                                                                                                  end else begin
                                                                                                    slave_in1_notify_r <= _GEN_720;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_in1_notify_r <= _GEN_720;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in1_notify_r <= _GEN_720;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_in1_notify_r <= _GEN_720;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_in1_notify_r <= _GEN_720;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  slave_in1_notify_r <= 1'h0;
                                                                                                end else begin
                                                                                                  slave_in1_notify_r <= _GEN_720;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in1_notify_r <= _GEN_720;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_in1_notify_r <= _GEN_720;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_in1_notify_r <= _GEN_720;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_in1_notify_r <= _GEN_720;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in1_notify_r <= _GEN_815;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            slave_in1_notify_r <= 1'h0;
                                                                                          end else begin
                                                                                            slave_in1_notify_r <= _GEN_815;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_in1_notify_r <= _GEN_815;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_in1_notify_r <= _GEN_815;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in1_notify_r <= _GEN_815;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_in1_notify_r <= _GEN_815;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          slave_in1_notify_r <= 1'h0;
                                                                                        end else begin
                                                                                          slave_in1_notify_r <= _GEN_815;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_in1_notify_r <= _GEN_815;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in1_notify_r <= _GEN_815;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_in1_notify_r <= _GEN_815;
                                                                                  end
                                                                                end else begin
                                                                                  slave_in1_notify_r <= _GEN_815;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        slave_in1_notify_r <= 1'h0;
                                                                                      end else begin
                                                                                        slave_in1_notify_r <= _GEN_815;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in1_notify_r <= _GEN_815;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_in1_notify_r <= _GEN_815;
                                                                                  end
                                                                                end else begin
                                                                                  slave_in1_notify_r <= _GEN_815;
                                                                                end
                                                                              end else begin
                                                                                slave_in1_notify_r <= _GEN_815;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            slave_in1_notify_r <= _GEN_910;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_in1_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_in1_notify_r <= _GEN_910;
                                                                                end
                                                                              end else begin
                                                                                slave_in1_notify_r <= _GEN_910;
                                                                              end
                                                                            end else begin
                                                                              slave_in1_notify_r <= _GEN_910;
                                                                            end
                                                                          end else begin
                                                                            slave_in1_notify_r <= _GEN_910;
                                                                          end
                                                                        end else begin
                                                                          slave_in1_notify_r <= _GEN_910;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_in1_notify_r <= 1'h0;
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_in1_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_in1_notify_r <= _GEN_910;
                                                                                end
                                                                              end else begin
                                                                                slave_in1_notify_r <= _GEN_910;
                                                                              end
                                                                            end else begin
                                                                              slave_in1_notify_r <= _GEN_910;
                                                                            end
                                                                          end else begin
                                                                            slave_in1_notify_r <= _GEN_910;
                                                                          end
                                                                        end else begin
                                                                          slave_in1_notify_r <= _GEN_910;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                slave_in1_notify_r <= 1'h0;
                                                                              end else begin
                                                                                slave_in1_notify_r <= _GEN_910;
                                                                              end
                                                                            end else begin
                                                                              slave_in1_notify_r <= _GEN_910;
                                                                            end
                                                                          end else begin
                                                                            slave_in1_notify_r <= _GEN_910;
                                                                          end
                                                                        end else begin
                                                                          slave_in1_notify_r <= _GEN_910;
                                                                        end
                                                                      end else begin
                                                                        slave_in1_notify_r <= _GEN_910;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (io_slave_out0_sync) begin
                                                                      slave_in1_notify_r <= 1'h0;
                                                                    end else begin
                                                                      slave_in1_notify_r <= _GEN_1005;
                                                                    end
                                                                  end else begin
                                                                    slave_in1_notify_r <= _GEN_1005;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_in1_notify_r <= 1'h0;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_in1_notify_r <= 1'h0;
                                                                      end else begin
                                                                        slave_in1_notify_r <= _GEN_1005;
                                                                      end
                                                                    end else begin
                                                                      slave_in1_notify_r <= _GEN_1005;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  slave_in1_notify_r <= _GEN_1037;
                                                                end
                                                              end else begin
                                                                slave_in1_notify_r <= _GEN_1037;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  slave_in1_notify_r <= 1'h0;
                                                                end else begin
                                                                  slave_in1_notify_r <= _GEN_1037;
                                                                end
                                                              end else begin
                                                                slave_in1_notify_r <= _GEN_1037;
                                                              end
                                                            end else begin
                                                              slave_in1_notify_r <= _GEN_1037;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_in1_notify_r <= 1'h0;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_in1_notify_r <= 1'h0;
                                                                  end else begin
                                                                    slave_in1_notify_r <= _GEN_1037;
                                                                  end
                                                                end else begin
                                                                  slave_in1_notify_r <= _GEN_1037;
                                                                end
                                                              end else begin
                                                                slave_in1_notify_r <= _GEN_1037;
                                                              end
                                                            end
                                                          end else begin
                                                            slave_in1_notify_r <= _GEN_1091;
                                                          end
                                                        end else begin
                                                          slave_in1_notify_r <= _GEN_1091;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_in1_notify_r <= 1'h0;
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_in1_notify_r <= 1'h0;
                                                            end else begin
                                                              slave_in1_notify_r <= _GEN_1091;
                                                            end
                                                          end else begin
                                                            slave_in1_notify_r <= _GEN_1091;
                                                          end
                                                        end else begin
                                                          slave_in1_notify_r <= _GEN_1091;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            slave_in1_notify_r <= 1'h0;
                                                          end else begin
                                                            slave_in1_notify_r <= _GEN_1091;
                                                          end
                                                        end else begin
                                                          slave_in1_notify_r <= _GEN_1091;
                                                        end
                                                      end else begin
                                                        slave_in1_notify_r <= _GEN_1091;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_in1_notify_r <= 1'h1;
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_in1_notify_r <= 1'h0;
                                                      end else begin
                                                        slave_in1_notify_r <= _GEN_1145;
                                                      end
                                                    end else begin
                                                      slave_in1_notify_r <= _GEN_1145;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (io_master_out_sync) begin
                                                      slave_in1_notify_r <= 1'h0;
                                                    end else begin
                                                      slave_in1_notify_r <= _GEN_1145;
                                                    end
                                                  end else begin
                                                    slave_in1_notify_r <= _GEN_1145;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (io_slave_out1_sync) begin
                                                  slave_in1_notify_r <= 1'h1;
                                                end else begin
                                                  slave_in1_notify_r <= _GEN_1177;
                                                end
                                              end else begin
                                                slave_in1_notify_r <= _GEN_1177;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_in1_notify_r <= 1'h0;
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_in1_notify_r <= 1'h1;
                                                  end else begin
                                                    slave_in1_notify_r <= _GEN_1177;
                                                  end
                                                end else begin
                                                  slave_in1_notify_r <= _GEN_1177;
                                                end
                                              end
                                            end else begin
                                              slave_in1_notify_r <= _GEN_1209;
                                            end
                                          end else begin
                                            slave_in1_notify_r <= _GEN_1209;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              slave_in1_notify_r <= 1'h0;
                                            end else begin
                                              slave_in1_notify_r <= _GEN_1209;
                                            end
                                          end else begin
                                            slave_in1_notify_r <= _GEN_1209;
                                          end
                                        end else begin
                                          slave_in1_notify_r <= _GEN_1209;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_in1_notify_r <= 1'h0;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_in1_notify_r <= 1'h0;
                                              end else begin
                                                slave_in1_notify_r <= _GEN_1209;
                                              end
                                            end else begin
                                              slave_in1_notify_r <= _GEN_1209;
                                            end
                                          end else begin
                                            slave_in1_notify_r <= _GEN_1209;
                                          end
                                        end
                                      end else begin
                                        slave_in1_notify_r <= _GEN_1263;
                                      end
                                    end else begin
                                      slave_in1_notify_r <= _GEN_1263;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_in1_notify_r <= 1'h0;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_in1_notify_r <= 1'h0;
                                        end else begin
                                          slave_in1_notify_r <= _GEN_1263;
                                        end
                                      end else begin
                                        slave_in1_notify_r <= _GEN_1263;
                                      end
                                    end else begin
                                      slave_in1_notify_r <= _GEN_1263;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        slave_in1_notify_r <= 1'h0;
                                      end else begin
                                        slave_in1_notify_r <= _GEN_1263;
                                      end
                                    end else begin
                                      slave_in1_notify_r <= _GEN_1263;
                                    end
                                  end else begin
                                    slave_in1_notify_r <= _GEN_1263;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (io_slave_out2_sync) begin
                                  slave_in1_notify_r <= 1'h0;
                                end else begin
                                  slave_in1_notify_r <= _GEN_1317;
                                end
                              end else begin
                                slave_in1_notify_r <= _GEN_1317;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_in1_notify_r <= 1'h0;
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_in1_notify_r <= 1'h0;
                                  end else begin
                                    slave_in1_notify_r <= _GEN_1317;
                                  end
                                end else begin
                                  slave_in1_notify_r <= _GEN_1317;
                                end
                              end
                            end else begin
                              slave_in1_notify_r <= _GEN_1349;
                            end
                          end else begin
                            slave_in1_notify_r <= _GEN_1349;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              slave_in1_notify_r <= 1'h0;
                            end else begin
                              slave_in1_notify_r <= _GEN_1349;
                            end
                          end else begin
                            slave_in1_notify_r <= _GEN_1349;
                          end
                        end else begin
                          slave_in1_notify_r <= _GEN_1349;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_in1_notify_r <= 1'h0;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_in1_notify_r <= 1'h0;
                              end else begin
                                slave_in1_notify_r <= _GEN_1349;
                              end
                            end else begin
                              slave_in1_notify_r <= _GEN_1349;
                            end
                          end else begin
                            slave_in1_notify_r <= _GEN_1349;
                          end
                        end
                      end else begin
                        slave_in1_notify_r <= _GEN_1403;
                      end
                    end else begin
                      slave_in1_notify_r <= _GEN_1403;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_in1_notify_r <= 1'h0;
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_in1_notify_r <= 1'h0;
                        end else begin
                          slave_in1_notify_r <= _GEN_1403;
                        end
                      end else begin
                        slave_in1_notify_r <= _GEN_1403;
                      end
                    end else begin
                      slave_in1_notify_r <= _GEN_1403;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        slave_in1_notify_r <= 1'h0;
                      end else begin
                        slave_in1_notify_r <= _GEN_1403;
                      end
                    end else begin
                      slave_in1_notify_r <= _GEN_1403;
                    end
                  end else begin
                    slave_in1_notify_r <= _GEN_1403;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (io_slave_out3_sync) begin
                  slave_in1_notify_r <= 1'h0;
                end else begin
                  slave_in1_notify_r <= _GEN_1457;
                end
              end else begin
                slave_in1_notify_r <= _GEN_1457;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                slave_in1_notify_r <= 1'h0;
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_in1_notify_r <= 1'h0;
                  end else begin
                    slave_in1_notify_r <= _GEN_1457;
                  end
                end else begin
                  slave_in1_notify_r <= _GEN_1457;
                end
              end
            end else begin
              slave_in1_notify_r <= _GEN_1489;
            end
          end else begin
            slave_in1_notify_r <= _GEN_1489;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              slave_in1_notify_r <= 1'h0;
            end else begin
              slave_in1_notify_r <= _GEN_1489;
            end
          end else begin
            slave_in1_notify_r <= _GEN_1489;
          end
        end else begin
          slave_in1_notify_r <= _GEN_1489;
        end
      end
    end
    if (reset) begin
      slave_in2_notify_r <= 1'h0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            slave_in2_notify_r <= 1'h0;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  slave_in2_notify_r <= 1'h0;
                end else begin
                  if (_T_518) begin
                    if (io_slave_out3_sync) begin
                      slave_in2_notify_r <= 1'h0;
                    end else begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            slave_in2_notify_r <= 1'h0;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  slave_in2_notify_r <= 1'h0;
                                end else begin
                                  if (_T_479) begin
                                    if (io_slave_out2_sync) begin
                                      slave_in2_notify_r <= 1'h1;
                                    end else begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            slave_in2_notify_r <= 1'h0;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  slave_in2_notify_r <= 1'h0;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (io_slave_out1_sync) begin
                                                      slave_in2_notify_r <= 1'h0;
                                                    end else begin
                                                      if (_T_429) begin
                                                        if (io_master_out_sync) begin
                                                          slave_in2_notify_r <= 1'h0;
                                                        end else begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                slave_in2_notify_r <= 1'h0;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      slave_in2_notify_r <= 1'h0;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (io_slave_out0_sync) begin
                                                                          slave_in2_notify_r <= 1'h0;
                                                                        end else begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    slave_in2_notify_r <= 1'h0;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              slave_in2_notify_r <= 1'h0;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        slave_in2_notify_r <= 1'h0;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  slave_in2_notify_r <= 1'h0;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            slave_in2_notify_r <= 1'h0;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      slave_in2_notify_r <= 1'h0;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    slave_in2_notify_r <= 1'h0;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  slave_in2_notify_r <= 1'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            slave_in2_notify_r <= 1'h0;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      slave_in2_notify_r <= 1'h0;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    slave_in2_notify_r <= 1'h0;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  slave_in2_notify_r <= 1'h0;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                slave_in2_notify_r <= 1'h0;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          slave_in2_notify_r <= 1'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                          slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        slave_in2_notify_r <= 1'h0;
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_in2_notify_r <= _GEN_89;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      slave_in2_notify_r <= 1'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_in2_notify_r <= _GEN_89;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_in2_notify_r <= _GEN_89;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_in2_notify_r <= _GEN_89;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in2_notify_r <= _GEN_184;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in2_notify_r <= _GEN_184;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in2_notify_r <= _GEN_184;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                slave_in2_notify_r <= 1'h0;
                                                                                                                                                              end else begin
                                                                                                                                                                slave_in2_notify_r <= _GEN_184;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_in2_notify_r <= _GEN_184;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_in2_notify_r <= _GEN_184;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in2_notify_r <= _GEN_184;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in2_notify_r <= _GEN_184;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in2_notify_r <= _GEN_184;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_in2_notify_r <= _GEN_184;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              slave_in2_notify_r <= 1'h0;
                                                                                                                                                            end else begin
                                                                                                                                                              slave_in2_notify_r <= _GEN_184;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_in2_notify_r <= _GEN_184;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in2_notify_r <= _GEN_184;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in2_notify_r <= _GEN_184;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in2_notify_r <= _GEN_184;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_in2_notify_r <= _GEN_184;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_in2_notify_r <= _GEN_184;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            slave_in2_notify_r <= 1'h0;
                                                                                                                                                          end else begin
                                                                                                                                                            slave_in2_notify_r <= _GEN_184;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in2_notify_r <= _GEN_184;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in2_notify_r <= _GEN_184;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in2_notify_r <= _GEN_184;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_in2_notify_r <= _GEN_184;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_in2_notify_r <= _GEN_184;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_in2_notify_r <= _GEN_184;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in2_notify_r <= _GEN_310;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in2_notify_r <= _GEN_310;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in2_notify_r <= _GEN_310;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  slave_in2_notify_r <= 1'h0;
                                                                                                                                                end else begin
                                                                                                                                                  slave_in2_notify_r <= _GEN_310;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_in2_notify_r <= _GEN_310;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_in2_notify_r <= _GEN_310;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in2_notify_r <= _GEN_310;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in2_notify_r <= _GEN_310;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in2_notify_r <= _GEN_310;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_in2_notify_r <= _GEN_310;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                slave_in2_notify_r <= 1'h0;
                                                                                                                                              end else begin
                                                                                                                                                slave_in2_notify_r <= _GEN_310;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_in2_notify_r <= _GEN_310;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in2_notify_r <= _GEN_310;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in2_notify_r <= _GEN_310;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in2_notify_r <= _GEN_310;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_in2_notify_r <= _GEN_310;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_in2_notify_r <= _GEN_310;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              slave_in2_notify_r <= 1'h0;
                                                                                                                                            end else begin
                                                                                                                                              slave_in2_notify_r <= _GEN_310;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in2_notify_r <= _GEN_310;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in2_notify_r <= _GEN_310;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in2_notify_r <= _GEN_310;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_in2_notify_r <= _GEN_310;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_in2_notify_r <= _GEN_310;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_in2_notify_r <= _GEN_310;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in2_notify_r <= _GEN_436;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    slave_in2_notify_r <= 1'h0;
                                                                                                                                  end else begin
                                                                                                                                    slave_in2_notify_r <= _GEN_436;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_in2_notify_r <= _GEN_436;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_in2_notify_r <= _GEN_436;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in2_notify_r <= _GEN_436;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_in2_notify_r <= _GEN_436;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  slave_in2_notify_r <= 1'h0;
                                                                                                                                end else begin
                                                                                                                                  slave_in2_notify_r <= _GEN_436;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_in2_notify_r <= _GEN_436;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in2_notify_r <= _GEN_436;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_in2_notify_r <= _GEN_436;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_in2_notify_r <= _GEN_436;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                slave_in2_notify_r <= 1'h0;
                                                                                                                              end else begin
                                                                                                                                slave_in2_notify_r <= _GEN_436;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in2_notify_r <= _GEN_436;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_in2_notify_r <= _GEN_436;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_in2_notify_r <= _GEN_436;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_in2_notify_r <= _GEN_436;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in2_notify_r <= _GEN_531;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          slave_in2_notify_r <= 1'h0;
                                                                                                                        end else begin
                                                                                                                          slave_in2_notify_r <= _GEN_531;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_in2_notify_r <= _GEN_531;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_in2_notify_r <= _GEN_531;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in2_notify_r <= _GEN_531;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_in2_notify_r <= _GEN_531;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        slave_in2_notify_r <= 1'h0;
                                                                                                                      end else begin
                                                                                                                        slave_in2_notify_r <= _GEN_531;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_in2_notify_r <= _GEN_531;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in2_notify_r <= _GEN_531;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_in2_notify_r <= _GEN_531;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_in2_notify_r <= _GEN_531;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      slave_in2_notify_r <= 1'h0;
                                                                                                                    end else begin
                                                                                                                      slave_in2_notify_r <= _GEN_531;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in2_notify_r <= _GEN_531;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_in2_notify_r <= _GEN_531;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_in2_notify_r <= _GEN_531;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_in2_notify_r <= _GEN_531;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in2_notify_r <= _GEN_626;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                slave_in2_notify_r <= 1'h0;
                                                                                                              end else begin
                                                                                                                slave_in2_notify_r <= _GEN_626;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_in2_notify_r <= _GEN_626;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_in2_notify_r <= _GEN_626;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in2_notify_r <= _GEN_626;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_in2_notify_r <= _GEN_626;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              slave_in2_notify_r <= 1'h0;
                                                                                                            end else begin
                                                                                                              slave_in2_notify_r <= _GEN_626;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_in2_notify_r <= _GEN_626;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in2_notify_r <= _GEN_626;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_in2_notify_r <= _GEN_626;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_in2_notify_r <= _GEN_626;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            slave_in2_notify_r <= 1'h0;
                                                                                                          end else begin
                                                                                                            slave_in2_notify_r <= _GEN_626;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in2_notify_r <= _GEN_626;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_in2_notify_r <= _GEN_626;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_in2_notify_r <= _GEN_626;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_in2_notify_r <= _GEN_626;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in2_notify_r <= _GEN_721;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      slave_in2_notify_r <= 1'h0;
                                                                                                    end else begin
                                                                                                      slave_in2_notify_r <= _GEN_721;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_in2_notify_r <= _GEN_721;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_in2_notify_r <= _GEN_721;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in2_notify_r <= _GEN_721;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_in2_notify_r <= _GEN_721;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    slave_in2_notify_r <= 1'h0;
                                                                                                  end else begin
                                                                                                    slave_in2_notify_r <= _GEN_721;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_in2_notify_r <= _GEN_721;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in2_notify_r <= _GEN_721;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_in2_notify_r <= _GEN_721;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_in2_notify_r <= _GEN_721;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  slave_in2_notify_r <= 1'h0;
                                                                                                end else begin
                                                                                                  slave_in2_notify_r <= _GEN_721;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in2_notify_r <= _GEN_721;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_in2_notify_r <= _GEN_721;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_in2_notify_r <= _GEN_721;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_in2_notify_r <= _GEN_721;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in2_notify_r <= _GEN_816;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            slave_in2_notify_r <= 1'h0;
                                                                                          end else begin
                                                                                            slave_in2_notify_r <= _GEN_816;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_in2_notify_r <= _GEN_816;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_in2_notify_r <= _GEN_816;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in2_notify_r <= _GEN_816;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_in2_notify_r <= _GEN_816;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          slave_in2_notify_r <= 1'h0;
                                                                                        end else begin
                                                                                          slave_in2_notify_r <= _GEN_816;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_in2_notify_r <= _GEN_816;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in2_notify_r <= _GEN_816;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_in2_notify_r <= _GEN_816;
                                                                                  end
                                                                                end else begin
                                                                                  slave_in2_notify_r <= _GEN_816;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        slave_in2_notify_r <= 1'h0;
                                                                                      end else begin
                                                                                        slave_in2_notify_r <= _GEN_816;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in2_notify_r <= _GEN_816;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_in2_notify_r <= _GEN_816;
                                                                                  end
                                                                                end else begin
                                                                                  slave_in2_notify_r <= _GEN_816;
                                                                                end
                                                                              end else begin
                                                                                slave_in2_notify_r <= _GEN_816;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            slave_in2_notify_r <= _GEN_911;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_in2_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_in2_notify_r <= _GEN_911;
                                                                                end
                                                                              end else begin
                                                                                slave_in2_notify_r <= _GEN_911;
                                                                              end
                                                                            end else begin
                                                                              slave_in2_notify_r <= _GEN_911;
                                                                            end
                                                                          end else begin
                                                                            slave_in2_notify_r <= _GEN_911;
                                                                          end
                                                                        end else begin
                                                                          slave_in2_notify_r <= _GEN_911;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_in2_notify_r <= 1'h0;
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_in2_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_in2_notify_r <= _GEN_911;
                                                                                end
                                                                              end else begin
                                                                                slave_in2_notify_r <= _GEN_911;
                                                                              end
                                                                            end else begin
                                                                              slave_in2_notify_r <= _GEN_911;
                                                                            end
                                                                          end else begin
                                                                            slave_in2_notify_r <= _GEN_911;
                                                                          end
                                                                        end else begin
                                                                          slave_in2_notify_r <= _GEN_911;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                slave_in2_notify_r <= 1'h0;
                                                                              end else begin
                                                                                slave_in2_notify_r <= _GEN_911;
                                                                              end
                                                                            end else begin
                                                                              slave_in2_notify_r <= _GEN_911;
                                                                            end
                                                                          end else begin
                                                                            slave_in2_notify_r <= _GEN_911;
                                                                          end
                                                                        end else begin
                                                                          slave_in2_notify_r <= _GEN_911;
                                                                        end
                                                                      end else begin
                                                                        slave_in2_notify_r <= _GEN_911;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (io_slave_out0_sync) begin
                                                                      slave_in2_notify_r <= 1'h0;
                                                                    end else begin
                                                                      slave_in2_notify_r <= _GEN_1006;
                                                                    end
                                                                  end else begin
                                                                    slave_in2_notify_r <= _GEN_1006;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_in2_notify_r <= 1'h0;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_in2_notify_r <= 1'h0;
                                                                      end else begin
                                                                        slave_in2_notify_r <= _GEN_1006;
                                                                      end
                                                                    end else begin
                                                                      slave_in2_notify_r <= _GEN_1006;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  slave_in2_notify_r <= _GEN_1038;
                                                                end
                                                              end else begin
                                                                slave_in2_notify_r <= _GEN_1038;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  slave_in2_notify_r <= 1'h0;
                                                                end else begin
                                                                  slave_in2_notify_r <= _GEN_1038;
                                                                end
                                                              end else begin
                                                                slave_in2_notify_r <= _GEN_1038;
                                                              end
                                                            end else begin
                                                              slave_in2_notify_r <= _GEN_1038;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_in2_notify_r <= 1'h0;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_in2_notify_r <= 1'h0;
                                                                  end else begin
                                                                    slave_in2_notify_r <= _GEN_1038;
                                                                  end
                                                                end else begin
                                                                  slave_in2_notify_r <= _GEN_1038;
                                                                end
                                                              end else begin
                                                                slave_in2_notify_r <= _GEN_1038;
                                                              end
                                                            end
                                                          end else begin
                                                            slave_in2_notify_r <= _GEN_1092;
                                                          end
                                                        end else begin
                                                          slave_in2_notify_r <= _GEN_1092;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_in2_notify_r <= 1'h0;
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_in2_notify_r <= 1'h0;
                                                            end else begin
                                                              slave_in2_notify_r <= _GEN_1092;
                                                            end
                                                          end else begin
                                                            slave_in2_notify_r <= _GEN_1092;
                                                          end
                                                        end else begin
                                                          slave_in2_notify_r <= _GEN_1092;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            slave_in2_notify_r <= 1'h0;
                                                          end else begin
                                                            slave_in2_notify_r <= _GEN_1092;
                                                          end
                                                        end else begin
                                                          slave_in2_notify_r <= _GEN_1092;
                                                        end
                                                      end else begin
                                                        slave_in2_notify_r <= _GEN_1092;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_in2_notify_r <= 1'h0;
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_in2_notify_r <= 1'h0;
                                                      end else begin
                                                        slave_in2_notify_r <= _GEN_1146;
                                                      end
                                                    end else begin
                                                      slave_in2_notify_r <= _GEN_1146;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (io_master_out_sync) begin
                                                      slave_in2_notify_r <= 1'h0;
                                                    end else begin
                                                      slave_in2_notify_r <= _GEN_1146;
                                                    end
                                                  end else begin
                                                    slave_in2_notify_r <= _GEN_1146;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (io_slave_out1_sync) begin
                                                  slave_in2_notify_r <= 1'h0;
                                                end else begin
                                                  slave_in2_notify_r <= _GEN_1178;
                                                end
                                              end else begin
                                                slave_in2_notify_r <= _GEN_1178;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_in2_notify_r <= 1'h0;
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_in2_notify_r <= 1'h0;
                                                  end else begin
                                                    slave_in2_notify_r <= _GEN_1178;
                                                  end
                                                end else begin
                                                  slave_in2_notify_r <= _GEN_1178;
                                                end
                                              end
                                            end else begin
                                              slave_in2_notify_r <= _GEN_1210;
                                            end
                                          end else begin
                                            slave_in2_notify_r <= _GEN_1210;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              slave_in2_notify_r <= 1'h0;
                                            end else begin
                                              slave_in2_notify_r <= _GEN_1210;
                                            end
                                          end else begin
                                            slave_in2_notify_r <= _GEN_1210;
                                          end
                                        end else begin
                                          slave_in2_notify_r <= _GEN_1210;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_in2_notify_r <= 1'h0;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_in2_notify_r <= 1'h0;
                                              end else begin
                                                slave_in2_notify_r <= _GEN_1210;
                                              end
                                            end else begin
                                              slave_in2_notify_r <= _GEN_1210;
                                            end
                                          end else begin
                                            slave_in2_notify_r <= _GEN_1210;
                                          end
                                        end
                                      end else begin
                                        slave_in2_notify_r <= _GEN_1264;
                                      end
                                    end else begin
                                      slave_in2_notify_r <= _GEN_1264;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_in2_notify_r <= 1'h1;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_in2_notify_r <= 1'h0;
                                        end else begin
                                          slave_in2_notify_r <= _GEN_1264;
                                        end
                                      end else begin
                                        slave_in2_notify_r <= _GEN_1264;
                                      end
                                    end else begin
                                      slave_in2_notify_r <= _GEN_1264;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        slave_in2_notify_r <= 1'h0;
                                      end else begin
                                        slave_in2_notify_r <= _GEN_1264;
                                      end
                                    end else begin
                                      slave_in2_notify_r <= _GEN_1264;
                                    end
                                  end else begin
                                    slave_in2_notify_r <= _GEN_1264;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (io_slave_out2_sync) begin
                                  slave_in2_notify_r <= 1'h1;
                                end else begin
                                  slave_in2_notify_r <= _GEN_1318;
                                end
                              end else begin
                                slave_in2_notify_r <= _GEN_1318;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_in2_notify_r <= 1'h0;
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_in2_notify_r <= 1'h1;
                                  end else begin
                                    slave_in2_notify_r <= _GEN_1318;
                                  end
                                end else begin
                                  slave_in2_notify_r <= _GEN_1318;
                                end
                              end
                            end else begin
                              slave_in2_notify_r <= _GEN_1350;
                            end
                          end else begin
                            slave_in2_notify_r <= _GEN_1350;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              slave_in2_notify_r <= 1'h0;
                            end else begin
                              slave_in2_notify_r <= _GEN_1350;
                            end
                          end else begin
                            slave_in2_notify_r <= _GEN_1350;
                          end
                        end else begin
                          slave_in2_notify_r <= _GEN_1350;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_in2_notify_r <= 1'h0;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_in2_notify_r <= 1'h0;
                              end else begin
                                slave_in2_notify_r <= _GEN_1350;
                              end
                            end else begin
                              slave_in2_notify_r <= _GEN_1350;
                            end
                          end else begin
                            slave_in2_notify_r <= _GEN_1350;
                          end
                        end
                      end else begin
                        slave_in2_notify_r <= _GEN_1404;
                      end
                    end else begin
                      slave_in2_notify_r <= _GEN_1404;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_in2_notify_r <= 1'h0;
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_in2_notify_r <= 1'h0;
                        end else begin
                          slave_in2_notify_r <= _GEN_1404;
                        end
                      end else begin
                        slave_in2_notify_r <= _GEN_1404;
                      end
                    end else begin
                      slave_in2_notify_r <= _GEN_1404;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        slave_in2_notify_r <= 1'h0;
                      end else begin
                        slave_in2_notify_r <= _GEN_1404;
                      end
                    end else begin
                      slave_in2_notify_r <= _GEN_1404;
                    end
                  end else begin
                    slave_in2_notify_r <= _GEN_1404;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (io_slave_out3_sync) begin
                  slave_in2_notify_r <= 1'h0;
                end else begin
                  slave_in2_notify_r <= _GEN_1458;
                end
              end else begin
                slave_in2_notify_r <= _GEN_1458;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                slave_in2_notify_r <= 1'h0;
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_in2_notify_r <= 1'h0;
                  end else begin
                    slave_in2_notify_r <= _GEN_1458;
                  end
                end else begin
                  slave_in2_notify_r <= _GEN_1458;
                end
              end
            end else begin
              slave_in2_notify_r <= _GEN_1490;
            end
          end else begin
            slave_in2_notify_r <= _GEN_1490;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              slave_in2_notify_r <= 1'h0;
            end else begin
              slave_in2_notify_r <= _GEN_1490;
            end
          end else begin
            slave_in2_notify_r <= _GEN_1490;
          end
        end else begin
          slave_in2_notify_r <= _GEN_1490;
        end
      end
    end
    if (reset) begin
      slave_in3_notify_r <= 1'h0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            slave_in3_notify_r <= 1'h0;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  slave_in3_notify_r <= 1'h0;
                end else begin
                  if (_T_518) begin
                    if (io_slave_out3_sync) begin
                      slave_in3_notify_r <= 1'h1;
                    end else begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            slave_in3_notify_r <= 1'h0;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  slave_in3_notify_r <= 1'h0;
                                end else begin
                                  if (_T_479) begin
                                    if (io_slave_out2_sync) begin
                                      slave_in3_notify_r <= 1'h0;
                                    end else begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            slave_in3_notify_r <= 1'h0;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  slave_in3_notify_r <= 1'h0;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (io_slave_out1_sync) begin
                                                      slave_in3_notify_r <= 1'h0;
                                                    end else begin
                                                      if (_T_429) begin
                                                        if (io_master_out_sync) begin
                                                          slave_in3_notify_r <= 1'h0;
                                                        end else begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                slave_in3_notify_r <= 1'h0;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      slave_in3_notify_r <= 1'h0;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (io_slave_out0_sync) begin
                                                                          slave_in3_notify_r <= 1'h0;
                                                                        end else begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    slave_in3_notify_r <= 1'h0;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              slave_in3_notify_r <= 1'h0;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        slave_in3_notify_r <= 1'h0;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  slave_in3_notify_r <= 1'h0;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            slave_in3_notify_r <= 1'h0;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      slave_in3_notify_r <= 1'h0;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    slave_in3_notify_r <= 1'h0;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  slave_in3_notify_r <= 1'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            slave_in3_notify_r <= 1'h0;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      slave_in3_notify_r <= 1'h0;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    slave_in3_notify_r <= 1'h0;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  slave_in3_notify_r <= 1'h0;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                slave_in3_notify_r <= 1'h0;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          slave_in3_notify_r <= 1'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                          slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        slave_in3_notify_r <= 1'h0;
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_in3_notify_r <= _GEN_90;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      slave_in3_notify_r <= 1'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_in3_notify_r <= _GEN_90;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_in3_notify_r <= _GEN_90;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_in3_notify_r <= _GEN_90;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in3_notify_r <= _GEN_185;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in3_notify_r <= _GEN_185;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in3_notify_r <= _GEN_185;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                slave_in3_notify_r <= 1'h0;
                                                                                                                                                              end else begin
                                                                                                                                                                slave_in3_notify_r <= _GEN_185;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_in3_notify_r <= _GEN_185;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_in3_notify_r <= _GEN_185;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in3_notify_r <= _GEN_185;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in3_notify_r <= _GEN_185;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in3_notify_r <= _GEN_185;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_in3_notify_r <= _GEN_185;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              slave_in3_notify_r <= 1'h0;
                                                                                                                                                            end else begin
                                                                                                                                                              slave_in3_notify_r <= _GEN_185;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_in3_notify_r <= _GEN_185;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in3_notify_r <= _GEN_185;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in3_notify_r <= _GEN_185;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in3_notify_r <= _GEN_185;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_in3_notify_r <= _GEN_185;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_in3_notify_r <= _GEN_185;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            slave_in3_notify_r <= 1'h0;
                                                                                                                                                          end else begin
                                                                                                                                                            slave_in3_notify_r <= _GEN_185;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_in3_notify_r <= _GEN_185;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_in3_notify_r <= _GEN_185;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_in3_notify_r <= _GEN_185;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_in3_notify_r <= _GEN_185;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_in3_notify_r <= _GEN_185;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_in3_notify_r <= _GEN_185;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in3_notify_r <= _GEN_311;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in3_notify_r <= _GEN_311;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in3_notify_r <= _GEN_311;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  slave_in3_notify_r <= 1'h0;
                                                                                                                                                end else begin
                                                                                                                                                  slave_in3_notify_r <= _GEN_311;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_in3_notify_r <= _GEN_311;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_in3_notify_r <= _GEN_311;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in3_notify_r <= _GEN_311;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in3_notify_r <= _GEN_311;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in3_notify_r <= _GEN_311;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_in3_notify_r <= _GEN_311;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                slave_in3_notify_r <= 1'h0;
                                                                                                                                              end else begin
                                                                                                                                                slave_in3_notify_r <= _GEN_311;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_in3_notify_r <= _GEN_311;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in3_notify_r <= _GEN_311;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in3_notify_r <= _GEN_311;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in3_notify_r <= _GEN_311;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_in3_notify_r <= _GEN_311;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_in3_notify_r <= _GEN_311;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              slave_in3_notify_r <= 1'h0;
                                                                                                                                            end else begin
                                                                                                                                              slave_in3_notify_r <= _GEN_311;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_in3_notify_r <= _GEN_311;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_in3_notify_r <= _GEN_311;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_in3_notify_r <= _GEN_311;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_in3_notify_r <= _GEN_311;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_in3_notify_r <= _GEN_311;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_in3_notify_r <= _GEN_311;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in3_notify_r <= _GEN_437;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    slave_in3_notify_r <= 1'h0;
                                                                                                                                  end else begin
                                                                                                                                    slave_in3_notify_r <= _GEN_437;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_in3_notify_r <= _GEN_437;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_in3_notify_r <= _GEN_437;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in3_notify_r <= _GEN_437;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_in3_notify_r <= _GEN_437;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  slave_in3_notify_r <= 1'h0;
                                                                                                                                end else begin
                                                                                                                                  slave_in3_notify_r <= _GEN_437;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_in3_notify_r <= _GEN_437;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in3_notify_r <= _GEN_437;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_in3_notify_r <= _GEN_437;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_in3_notify_r <= _GEN_437;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                slave_in3_notify_r <= 1'h0;
                                                                                                                              end else begin
                                                                                                                                slave_in3_notify_r <= _GEN_437;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_in3_notify_r <= _GEN_437;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_in3_notify_r <= _GEN_437;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_in3_notify_r <= _GEN_437;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_in3_notify_r <= _GEN_437;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in3_notify_r <= _GEN_532;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          slave_in3_notify_r <= 1'h0;
                                                                                                                        end else begin
                                                                                                                          slave_in3_notify_r <= _GEN_532;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_in3_notify_r <= _GEN_532;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_in3_notify_r <= _GEN_532;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in3_notify_r <= _GEN_532;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_in3_notify_r <= _GEN_532;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        slave_in3_notify_r <= 1'h0;
                                                                                                                      end else begin
                                                                                                                        slave_in3_notify_r <= _GEN_532;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_in3_notify_r <= _GEN_532;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in3_notify_r <= _GEN_532;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_in3_notify_r <= _GEN_532;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_in3_notify_r <= _GEN_532;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      slave_in3_notify_r <= 1'h0;
                                                                                                                    end else begin
                                                                                                                      slave_in3_notify_r <= _GEN_532;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_in3_notify_r <= _GEN_532;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_in3_notify_r <= _GEN_532;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_in3_notify_r <= _GEN_532;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_in3_notify_r <= _GEN_532;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in3_notify_r <= _GEN_627;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                slave_in3_notify_r <= 1'h0;
                                                                                                              end else begin
                                                                                                                slave_in3_notify_r <= _GEN_627;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_in3_notify_r <= _GEN_627;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_in3_notify_r <= _GEN_627;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in3_notify_r <= _GEN_627;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_in3_notify_r <= _GEN_627;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              slave_in3_notify_r <= 1'h0;
                                                                                                            end else begin
                                                                                                              slave_in3_notify_r <= _GEN_627;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_in3_notify_r <= _GEN_627;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in3_notify_r <= _GEN_627;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_in3_notify_r <= _GEN_627;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_in3_notify_r <= _GEN_627;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            slave_in3_notify_r <= 1'h0;
                                                                                                          end else begin
                                                                                                            slave_in3_notify_r <= _GEN_627;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_in3_notify_r <= _GEN_627;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_in3_notify_r <= _GEN_627;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_in3_notify_r <= _GEN_627;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_in3_notify_r <= _GEN_627;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in3_notify_r <= _GEN_722;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      slave_in3_notify_r <= 1'h0;
                                                                                                    end else begin
                                                                                                      slave_in3_notify_r <= _GEN_722;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_in3_notify_r <= _GEN_722;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_in3_notify_r <= _GEN_722;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in3_notify_r <= _GEN_722;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_in3_notify_r <= _GEN_722;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    slave_in3_notify_r <= 1'h0;
                                                                                                  end else begin
                                                                                                    slave_in3_notify_r <= _GEN_722;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_in3_notify_r <= _GEN_722;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in3_notify_r <= _GEN_722;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_in3_notify_r <= _GEN_722;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_in3_notify_r <= _GEN_722;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  slave_in3_notify_r <= 1'h0;
                                                                                                end else begin
                                                                                                  slave_in3_notify_r <= _GEN_722;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_in3_notify_r <= _GEN_722;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_in3_notify_r <= _GEN_722;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_in3_notify_r <= _GEN_722;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_in3_notify_r <= _GEN_722;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in3_notify_r <= _GEN_817;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            slave_in3_notify_r <= 1'h0;
                                                                                          end else begin
                                                                                            slave_in3_notify_r <= _GEN_817;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_in3_notify_r <= _GEN_817;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_in3_notify_r <= _GEN_817;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in3_notify_r <= _GEN_817;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_in3_notify_r <= _GEN_817;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          slave_in3_notify_r <= 1'h0;
                                                                                        end else begin
                                                                                          slave_in3_notify_r <= _GEN_817;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_in3_notify_r <= _GEN_817;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in3_notify_r <= _GEN_817;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_in3_notify_r <= _GEN_817;
                                                                                  end
                                                                                end else begin
                                                                                  slave_in3_notify_r <= _GEN_817;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        slave_in3_notify_r <= 1'h0;
                                                                                      end else begin
                                                                                        slave_in3_notify_r <= _GEN_817;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_in3_notify_r <= _GEN_817;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_in3_notify_r <= _GEN_817;
                                                                                  end
                                                                                end else begin
                                                                                  slave_in3_notify_r <= _GEN_817;
                                                                                end
                                                                              end else begin
                                                                                slave_in3_notify_r <= _GEN_817;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            slave_in3_notify_r <= _GEN_912;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_in3_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_in3_notify_r <= _GEN_912;
                                                                                end
                                                                              end else begin
                                                                                slave_in3_notify_r <= _GEN_912;
                                                                              end
                                                                            end else begin
                                                                              slave_in3_notify_r <= _GEN_912;
                                                                            end
                                                                          end else begin
                                                                            slave_in3_notify_r <= _GEN_912;
                                                                          end
                                                                        end else begin
                                                                          slave_in3_notify_r <= _GEN_912;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_in3_notify_r <= 1'h0;
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_in3_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_in3_notify_r <= _GEN_912;
                                                                                end
                                                                              end else begin
                                                                                slave_in3_notify_r <= _GEN_912;
                                                                              end
                                                                            end else begin
                                                                              slave_in3_notify_r <= _GEN_912;
                                                                            end
                                                                          end else begin
                                                                            slave_in3_notify_r <= _GEN_912;
                                                                          end
                                                                        end else begin
                                                                          slave_in3_notify_r <= _GEN_912;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                slave_in3_notify_r <= 1'h0;
                                                                              end else begin
                                                                                slave_in3_notify_r <= _GEN_912;
                                                                              end
                                                                            end else begin
                                                                              slave_in3_notify_r <= _GEN_912;
                                                                            end
                                                                          end else begin
                                                                            slave_in3_notify_r <= _GEN_912;
                                                                          end
                                                                        end else begin
                                                                          slave_in3_notify_r <= _GEN_912;
                                                                        end
                                                                      end else begin
                                                                        slave_in3_notify_r <= _GEN_912;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (io_slave_out0_sync) begin
                                                                      slave_in3_notify_r <= 1'h0;
                                                                    end else begin
                                                                      slave_in3_notify_r <= _GEN_1007;
                                                                    end
                                                                  end else begin
                                                                    slave_in3_notify_r <= _GEN_1007;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_in3_notify_r <= 1'h0;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_in3_notify_r <= 1'h0;
                                                                      end else begin
                                                                        slave_in3_notify_r <= _GEN_1007;
                                                                      end
                                                                    end else begin
                                                                      slave_in3_notify_r <= _GEN_1007;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  slave_in3_notify_r <= _GEN_1039;
                                                                end
                                                              end else begin
                                                                slave_in3_notify_r <= _GEN_1039;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  slave_in3_notify_r <= 1'h0;
                                                                end else begin
                                                                  slave_in3_notify_r <= _GEN_1039;
                                                                end
                                                              end else begin
                                                                slave_in3_notify_r <= _GEN_1039;
                                                              end
                                                            end else begin
                                                              slave_in3_notify_r <= _GEN_1039;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_in3_notify_r <= 1'h0;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_in3_notify_r <= 1'h0;
                                                                  end else begin
                                                                    slave_in3_notify_r <= _GEN_1039;
                                                                  end
                                                                end else begin
                                                                  slave_in3_notify_r <= _GEN_1039;
                                                                end
                                                              end else begin
                                                                slave_in3_notify_r <= _GEN_1039;
                                                              end
                                                            end
                                                          end else begin
                                                            slave_in3_notify_r <= _GEN_1093;
                                                          end
                                                        end else begin
                                                          slave_in3_notify_r <= _GEN_1093;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_in3_notify_r <= 1'h0;
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_in3_notify_r <= 1'h0;
                                                            end else begin
                                                              slave_in3_notify_r <= _GEN_1093;
                                                            end
                                                          end else begin
                                                            slave_in3_notify_r <= _GEN_1093;
                                                          end
                                                        end else begin
                                                          slave_in3_notify_r <= _GEN_1093;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            slave_in3_notify_r <= 1'h0;
                                                          end else begin
                                                            slave_in3_notify_r <= _GEN_1093;
                                                          end
                                                        end else begin
                                                          slave_in3_notify_r <= _GEN_1093;
                                                        end
                                                      end else begin
                                                        slave_in3_notify_r <= _GEN_1093;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_in3_notify_r <= 1'h0;
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_in3_notify_r <= 1'h0;
                                                      end else begin
                                                        slave_in3_notify_r <= _GEN_1147;
                                                      end
                                                    end else begin
                                                      slave_in3_notify_r <= _GEN_1147;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (io_master_out_sync) begin
                                                      slave_in3_notify_r <= 1'h0;
                                                    end else begin
                                                      slave_in3_notify_r <= _GEN_1147;
                                                    end
                                                  end else begin
                                                    slave_in3_notify_r <= _GEN_1147;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (io_slave_out1_sync) begin
                                                  slave_in3_notify_r <= 1'h0;
                                                end else begin
                                                  slave_in3_notify_r <= _GEN_1179;
                                                end
                                              end else begin
                                                slave_in3_notify_r <= _GEN_1179;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_in3_notify_r <= 1'h0;
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_in3_notify_r <= 1'h0;
                                                  end else begin
                                                    slave_in3_notify_r <= _GEN_1179;
                                                  end
                                                end else begin
                                                  slave_in3_notify_r <= _GEN_1179;
                                                end
                                              end
                                            end else begin
                                              slave_in3_notify_r <= _GEN_1211;
                                            end
                                          end else begin
                                            slave_in3_notify_r <= _GEN_1211;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              slave_in3_notify_r <= 1'h0;
                                            end else begin
                                              slave_in3_notify_r <= _GEN_1211;
                                            end
                                          end else begin
                                            slave_in3_notify_r <= _GEN_1211;
                                          end
                                        end else begin
                                          slave_in3_notify_r <= _GEN_1211;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_in3_notify_r <= 1'h0;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_in3_notify_r <= 1'h0;
                                              end else begin
                                                slave_in3_notify_r <= _GEN_1211;
                                              end
                                            end else begin
                                              slave_in3_notify_r <= _GEN_1211;
                                            end
                                          end else begin
                                            slave_in3_notify_r <= _GEN_1211;
                                          end
                                        end
                                      end else begin
                                        slave_in3_notify_r <= _GEN_1265;
                                      end
                                    end else begin
                                      slave_in3_notify_r <= _GEN_1265;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_in3_notify_r <= 1'h0;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_in3_notify_r <= 1'h0;
                                        end else begin
                                          slave_in3_notify_r <= _GEN_1265;
                                        end
                                      end else begin
                                        slave_in3_notify_r <= _GEN_1265;
                                      end
                                    end else begin
                                      slave_in3_notify_r <= _GEN_1265;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        slave_in3_notify_r <= 1'h0;
                                      end else begin
                                        slave_in3_notify_r <= _GEN_1265;
                                      end
                                    end else begin
                                      slave_in3_notify_r <= _GEN_1265;
                                    end
                                  end else begin
                                    slave_in3_notify_r <= _GEN_1265;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (io_slave_out2_sync) begin
                                  slave_in3_notify_r <= 1'h0;
                                end else begin
                                  slave_in3_notify_r <= _GEN_1319;
                                end
                              end else begin
                                slave_in3_notify_r <= _GEN_1319;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_in3_notify_r <= 1'h0;
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_in3_notify_r <= 1'h0;
                                  end else begin
                                    slave_in3_notify_r <= _GEN_1319;
                                  end
                                end else begin
                                  slave_in3_notify_r <= _GEN_1319;
                                end
                              end
                            end else begin
                              slave_in3_notify_r <= _GEN_1351;
                            end
                          end else begin
                            slave_in3_notify_r <= _GEN_1351;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              slave_in3_notify_r <= 1'h0;
                            end else begin
                              slave_in3_notify_r <= _GEN_1351;
                            end
                          end else begin
                            slave_in3_notify_r <= _GEN_1351;
                          end
                        end else begin
                          slave_in3_notify_r <= _GEN_1351;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_in3_notify_r <= 1'h0;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_in3_notify_r <= 1'h0;
                              end else begin
                                slave_in3_notify_r <= _GEN_1351;
                              end
                            end else begin
                              slave_in3_notify_r <= _GEN_1351;
                            end
                          end else begin
                            slave_in3_notify_r <= _GEN_1351;
                          end
                        end
                      end else begin
                        slave_in3_notify_r <= _GEN_1405;
                      end
                    end else begin
                      slave_in3_notify_r <= _GEN_1405;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_in3_notify_r <= 1'h1;
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_in3_notify_r <= 1'h0;
                        end else begin
                          slave_in3_notify_r <= _GEN_1405;
                        end
                      end else begin
                        slave_in3_notify_r <= _GEN_1405;
                      end
                    end else begin
                      slave_in3_notify_r <= _GEN_1405;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        slave_in3_notify_r <= 1'h0;
                      end else begin
                        slave_in3_notify_r <= _GEN_1405;
                      end
                    end else begin
                      slave_in3_notify_r <= _GEN_1405;
                    end
                  end else begin
                    slave_in3_notify_r <= _GEN_1405;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (io_slave_out3_sync) begin
                  slave_in3_notify_r <= 1'h1;
                end else begin
                  slave_in3_notify_r <= _GEN_1459;
                end
              end else begin
                slave_in3_notify_r <= _GEN_1459;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                slave_in3_notify_r <= 1'h0;
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_in3_notify_r <= 1'h1;
                  end else begin
                    slave_in3_notify_r <= _GEN_1459;
                  end
                end else begin
                  slave_in3_notify_r <= _GEN_1459;
                end
              end
            end else begin
              slave_in3_notify_r <= _GEN_1491;
            end
          end else begin
            slave_in3_notify_r <= _GEN_1491;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              slave_in3_notify_r <= 1'h0;
            end else begin
              slave_in3_notify_r <= _GEN_1491;
            end
          end else begin
            slave_in3_notify_r <= _GEN_1491;
          end
        end else begin
          slave_in3_notify_r <= _GEN_1491;
        end
      end
    end
    if (reset) begin
      slave_out0_notify_r <= 1'h0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            slave_out0_notify_r <= 1'h0;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  slave_out0_notify_r <= 1'h0;
                end else begin
                  if (_T_518) begin
                    if (io_slave_out3_sync) begin
                      slave_out0_notify_r <= 1'h0;
                    end else begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            slave_out0_notify_r <= 1'h0;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  slave_out0_notify_r <= 1'h0;
                                end else begin
                                  if (_T_479) begin
                                    if (io_slave_out2_sync) begin
                                      slave_out0_notify_r <= 1'h0;
                                    end else begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            slave_out0_notify_r <= 1'h0;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  slave_out0_notify_r <= 1'h0;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (io_slave_out1_sync) begin
                                                      slave_out0_notify_r <= 1'h0;
                                                    end else begin
                                                      if (_T_429) begin
                                                        if (io_master_out_sync) begin
                                                          slave_out0_notify_r <= 1'h0;
                                                        end else begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                slave_out0_notify_r <= 1'h0;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      slave_out0_notify_r <= 1'h0;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (io_slave_out0_sync) begin
                                                                          slave_out0_notify_r <= 1'h0;
                                                                        end else begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    slave_out0_notify_r <= 1'h0;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              slave_out0_notify_r <= 1'h0;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        slave_out0_notify_r <= 1'h0;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  slave_out0_notify_r <= 1'h0;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            slave_out0_notify_r <= 1'h0;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      slave_out0_notify_r <= 1'h0;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    slave_out0_notify_r <= 1'h0;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  slave_out0_notify_r <= 1'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            slave_out0_notify_r <= 1'h1;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      slave_out0_notify_r <= 1'h1;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    slave_out0_notify_r <= 1'h1;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  slave_out0_notify_r <= 1'h1;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                slave_out0_notify_r <= 1'h1;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          slave_out0_notify_r <= 1'h1;
                                                                                                                                                                        end else begin
                                                                                                                                                                          slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        slave_out0_notify_r <= 1'h1;
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_out0_notify_r <= _GEN_91;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      slave_out0_notify_r <= 1'h1;
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_out0_notify_r <= _GEN_91;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_out0_notify_r <= _GEN_91;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_out0_notify_r <= _GEN_91;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out0_notify_r <= _GEN_186;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out0_notify_r <= _GEN_186;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out0_notify_r <= _GEN_186;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                slave_out0_notify_r <= 1'h0;
                                                                                                                                                              end else begin
                                                                                                                                                                slave_out0_notify_r <= _GEN_186;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_out0_notify_r <= _GEN_186;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_out0_notify_r <= _GEN_186;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out0_notify_r <= _GEN_186;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out0_notify_r <= _GEN_186;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out0_notify_r <= _GEN_186;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_out0_notify_r <= _GEN_186;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              slave_out0_notify_r <= 1'h0;
                                                                                                                                                            end else begin
                                                                                                                                                              slave_out0_notify_r <= _GEN_186;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_out0_notify_r <= _GEN_186;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out0_notify_r <= _GEN_186;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out0_notify_r <= _GEN_186;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out0_notify_r <= _GEN_186;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_out0_notify_r <= _GEN_186;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_out0_notify_r <= _GEN_186;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            slave_out0_notify_r <= 1'h0;
                                                                                                                                                          end else begin
                                                                                                                                                            slave_out0_notify_r <= _GEN_186;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out0_notify_r <= _GEN_186;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out0_notify_r <= _GEN_186;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out0_notify_r <= _GEN_186;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_out0_notify_r <= _GEN_186;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_out0_notify_r <= _GEN_186;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_out0_notify_r <= _GEN_186;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out0_notify_r <= _GEN_312;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out0_notify_r <= _GEN_312;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out0_notify_r <= _GEN_312;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  slave_out0_notify_r <= 1'h0;
                                                                                                                                                end else begin
                                                                                                                                                  slave_out0_notify_r <= _GEN_312;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_out0_notify_r <= _GEN_312;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_out0_notify_r <= _GEN_312;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out0_notify_r <= _GEN_312;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out0_notify_r <= _GEN_312;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out0_notify_r <= _GEN_312;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_out0_notify_r <= _GEN_312;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                slave_out0_notify_r <= 1'h0;
                                                                                                                                              end else begin
                                                                                                                                                slave_out0_notify_r <= _GEN_312;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_out0_notify_r <= _GEN_312;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out0_notify_r <= _GEN_312;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out0_notify_r <= _GEN_312;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out0_notify_r <= _GEN_312;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_out0_notify_r <= _GEN_312;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_out0_notify_r <= _GEN_312;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              slave_out0_notify_r <= 1'h0;
                                                                                                                                            end else begin
                                                                                                                                              slave_out0_notify_r <= _GEN_312;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out0_notify_r <= _GEN_312;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out0_notify_r <= _GEN_312;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out0_notify_r <= _GEN_312;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_out0_notify_r <= _GEN_312;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_out0_notify_r <= _GEN_312;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_out0_notify_r <= _GEN_312;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out0_notify_r <= _GEN_438;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    slave_out0_notify_r <= 1'h0;
                                                                                                                                  end else begin
                                                                                                                                    slave_out0_notify_r <= _GEN_438;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_out0_notify_r <= _GEN_438;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_out0_notify_r <= _GEN_438;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out0_notify_r <= _GEN_438;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_out0_notify_r <= _GEN_438;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  slave_out0_notify_r <= 1'h0;
                                                                                                                                end else begin
                                                                                                                                  slave_out0_notify_r <= _GEN_438;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_out0_notify_r <= _GEN_438;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out0_notify_r <= _GEN_438;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_out0_notify_r <= _GEN_438;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_out0_notify_r <= _GEN_438;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                slave_out0_notify_r <= 1'h0;
                                                                                                                              end else begin
                                                                                                                                slave_out0_notify_r <= _GEN_438;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out0_notify_r <= _GEN_438;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_out0_notify_r <= _GEN_438;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_out0_notify_r <= _GEN_438;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_out0_notify_r <= _GEN_438;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out0_notify_r <= _GEN_533;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          slave_out0_notify_r <= 1'h0;
                                                                                                                        end else begin
                                                                                                                          slave_out0_notify_r <= _GEN_533;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_out0_notify_r <= _GEN_533;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_out0_notify_r <= _GEN_533;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out0_notify_r <= _GEN_533;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_out0_notify_r <= _GEN_533;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        slave_out0_notify_r <= 1'h0;
                                                                                                                      end else begin
                                                                                                                        slave_out0_notify_r <= _GEN_533;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_out0_notify_r <= _GEN_533;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out0_notify_r <= _GEN_533;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_out0_notify_r <= _GEN_533;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_out0_notify_r <= _GEN_533;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      slave_out0_notify_r <= 1'h0;
                                                                                                                    end else begin
                                                                                                                      slave_out0_notify_r <= _GEN_533;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out0_notify_r <= _GEN_533;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_out0_notify_r <= _GEN_533;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_out0_notify_r <= _GEN_533;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_out0_notify_r <= _GEN_533;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out0_notify_r <= _GEN_628;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                slave_out0_notify_r <= 1'h0;
                                                                                                              end else begin
                                                                                                                slave_out0_notify_r <= _GEN_628;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_out0_notify_r <= _GEN_628;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_out0_notify_r <= _GEN_628;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out0_notify_r <= _GEN_628;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_out0_notify_r <= _GEN_628;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              slave_out0_notify_r <= 1'h0;
                                                                                                            end else begin
                                                                                                              slave_out0_notify_r <= _GEN_628;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_out0_notify_r <= _GEN_628;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out0_notify_r <= _GEN_628;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_out0_notify_r <= _GEN_628;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_out0_notify_r <= _GEN_628;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            slave_out0_notify_r <= 1'h0;
                                                                                                          end else begin
                                                                                                            slave_out0_notify_r <= _GEN_628;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out0_notify_r <= _GEN_628;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_out0_notify_r <= _GEN_628;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_out0_notify_r <= _GEN_628;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_out0_notify_r <= _GEN_628;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out0_notify_r <= _GEN_723;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      slave_out0_notify_r <= 1'h0;
                                                                                                    end else begin
                                                                                                      slave_out0_notify_r <= _GEN_723;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_out0_notify_r <= _GEN_723;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_out0_notify_r <= _GEN_723;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out0_notify_r <= _GEN_723;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_out0_notify_r <= _GEN_723;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    slave_out0_notify_r <= 1'h0;
                                                                                                  end else begin
                                                                                                    slave_out0_notify_r <= _GEN_723;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_out0_notify_r <= _GEN_723;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out0_notify_r <= _GEN_723;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_out0_notify_r <= _GEN_723;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_out0_notify_r <= _GEN_723;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  slave_out0_notify_r <= 1'h0;
                                                                                                end else begin
                                                                                                  slave_out0_notify_r <= _GEN_723;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out0_notify_r <= _GEN_723;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_out0_notify_r <= _GEN_723;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_out0_notify_r <= _GEN_723;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_out0_notify_r <= _GEN_723;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out0_notify_r <= _GEN_818;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            slave_out0_notify_r <= 1'h0;
                                                                                          end else begin
                                                                                            slave_out0_notify_r <= _GEN_818;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_out0_notify_r <= _GEN_818;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_out0_notify_r <= _GEN_818;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out0_notify_r <= _GEN_818;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_out0_notify_r <= _GEN_818;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          slave_out0_notify_r <= 1'h0;
                                                                                        end else begin
                                                                                          slave_out0_notify_r <= _GEN_818;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_out0_notify_r <= _GEN_818;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out0_notify_r <= _GEN_818;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_out0_notify_r <= _GEN_818;
                                                                                  end
                                                                                end else begin
                                                                                  slave_out0_notify_r <= _GEN_818;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        slave_out0_notify_r <= 1'h0;
                                                                                      end else begin
                                                                                        slave_out0_notify_r <= _GEN_818;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out0_notify_r <= _GEN_818;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_out0_notify_r <= _GEN_818;
                                                                                  end
                                                                                end else begin
                                                                                  slave_out0_notify_r <= _GEN_818;
                                                                                end
                                                                              end else begin
                                                                                slave_out0_notify_r <= _GEN_818;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            slave_out0_notify_r <= _GEN_913;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_out0_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_out0_notify_r <= _GEN_913;
                                                                                end
                                                                              end else begin
                                                                                slave_out0_notify_r <= _GEN_913;
                                                                              end
                                                                            end else begin
                                                                              slave_out0_notify_r <= _GEN_913;
                                                                            end
                                                                          end else begin
                                                                            slave_out0_notify_r <= _GEN_913;
                                                                          end
                                                                        end else begin
                                                                          slave_out0_notify_r <= _GEN_913;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_out0_notify_r <= 1'h0;
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_out0_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_out0_notify_r <= _GEN_913;
                                                                                end
                                                                              end else begin
                                                                                slave_out0_notify_r <= _GEN_913;
                                                                              end
                                                                            end else begin
                                                                              slave_out0_notify_r <= _GEN_913;
                                                                            end
                                                                          end else begin
                                                                            slave_out0_notify_r <= _GEN_913;
                                                                          end
                                                                        end else begin
                                                                          slave_out0_notify_r <= _GEN_913;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                slave_out0_notify_r <= 1'h0;
                                                                              end else begin
                                                                                slave_out0_notify_r <= _GEN_913;
                                                                              end
                                                                            end else begin
                                                                              slave_out0_notify_r <= _GEN_913;
                                                                            end
                                                                          end else begin
                                                                            slave_out0_notify_r <= _GEN_913;
                                                                          end
                                                                        end else begin
                                                                          slave_out0_notify_r <= _GEN_913;
                                                                        end
                                                                      end else begin
                                                                        slave_out0_notify_r <= _GEN_913;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (io_slave_out0_sync) begin
                                                                      slave_out0_notify_r <= 1'h0;
                                                                    end else begin
                                                                      slave_out0_notify_r <= _GEN_1008;
                                                                    end
                                                                  end else begin
                                                                    slave_out0_notify_r <= _GEN_1008;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_out0_notify_r <= 1'h0;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_out0_notify_r <= 1'h0;
                                                                      end else begin
                                                                        slave_out0_notify_r <= _GEN_1008;
                                                                      end
                                                                    end else begin
                                                                      slave_out0_notify_r <= _GEN_1008;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  slave_out0_notify_r <= _GEN_1040;
                                                                end
                                                              end else begin
                                                                slave_out0_notify_r <= _GEN_1040;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  slave_out0_notify_r <= 1'h0;
                                                                end else begin
                                                                  slave_out0_notify_r <= _GEN_1040;
                                                                end
                                                              end else begin
                                                                slave_out0_notify_r <= _GEN_1040;
                                                              end
                                                            end else begin
                                                              slave_out0_notify_r <= _GEN_1040;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_out0_notify_r <= 1'h0;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_out0_notify_r <= 1'h0;
                                                                  end else begin
                                                                    slave_out0_notify_r <= _GEN_1040;
                                                                  end
                                                                end else begin
                                                                  slave_out0_notify_r <= _GEN_1040;
                                                                end
                                                              end else begin
                                                                slave_out0_notify_r <= _GEN_1040;
                                                              end
                                                            end
                                                          end else begin
                                                            slave_out0_notify_r <= _GEN_1094;
                                                          end
                                                        end else begin
                                                          slave_out0_notify_r <= _GEN_1094;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_out0_notify_r <= 1'h0;
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_out0_notify_r <= 1'h0;
                                                            end else begin
                                                              slave_out0_notify_r <= _GEN_1094;
                                                            end
                                                          end else begin
                                                            slave_out0_notify_r <= _GEN_1094;
                                                          end
                                                        end else begin
                                                          slave_out0_notify_r <= _GEN_1094;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            slave_out0_notify_r <= 1'h0;
                                                          end else begin
                                                            slave_out0_notify_r <= _GEN_1094;
                                                          end
                                                        end else begin
                                                          slave_out0_notify_r <= _GEN_1094;
                                                        end
                                                      end else begin
                                                        slave_out0_notify_r <= _GEN_1094;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_out0_notify_r <= 1'h0;
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_out0_notify_r <= 1'h0;
                                                      end else begin
                                                        slave_out0_notify_r <= _GEN_1148;
                                                      end
                                                    end else begin
                                                      slave_out0_notify_r <= _GEN_1148;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (io_master_out_sync) begin
                                                      slave_out0_notify_r <= 1'h0;
                                                    end else begin
                                                      slave_out0_notify_r <= _GEN_1148;
                                                    end
                                                  end else begin
                                                    slave_out0_notify_r <= _GEN_1148;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (io_slave_out1_sync) begin
                                                  slave_out0_notify_r <= 1'h0;
                                                end else begin
                                                  slave_out0_notify_r <= _GEN_1180;
                                                end
                                              end else begin
                                                slave_out0_notify_r <= _GEN_1180;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_out0_notify_r <= 1'h0;
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_out0_notify_r <= 1'h0;
                                                  end else begin
                                                    slave_out0_notify_r <= _GEN_1180;
                                                  end
                                                end else begin
                                                  slave_out0_notify_r <= _GEN_1180;
                                                end
                                              end
                                            end else begin
                                              slave_out0_notify_r <= _GEN_1212;
                                            end
                                          end else begin
                                            slave_out0_notify_r <= _GEN_1212;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              slave_out0_notify_r <= 1'h0;
                                            end else begin
                                              slave_out0_notify_r <= _GEN_1212;
                                            end
                                          end else begin
                                            slave_out0_notify_r <= _GEN_1212;
                                          end
                                        end else begin
                                          slave_out0_notify_r <= _GEN_1212;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_out0_notify_r <= 1'h0;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_out0_notify_r <= 1'h0;
                                              end else begin
                                                slave_out0_notify_r <= _GEN_1212;
                                              end
                                            end else begin
                                              slave_out0_notify_r <= _GEN_1212;
                                            end
                                          end else begin
                                            slave_out0_notify_r <= _GEN_1212;
                                          end
                                        end
                                      end else begin
                                        slave_out0_notify_r <= _GEN_1266;
                                      end
                                    end else begin
                                      slave_out0_notify_r <= _GEN_1266;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_out0_notify_r <= 1'h0;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_out0_notify_r <= 1'h0;
                                        end else begin
                                          slave_out0_notify_r <= _GEN_1266;
                                        end
                                      end else begin
                                        slave_out0_notify_r <= _GEN_1266;
                                      end
                                    end else begin
                                      slave_out0_notify_r <= _GEN_1266;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        slave_out0_notify_r <= 1'h0;
                                      end else begin
                                        slave_out0_notify_r <= _GEN_1266;
                                      end
                                    end else begin
                                      slave_out0_notify_r <= _GEN_1266;
                                    end
                                  end else begin
                                    slave_out0_notify_r <= _GEN_1266;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (io_slave_out2_sync) begin
                                  slave_out0_notify_r <= 1'h0;
                                end else begin
                                  slave_out0_notify_r <= _GEN_1320;
                                end
                              end else begin
                                slave_out0_notify_r <= _GEN_1320;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_out0_notify_r <= 1'h0;
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_out0_notify_r <= 1'h0;
                                  end else begin
                                    slave_out0_notify_r <= _GEN_1320;
                                  end
                                end else begin
                                  slave_out0_notify_r <= _GEN_1320;
                                end
                              end
                            end else begin
                              slave_out0_notify_r <= _GEN_1352;
                            end
                          end else begin
                            slave_out0_notify_r <= _GEN_1352;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              slave_out0_notify_r <= 1'h0;
                            end else begin
                              slave_out0_notify_r <= _GEN_1352;
                            end
                          end else begin
                            slave_out0_notify_r <= _GEN_1352;
                          end
                        end else begin
                          slave_out0_notify_r <= _GEN_1352;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_out0_notify_r <= 1'h0;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_out0_notify_r <= 1'h0;
                              end else begin
                                slave_out0_notify_r <= _GEN_1352;
                              end
                            end else begin
                              slave_out0_notify_r <= _GEN_1352;
                            end
                          end else begin
                            slave_out0_notify_r <= _GEN_1352;
                          end
                        end
                      end else begin
                        slave_out0_notify_r <= _GEN_1406;
                      end
                    end else begin
                      slave_out0_notify_r <= _GEN_1406;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_out0_notify_r <= 1'h0;
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_out0_notify_r <= 1'h0;
                        end else begin
                          slave_out0_notify_r <= _GEN_1406;
                        end
                      end else begin
                        slave_out0_notify_r <= _GEN_1406;
                      end
                    end else begin
                      slave_out0_notify_r <= _GEN_1406;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        slave_out0_notify_r <= 1'h0;
                      end else begin
                        slave_out0_notify_r <= _GEN_1406;
                      end
                    end else begin
                      slave_out0_notify_r <= _GEN_1406;
                    end
                  end else begin
                    slave_out0_notify_r <= _GEN_1406;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (io_slave_out3_sync) begin
                  slave_out0_notify_r <= 1'h0;
                end else begin
                  slave_out0_notify_r <= _GEN_1460;
                end
              end else begin
                slave_out0_notify_r <= _GEN_1460;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                slave_out0_notify_r <= 1'h0;
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_out0_notify_r <= 1'h0;
                  end else begin
                    slave_out0_notify_r <= _GEN_1460;
                  end
                end else begin
                  slave_out0_notify_r <= _GEN_1460;
                end
              end
            end else begin
              slave_out0_notify_r <= _GEN_1492;
            end
          end else begin
            slave_out0_notify_r <= _GEN_1492;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              slave_out0_notify_r <= 1'h0;
            end else begin
              slave_out0_notify_r <= _GEN_1492;
            end
          end else begin
            slave_out0_notify_r <= _GEN_1492;
          end
        end else begin
          slave_out0_notify_r <= _GEN_1492;
        end
      end
    end
    if (reset) begin
      slave_out1_notify_r <= 1'h0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            slave_out1_notify_r <= 1'h0;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  slave_out1_notify_r <= 1'h0;
                end else begin
                  if (_T_518) begin
                    if (io_slave_out3_sync) begin
                      slave_out1_notify_r <= 1'h0;
                    end else begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            slave_out1_notify_r <= 1'h0;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  slave_out1_notify_r <= 1'h0;
                                end else begin
                                  if (_T_479) begin
                                    if (io_slave_out2_sync) begin
                                      slave_out1_notify_r <= 1'h0;
                                    end else begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            slave_out1_notify_r <= 1'h0;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  slave_out1_notify_r <= 1'h0;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (io_slave_out1_sync) begin
                                                      slave_out1_notify_r <= 1'h0;
                                                    end else begin
                                                      if (_T_429) begin
                                                        if (io_master_out_sync) begin
                                                          slave_out1_notify_r <= 1'h0;
                                                        end else begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                slave_out1_notify_r <= 1'h0;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      slave_out1_notify_r <= 1'h0;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (io_slave_out0_sync) begin
                                                                          slave_out1_notify_r <= 1'h0;
                                                                        end else begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    slave_out1_notify_r <= 1'h0;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              slave_out1_notify_r <= 1'h0;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        slave_out1_notify_r <= 1'h0;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  slave_out1_notify_r <= 1'h0;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            slave_out1_notify_r <= 1'h1;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      slave_out1_notify_r <= 1'h1;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    slave_out1_notify_r <= 1'h0;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  slave_out1_notify_r <= 1'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            slave_out1_notify_r <= 1'h0;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      slave_out1_notify_r <= 1'h0;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    slave_out1_notify_r <= 1'h0;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  slave_out1_notify_r <= 1'h0;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                slave_out1_notify_r <= 1'h0;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          slave_out1_notify_r <= 1'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                          slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        slave_out1_notify_r <= 1'h0;
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_out1_notify_r <= _GEN_92;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      slave_out1_notify_r <= 1'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_out1_notify_r <= _GEN_92;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_out1_notify_r <= _GEN_92;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_out1_notify_r <= _GEN_92;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out1_notify_r <= _GEN_187;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out1_notify_r <= _GEN_187;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out1_notify_r <= _GEN_187;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                slave_out1_notify_r <= 1'h0;
                                                                                                                                                              end else begin
                                                                                                                                                                slave_out1_notify_r <= _GEN_187;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_out1_notify_r <= _GEN_187;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_out1_notify_r <= _GEN_187;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out1_notify_r <= _GEN_187;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out1_notify_r <= _GEN_187;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out1_notify_r <= _GEN_187;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_out1_notify_r <= _GEN_187;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              slave_out1_notify_r <= 1'h0;
                                                                                                                                                            end else begin
                                                                                                                                                              slave_out1_notify_r <= _GEN_187;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_out1_notify_r <= _GEN_187;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out1_notify_r <= _GEN_187;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out1_notify_r <= _GEN_187;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out1_notify_r <= _GEN_187;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_out1_notify_r <= _GEN_187;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_out1_notify_r <= _GEN_187;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            slave_out1_notify_r <= 1'h0;
                                                                                                                                                          end else begin
                                                                                                                                                            slave_out1_notify_r <= _GEN_187;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out1_notify_r <= _GEN_187;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out1_notify_r <= _GEN_187;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out1_notify_r <= _GEN_187;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_out1_notify_r <= _GEN_187;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_out1_notify_r <= _GEN_187;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_out1_notify_r <= _GEN_187;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out1_notify_r <= _GEN_313;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out1_notify_r <= _GEN_313;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out1_notify_r <= _GEN_313;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  slave_out1_notify_r <= 1'h0;
                                                                                                                                                end else begin
                                                                                                                                                  slave_out1_notify_r <= _GEN_313;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_out1_notify_r <= _GEN_313;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_out1_notify_r <= _GEN_313;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out1_notify_r <= _GEN_313;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out1_notify_r <= _GEN_313;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out1_notify_r <= _GEN_313;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_out1_notify_r <= _GEN_313;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                slave_out1_notify_r <= 1'h0;
                                                                                                                                              end else begin
                                                                                                                                                slave_out1_notify_r <= _GEN_313;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_out1_notify_r <= _GEN_313;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out1_notify_r <= _GEN_313;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out1_notify_r <= _GEN_313;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out1_notify_r <= _GEN_313;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_out1_notify_r <= _GEN_313;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_out1_notify_r <= _GEN_313;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              slave_out1_notify_r <= 1'h0;
                                                                                                                                            end else begin
                                                                                                                                              slave_out1_notify_r <= _GEN_313;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out1_notify_r <= _GEN_313;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out1_notify_r <= _GEN_313;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out1_notify_r <= _GEN_313;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_out1_notify_r <= _GEN_313;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_out1_notify_r <= _GEN_313;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_out1_notify_r <= _GEN_313;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out1_notify_r <= _GEN_439;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    slave_out1_notify_r <= 1'h1;
                                                                                                                                  end else begin
                                                                                                                                    slave_out1_notify_r <= _GEN_439;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_out1_notify_r <= _GEN_439;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_out1_notify_r <= _GEN_439;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out1_notify_r <= _GEN_439;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_out1_notify_r <= _GEN_439;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  slave_out1_notify_r <= 1'h1;
                                                                                                                                end else begin
                                                                                                                                  slave_out1_notify_r <= _GEN_439;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_out1_notify_r <= _GEN_439;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out1_notify_r <= _GEN_439;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_out1_notify_r <= _GEN_439;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_out1_notify_r <= _GEN_439;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                slave_out1_notify_r <= 1'h1;
                                                                                                                              end else begin
                                                                                                                                slave_out1_notify_r <= _GEN_439;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out1_notify_r <= _GEN_439;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_out1_notify_r <= _GEN_439;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_out1_notify_r <= _GEN_439;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_out1_notify_r <= _GEN_439;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out1_notify_r <= _GEN_534;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          slave_out1_notify_r <= 1'h1;
                                                                                                                        end else begin
                                                                                                                          slave_out1_notify_r <= _GEN_534;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_out1_notify_r <= _GEN_534;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_out1_notify_r <= _GEN_534;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out1_notify_r <= _GEN_534;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_out1_notify_r <= _GEN_534;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        slave_out1_notify_r <= 1'h1;
                                                                                                                      end else begin
                                                                                                                        slave_out1_notify_r <= _GEN_534;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_out1_notify_r <= _GEN_534;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out1_notify_r <= _GEN_534;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_out1_notify_r <= _GEN_534;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_out1_notify_r <= _GEN_534;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      slave_out1_notify_r <= 1'h1;
                                                                                                                    end else begin
                                                                                                                      slave_out1_notify_r <= _GEN_534;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out1_notify_r <= _GEN_534;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_out1_notify_r <= _GEN_534;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_out1_notify_r <= _GEN_534;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_out1_notify_r <= _GEN_534;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out1_notify_r <= _GEN_629;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                slave_out1_notify_r <= 1'h0;
                                                                                                              end else begin
                                                                                                                slave_out1_notify_r <= _GEN_629;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_out1_notify_r <= _GEN_629;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_out1_notify_r <= _GEN_629;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out1_notify_r <= _GEN_629;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_out1_notify_r <= _GEN_629;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              slave_out1_notify_r <= 1'h0;
                                                                                                            end else begin
                                                                                                              slave_out1_notify_r <= _GEN_629;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_out1_notify_r <= _GEN_629;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out1_notify_r <= _GEN_629;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_out1_notify_r <= _GEN_629;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_out1_notify_r <= _GEN_629;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            slave_out1_notify_r <= 1'h0;
                                                                                                          end else begin
                                                                                                            slave_out1_notify_r <= _GEN_629;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out1_notify_r <= _GEN_629;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_out1_notify_r <= _GEN_629;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_out1_notify_r <= _GEN_629;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_out1_notify_r <= _GEN_629;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out1_notify_r <= _GEN_724;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      slave_out1_notify_r <= 1'h0;
                                                                                                    end else begin
                                                                                                      slave_out1_notify_r <= _GEN_724;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_out1_notify_r <= _GEN_724;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_out1_notify_r <= _GEN_724;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out1_notify_r <= _GEN_724;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_out1_notify_r <= _GEN_724;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    slave_out1_notify_r <= 1'h0;
                                                                                                  end else begin
                                                                                                    slave_out1_notify_r <= _GEN_724;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_out1_notify_r <= _GEN_724;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out1_notify_r <= _GEN_724;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_out1_notify_r <= _GEN_724;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_out1_notify_r <= _GEN_724;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  slave_out1_notify_r <= 1'h0;
                                                                                                end else begin
                                                                                                  slave_out1_notify_r <= _GEN_724;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out1_notify_r <= _GEN_724;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_out1_notify_r <= _GEN_724;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_out1_notify_r <= _GEN_724;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_out1_notify_r <= _GEN_724;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out1_notify_r <= _GEN_819;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            slave_out1_notify_r <= 1'h0;
                                                                                          end else begin
                                                                                            slave_out1_notify_r <= _GEN_819;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_out1_notify_r <= _GEN_819;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_out1_notify_r <= _GEN_819;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out1_notify_r <= _GEN_819;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_out1_notify_r <= _GEN_819;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          slave_out1_notify_r <= 1'h0;
                                                                                        end else begin
                                                                                          slave_out1_notify_r <= _GEN_819;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_out1_notify_r <= _GEN_819;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out1_notify_r <= _GEN_819;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_out1_notify_r <= _GEN_819;
                                                                                  end
                                                                                end else begin
                                                                                  slave_out1_notify_r <= _GEN_819;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        slave_out1_notify_r <= 1'h0;
                                                                                      end else begin
                                                                                        slave_out1_notify_r <= _GEN_819;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out1_notify_r <= _GEN_819;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_out1_notify_r <= _GEN_819;
                                                                                  end
                                                                                end else begin
                                                                                  slave_out1_notify_r <= _GEN_819;
                                                                                end
                                                                              end else begin
                                                                                slave_out1_notify_r <= _GEN_819;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            slave_out1_notify_r <= _GEN_914;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_out1_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_out1_notify_r <= _GEN_914;
                                                                                end
                                                                              end else begin
                                                                                slave_out1_notify_r <= _GEN_914;
                                                                              end
                                                                            end else begin
                                                                              slave_out1_notify_r <= _GEN_914;
                                                                            end
                                                                          end else begin
                                                                            slave_out1_notify_r <= _GEN_914;
                                                                          end
                                                                        end else begin
                                                                          slave_out1_notify_r <= _GEN_914;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_out1_notify_r <= 1'h0;
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_out1_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_out1_notify_r <= _GEN_914;
                                                                                end
                                                                              end else begin
                                                                                slave_out1_notify_r <= _GEN_914;
                                                                              end
                                                                            end else begin
                                                                              slave_out1_notify_r <= _GEN_914;
                                                                            end
                                                                          end else begin
                                                                            slave_out1_notify_r <= _GEN_914;
                                                                          end
                                                                        end else begin
                                                                          slave_out1_notify_r <= _GEN_914;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                slave_out1_notify_r <= 1'h0;
                                                                              end else begin
                                                                                slave_out1_notify_r <= _GEN_914;
                                                                              end
                                                                            end else begin
                                                                              slave_out1_notify_r <= _GEN_914;
                                                                            end
                                                                          end else begin
                                                                            slave_out1_notify_r <= _GEN_914;
                                                                          end
                                                                        end else begin
                                                                          slave_out1_notify_r <= _GEN_914;
                                                                        end
                                                                      end else begin
                                                                        slave_out1_notify_r <= _GEN_914;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (io_slave_out0_sync) begin
                                                                      slave_out1_notify_r <= 1'h0;
                                                                    end else begin
                                                                      slave_out1_notify_r <= _GEN_1009;
                                                                    end
                                                                  end else begin
                                                                    slave_out1_notify_r <= _GEN_1009;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_out1_notify_r <= 1'h0;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_out1_notify_r <= 1'h0;
                                                                      end else begin
                                                                        slave_out1_notify_r <= _GEN_1009;
                                                                      end
                                                                    end else begin
                                                                      slave_out1_notify_r <= _GEN_1009;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  slave_out1_notify_r <= _GEN_1041;
                                                                end
                                                              end else begin
                                                                slave_out1_notify_r <= _GEN_1041;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  slave_out1_notify_r <= 1'h0;
                                                                end else begin
                                                                  slave_out1_notify_r <= _GEN_1041;
                                                                end
                                                              end else begin
                                                                slave_out1_notify_r <= _GEN_1041;
                                                              end
                                                            end else begin
                                                              slave_out1_notify_r <= _GEN_1041;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_out1_notify_r <= 1'h0;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_out1_notify_r <= 1'h0;
                                                                  end else begin
                                                                    slave_out1_notify_r <= _GEN_1041;
                                                                  end
                                                                end else begin
                                                                  slave_out1_notify_r <= _GEN_1041;
                                                                end
                                                              end else begin
                                                                slave_out1_notify_r <= _GEN_1041;
                                                              end
                                                            end
                                                          end else begin
                                                            slave_out1_notify_r <= _GEN_1095;
                                                          end
                                                        end else begin
                                                          slave_out1_notify_r <= _GEN_1095;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_out1_notify_r <= 1'h0;
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_out1_notify_r <= 1'h0;
                                                            end else begin
                                                              slave_out1_notify_r <= _GEN_1095;
                                                            end
                                                          end else begin
                                                            slave_out1_notify_r <= _GEN_1095;
                                                          end
                                                        end else begin
                                                          slave_out1_notify_r <= _GEN_1095;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            slave_out1_notify_r <= 1'h0;
                                                          end else begin
                                                            slave_out1_notify_r <= _GEN_1095;
                                                          end
                                                        end else begin
                                                          slave_out1_notify_r <= _GEN_1095;
                                                        end
                                                      end else begin
                                                        slave_out1_notify_r <= _GEN_1095;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_out1_notify_r <= 1'h0;
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_out1_notify_r <= 1'h0;
                                                      end else begin
                                                        slave_out1_notify_r <= _GEN_1149;
                                                      end
                                                    end else begin
                                                      slave_out1_notify_r <= _GEN_1149;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (io_master_out_sync) begin
                                                      slave_out1_notify_r <= 1'h0;
                                                    end else begin
                                                      slave_out1_notify_r <= _GEN_1149;
                                                    end
                                                  end else begin
                                                    slave_out1_notify_r <= _GEN_1149;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (io_slave_out1_sync) begin
                                                  slave_out1_notify_r <= 1'h0;
                                                end else begin
                                                  slave_out1_notify_r <= _GEN_1181;
                                                end
                                              end else begin
                                                slave_out1_notify_r <= _GEN_1181;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_out1_notify_r <= 1'h0;
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_out1_notify_r <= 1'h0;
                                                  end else begin
                                                    slave_out1_notify_r <= _GEN_1181;
                                                  end
                                                end else begin
                                                  slave_out1_notify_r <= _GEN_1181;
                                                end
                                              end
                                            end else begin
                                              slave_out1_notify_r <= _GEN_1213;
                                            end
                                          end else begin
                                            slave_out1_notify_r <= _GEN_1213;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              slave_out1_notify_r <= 1'h0;
                                            end else begin
                                              slave_out1_notify_r <= _GEN_1213;
                                            end
                                          end else begin
                                            slave_out1_notify_r <= _GEN_1213;
                                          end
                                        end else begin
                                          slave_out1_notify_r <= _GEN_1213;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_out1_notify_r <= 1'h0;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_out1_notify_r <= 1'h0;
                                              end else begin
                                                slave_out1_notify_r <= _GEN_1213;
                                              end
                                            end else begin
                                              slave_out1_notify_r <= _GEN_1213;
                                            end
                                          end else begin
                                            slave_out1_notify_r <= _GEN_1213;
                                          end
                                        end
                                      end else begin
                                        slave_out1_notify_r <= _GEN_1267;
                                      end
                                    end else begin
                                      slave_out1_notify_r <= _GEN_1267;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_out1_notify_r <= 1'h0;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_out1_notify_r <= 1'h0;
                                        end else begin
                                          slave_out1_notify_r <= _GEN_1267;
                                        end
                                      end else begin
                                        slave_out1_notify_r <= _GEN_1267;
                                      end
                                    end else begin
                                      slave_out1_notify_r <= _GEN_1267;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        slave_out1_notify_r <= 1'h0;
                                      end else begin
                                        slave_out1_notify_r <= _GEN_1267;
                                      end
                                    end else begin
                                      slave_out1_notify_r <= _GEN_1267;
                                    end
                                  end else begin
                                    slave_out1_notify_r <= _GEN_1267;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (io_slave_out2_sync) begin
                                  slave_out1_notify_r <= 1'h0;
                                end else begin
                                  slave_out1_notify_r <= _GEN_1321;
                                end
                              end else begin
                                slave_out1_notify_r <= _GEN_1321;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_out1_notify_r <= 1'h0;
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_out1_notify_r <= 1'h0;
                                  end else begin
                                    slave_out1_notify_r <= _GEN_1321;
                                  end
                                end else begin
                                  slave_out1_notify_r <= _GEN_1321;
                                end
                              end
                            end else begin
                              slave_out1_notify_r <= _GEN_1353;
                            end
                          end else begin
                            slave_out1_notify_r <= _GEN_1353;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              slave_out1_notify_r <= 1'h0;
                            end else begin
                              slave_out1_notify_r <= _GEN_1353;
                            end
                          end else begin
                            slave_out1_notify_r <= _GEN_1353;
                          end
                        end else begin
                          slave_out1_notify_r <= _GEN_1353;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_out1_notify_r <= 1'h0;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_out1_notify_r <= 1'h0;
                              end else begin
                                slave_out1_notify_r <= _GEN_1353;
                              end
                            end else begin
                              slave_out1_notify_r <= _GEN_1353;
                            end
                          end else begin
                            slave_out1_notify_r <= _GEN_1353;
                          end
                        end
                      end else begin
                        slave_out1_notify_r <= _GEN_1407;
                      end
                    end else begin
                      slave_out1_notify_r <= _GEN_1407;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_out1_notify_r <= 1'h0;
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_out1_notify_r <= 1'h0;
                        end else begin
                          slave_out1_notify_r <= _GEN_1407;
                        end
                      end else begin
                        slave_out1_notify_r <= _GEN_1407;
                      end
                    end else begin
                      slave_out1_notify_r <= _GEN_1407;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        slave_out1_notify_r <= 1'h0;
                      end else begin
                        slave_out1_notify_r <= _GEN_1407;
                      end
                    end else begin
                      slave_out1_notify_r <= _GEN_1407;
                    end
                  end else begin
                    slave_out1_notify_r <= _GEN_1407;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (io_slave_out3_sync) begin
                  slave_out1_notify_r <= 1'h0;
                end else begin
                  slave_out1_notify_r <= _GEN_1461;
                end
              end else begin
                slave_out1_notify_r <= _GEN_1461;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                slave_out1_notify_r <= 1'h0;
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_out1_notify_r <= 1'h0;
                  end else begin
                    slave_out1_notify_r <= _GEN_1461;
                  end
                end else begin
                  slave_out1_notify_r <= _GEN_1461;
                end
              end
            end else begin
              slave_out1_notify_r <= _GEN_1493;
            end
          end else begin
            slave_out1_notify_r <= _GEN_1493;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              slave_out1_notify_r <= 1'h0;
            end else begin
              slave_out1_notify_r <= _GEN_1493;
            end
          end else begin
            slave_out1_notify_r <= _GEN_1493;
          end
        end else begin
          slave_out1_notify_r <= _GEN_1493;
        end
      end
    end
    if (reset) begin
      slave_out2_notify_r <= 1'h0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            slave_out2_notify_r <= 1'h0;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  slave_out2_notify_r <= 1'h0;
                end else begin
                  if (_T_518) begin
                    if (io_slave_out3_sync) begin
                      slave_out2_notify_r <= 1'h0;
                    end else begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            slave_out2_notify_r <= 1'h0;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  slave_out2_notify_r <= 1'h0;
                                end else begin
                                  if (_T_479) begin
                                    if (io_slave_out2_sync) begin
                                      slave_out2_notify_r <= 1'h0;
                                    end else begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            slave_out2_notify_r <= 1'h0;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  slave_out2_notify_r <= 1'h0;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (io_slave_out1_sync) begin
                                                      slave_out2_notify_r <= 1'h0;
                                                    end else begin
                                                      if (_T_429) begin
                                                        if (io_master_out_sync) begin
                                                          slave_out2_notify_r <= 1'h0;
                                                        end else begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                slave_out2_notify_r <= 1'h0;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      slave_out2_notify_r <= 1'h0;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (io_slave_out0_sync) begin
                                                                          slave_out2_notify_r <= 1'h0;
                                                                        end else begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    slave_out2_notify_r <= 1'h0;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              slave_out2_notify_r <= 1'h0;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        slave_out2_notify_r <= 1'h1;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  slave_out2_notify_r <= 1'h1;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            slave_out2_notify_r <= 1'h0;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      slave_out2_notify_r <= 1'h0;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    slave_out2_notify_r <= 1'h0;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  slave_out2_notify_r <= 1'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            slave_out2_notify_r <= 1'h0;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      slave_out2_notify_r <= 1'h0;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    slave_out2_notify_r <= 1'h0;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  slave_out2_notify_r <= 1'h0;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                slave_out2_notify_r <= 1'h0;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          slave_out2_notify_r <= 1'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                          slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        slave_out2_notify_r <= 1'h0;
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_out2_notify_r <= _GEN_93;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      slave_out2_notify_r <= 1'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_out2_notify_r <= _GEN_93;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_out2_notify_r <= _GEN_93;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_out2_notify_r <= _GEN_93;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out2_notify_r <= _GEN_188;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out2_notify_r <= _GEN_188;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out2_notify_r <= _GEN_188;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                slave_out2_notify_r <= 1'h0;
                                                                                                                                                              end else begin
                                                                                                                                                                slave_out2_notify_r <= _GEN_188;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_out2_notify_r <= _GEN_188;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_out2_notify_r <= _GEN_188;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out2_notify_r <= _GEN_188;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out2_notify_r <= _GEN_188;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out2_notify_r <= _GEN_188;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_out2_notify_r <= _GEN_188;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              slave_out2_notify_r <= 1'h0;
                                                                                                                                                            end else begin
                                                                                                                                                              slave_out2_notify_r <= _GEN_188;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_out2_notify_r <= _GEN_188;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out2_notify_r <= _GEN_188;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out2_notify_r <= _GEN_188;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out2_notify_r <= _GEN_188;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_out2_notify_r <= _GEN_188;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_out2_notify_r <= _GEN_188;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            slave_out2_notify_r <= 1'h0;
                                                                                                                                                          end else begin
                                                                                                                                                            slave_out2_notify_r <= _GEN_188;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out2_notify_r <= _GEN_188;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out2_notify_r <= _GEN_188;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out2_notify_r <= _GEN_188;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_out2_notify_r <= _GEN_188;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_out2_notify_r <= _GEN_188;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_out2_notify_r <= _GEN_188;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out2_notify_r <= _GEN_314;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out2_notify_r <= _GEN_314;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out2_notify_r <= _GEN_314;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  slave_out2_notify_r <= 1'h0;
                                                                                                                                                end else begin
                                                                                                                                                  slave_out2_notify_r <= _GEN_314;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_out2_notify_r <= _GEN_314;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_out2_notify_r <= _GEN_314;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out2_notify_r <= _GEN_314;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out2_notify_r <= _GEN_314;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out2_notify_r <= _GEN_314;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_out2_notify_r <= _GEN_314;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                slave_out2_notify_r <= 1'h0;
                                                                                                                                              end else begin
                                                                                                                                                slave_out2_notify_r <= _GEN_314;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_out2_notify_r <= _GEN_314;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out2_notify_r <= _GEN_314;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out2_notify_r <= _GEN_314;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out2_notify_r <= _GEN_314;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_out2_notify_r <= _GEN_314;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_out2_notify_r <= _GEN_314;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              slave_out2_notify_r <= 1'h0;
                                                                                                                                            end else begin
                                                                                                                                              slave_out2_notify_r <= _GEN_314;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out2_notify_r <= _GEN_314;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out2_notify_r <= _GEN_314;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out2_notify_r <= _GEN_314;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_out2_notify_r <= _GEN_314;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_out2_notify_r <= _GEN_314;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_out2_notify_r <= _GEN_314;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out2_notify_r <= _GEN_440;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    slave_out2_notify_r <= 1'h0;
                                                                                                                                  end else begin
                                                                                                                                    slave_out2_notify_r <= _GEN_440;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_out2_notify_r <= _GEN_440;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_out2_notify_r <= _GEN_440;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out2_notify_r <= _GEN_440;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_out2_notify_r <= _GEN_440;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  slave_out2_notify_r <= 1'h0;
                                                                                                                                end else begin
                                                                                                                                  slave_out2_notify_r <= _GEN_440;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_out2_notify_r <= _GEN_440;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out2_notify_r <= _GEN_440;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_out2_notify_r <= _GEN_440;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_out2_notify_r <= _GEN_440;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                slave_out2_notify_r <= 1'h0;
                                                                                                                              end else begin
                                                                                                                                slave_out2_notify_r <= _GEN_440;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out2_notify_r <= _GEN_440;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_out2_notify_r <= _GEN_440;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_out2_notify_r <= _GEN_440;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_out2_notify_r <= _GEN_440;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out2_notify_r <= _GEN_535;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          slave_out2_notify_r <= 1'h0;
                                                                                                                        end else begin
                                                                                                                          slave_out2_notify_r <= _GEN_535;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_out2_notify_r <= _GEN_535;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_out2_notify_r <= _GEN_535;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out2_notify_r <= _GEN_535;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_out2_notify_r <= _GEN_535;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        slave_out2_notify_r <= 1'h0;
                                                                                                                      end else begin
                                                                                                                        slave_out2_notify_r <= _GEN_535;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_out2_notify_r <= _GEN_535;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out2_notify_r <= _GEN_535;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_out2_notify_r <= _GEN_535;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_out2_notify_r <= _GEN_535;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      slave_out2_notify_r <= 1'h0;
                                                                                                                    end else begin
                                                                                                                      slave_out2_notify_r <= _GEN_535;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out2_notify_r <= _GEN_535;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_out2_notify_r <= _GEN_535;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_out2_notify_r <= _GEN_535;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_out2_notify_r <= _GEN_535;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out2_notify_r <= _GEN_630;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                slave_out2_notify_r <= 1'h1;
                                                                                                              end else begin
                                                                                                                slave_out2_notify_r <= _GEN_630;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_out2_notify_r <= _GEN_630;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_out2_notify_r <= _GEN_630;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out2_notify_r <= _GEN_630;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_out2_notify_r <= _GEN_630;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              slave_out2_notify_r <= 1'h1;
                                                                                                            end else begin
                                                                                                              slave_out2_notify_r <= _GEN_630;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_out2_notify_r <= _GEN_630;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out2_notify_r <= _GEN_630;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_out2_notify_r <= _GEN_630;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_out2_notify_r <= _GEN_630;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            slave_out2_notify_r <= 1'h1;
                                                                                                          end else begin
                                                                                                            slave_out2_notify_r <= _GEN_630;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out2_notify_r <= _GEN_630;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_out2_notify_r <= _GEN_630;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_out2_notify_r <= _GEN_630;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_out2_notify_r <= _GEN_630;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out2_notify_r <= _GEN_725;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      slave_out2_notify_r <= 1'h1;
                                                                                                    end else begin
                                                                                                      slave_out2_notify_r <= _GEN_725;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_out2_notify_r <= _GEN_725;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_out2_notify_r <= _GEN_725;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out2_notify_r <= _GEN_725;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_out2_notify_r <= _GEN_725;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    slave_out2_notify_r <= 1'h1;
                                                                                                  end else begin
                                                                                                    slave_out2_notify_r <= _GEN_725;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_out2_notify_r <= _GEN_725;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out2_notify_r <= _GEN_725;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_out2_notify_r <= _GEN_725;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_out2_notify_r <= _GEN_725;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  slave_out2_notify_r <= 1'h1;
                                                                                                end else begin
                                                                                                  slave_out2_notify_r <= _GEN_725;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out2_notify_r <= _GEN_725;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_out2_notify_r <= _GEN_725;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_out2_notify_r <= _GEN_725;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_out2_notify_r <= _GEN_725;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out2_notify_r <= _GEN_820;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            slave_out2_notify_r <= 1'h0;
                                                                                          end else begin
                                                                                            slave_out2_notify_r <= _GEN_820;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_out2_notify_r <= _GEN_820;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_out2_notify_r <= _GEN_820;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out2_notify_r <= _GEN_820;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_out2_notify_r <= _GEN_820;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          slave_out2_notify_r <= 1'h0;
                                                                                        end else begin
                                                                                          slave_out2_notify_r <= _GEN_820;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_out2_notify_r <= _GEN_820;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out2_notify_r <= _GEN_820;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_out2_notify_r <= _GEN_820;
                                                                                  end
                                                                                end else begin
                                                                                  slave_out2_notify_r <= _GEN_820;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        slave_out2_notify_r <= 1'h0;
                                                                                      end else begin
                                                                                        slave_out2_notify_r <= _GEN_820;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out2_notify_r <= _GEN_820;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_out2_notify_r <= _GEN_820;
                                                                                  end
                                                                                end else begin
                                                                                  slave_out2_notify_r <= _GEN_820;
                                                                                end
                                                                              end else begin
                                                                                slave_out2_notify_r <= _GEN_820;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            slave_out2_notify_r <= _GEN_915;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_out2_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_out2_notify_r <= _GEN_915;
                                                                                end
                                                                              end else begin
                                                                                slave_out2_notify_r <= _GEN_915;
                                                                              end
                                                                            end else begin
                                                                              slave_out2_notify_r <= _GEN_915;
                                                                            end
                                                                          end else begin
                                                                            slave_out2_notify_r <= _GEN_915;
                                                                          end
                                                                        end else begin
                                                                          slave_out2_notify_r <= _GEN_915;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_out2_notify_r <= 1'h0;
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_out2_notify_r <= 1'h0;
                                                                                end else begin
                                                                                  slave_out2_notify_r <= _GEN_915;
                                                                                end
                                                                              end else begin
                                                                                slave_out2_notify_r <= _GEN_915;
                                                                              end
                                                                            end else begin
                                                                              slave_out2_notify_r <= _GEN_915;
                                                                            end
                                                                          end else begin
                                                                            slave_out2_notify_r <= _GEN_915;
                                                                          end
                                                                        end else begin
                                                                          slave_out2_notify_r <= _GEN_915;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                slave_out2_notify_r <= 1'h0;
                                                                              end else begin
                                                                                slave_out2_notify_r <= _GEN_915;
                                                                              end
                                                                            end else begin
                                                                              slave_out2_notify_r <= _GEN_915;
                                                                            end
                                                                          end else begin
                                                                            slave_out2_notify_r <= _GEN_915;
                                                                          end
                                                                        end else begin
                                                                          slave_out2_notify_r <= _GEN_915;
                                                                        end
                                                                      end else begin
                                                                        slave_out2_notify_r <= _GEN_915;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (io_slave_out0_sync) begin
                                                                      slave_out2_notify_r <= 1'h0;
                                                                    end else begin
                                                                      slave_out2_notify_r <= _GEN_1010;
                                                                    end
                                                                  end else begin
                                                                    slave_out2_notify_r <= _GEN_1010;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_out2_notify_r <= 1'h0;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_out2_notify_r <= 1'h0;
                                                                      end else begin
                                                                        slave_out2_notify_r <= _GEN_1010;
                                                                      end
                                                                    end else begin
                                                                      slave_out2_notify_r <= _GEN_1010;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  slave_out2_notify_r <= _GEN_1042;
                                                                end
                                                              end else begin
                                                                slave_out2_notify_r <= _GEN_1042;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  slave_out2_notify_r <= 1'h0;
                                                                end else begin
                                                                  slave_out2_notify_r <= _GEN_1042;
                                                                end
                                                              end else begin
                                                                slave_out2_notify_r <= _GEN_1042;
                                                              end
                                                            end else begin
                                                              slave_out2_notify_r <= _GEN_1042;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_out2_notify_r <= 1'h0;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_out2_notify_r <= 1'h0;
                                                                  end else begin
                                                                    slave_out2_notify_r <= _GEN_1042;
                                                                  end
                                                                end else begin
                                                                  slave_out2_notify_r <= _GEN_1042;
                                                                end
                                                              end else begin
                                                                slave_out2_notify_r <= _GEN_1042;
                                                              end
                                                            end
                                                          end else begin
                                                            slave_out2_notify_r <= _GEN_1096;
                                                          end
                                                        end else begin
                                                          slave_out2_notify_r <= _GEN_1096;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_out2_notify_r <= 1'h0;
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_out2_notify_r <= 1'h0;
                                                            end else begin
                                                              slave_out2_notify_r <= _GEN_1096;
                                                            end
                                                          end else begin
                                                            slave_out2_notify_r <= _GEN_1096;
                                                          end
                                                        end else begin
                                                          slave_out2_notify_r <= _GEN_1096;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            slave_out2_notify_r <= 1'h0;
                                                          end else begin
                                                            slave_out2_notify_r <= _GEN_1096;
                                                          end
                                                        end else begin
                                                          slave_out2_notify_r <= _GEN_1096;
                                                        end
                                                      end else begin
                                                        slave_out2_notify_r <= _GEN_1096;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_out2_notify_r <= 1'h0;
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_out2_notify_r <= 1'h0;
                                                      end else begin
                                                        slave_out2_notify_r <= _GEN_1150;
                                                      end
                                                    end else begin
                                                      slave_out2_notify_r <= _GEN_1150;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (io_master_out_sync) begin
                                                      slave_out2_notify_r <= 1'h0;
                                                    end else begin
                                                      slave_out2_notify_r <= _GEN_1150;
                                                    end
                                                  end else begin
                                                    slave_out2_notify_r <= _GEN_1150;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (io_slave_out1_sync) begin
                                                  slave_out2_notify_r <= 1'h0;
                                                end else begin
                                                  slave_out2_notify_r <= _GEN_1182;
                                                end
                                              end else begin
                                                slave_out2_notify_r <= _GEN_1182;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_out2_notify_r <= 1'h0;
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_out2_notify_r <= 1'h0;
                                                  end else begin
                                                    slave_out2_notify_r <= _GEN_1182;
                                                  end
                                                end else begin
                                                  slave_out2_notify_r <= _GEN_1182;
                                                end
                                              end
                                            end else begin
                                              slave_out2_notify_r <= _GEN_1214;
                                            end
                                          end else begin
                                            slave_out2_notify_r <= _GEN_1214;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              slave_out2_notify_r <= 1'h0;
                                            end else begin
                                              slave_out2_notify_r <= _GEN_1214;
                                            end
                                          end else begin
                                            slave_out2_notify_r <= _GEN_1214;
                                          end
                                        end else begin
                                          slave_out2_notify_r <= _GEN_1214;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_out2_notify_r <= 1'h0;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_out2_notify_r <= 1'h0;
                                              end else begin
                                                slave_out2_notify_r <= _GEN_1214;
                                              end
                                            end else begin
                                              slave_out2_notify_r <= _GEN_1214;
                                            end
                                          end else begin
                                            slave_out2_notify_r <= _GEN_1214;
                                          end
                                        end
                                      end else begin
                                        slave_out2_notify_r <= _GEN_1268;
                                      end
                                    end else begin
                                      slave_out2_notify_r <= _GEN_1268;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_out2_notify_r <= 1'h0;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_out2_notify_r <= 1'h0;
                                        end else begin
                                          slave_out2_notify_r <= _GEN_1268;
                                        end
                                      end else begin
                                        slave_out2_notify_r <= _GEN_1268;
                                      end
                                    end else begin
                                      slave_out2_notify_r <= _GEN_1268;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        slave_out2_notify_r <= 1'h0;
                                      end else begin
                                        slave_out2_notify_r <= _GEN_1268;
                                      end
                                    end else begin
                                      slave_out2_notify_r <= _GEN_1268;
                                    end
                                  end else begin
                                    slave_out2_notify_r <= _GEN_1268;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (io_slave_out2_sync) begin
                                  slave_out2_notify_r <= 1'h0;
                                end else begin
                                  slave_out2_notify_r <= _GEN_1322;
                                end
                              end else begin
                                slave_out2_notify_r <= _GEN_1322;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_out2_notify_r <= 1'h0;
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_out2_notify_r <= 1'h0;
                                  end else begin
                                    slave_out2_notify_r <= _GEN_1322;
                                  end
                                end else begin
                                  slave_out2_notify_r <= _GEN_1322;
                                end
                              end
                            end else begin
                              slave_out2_notify_r <= _GEN_1354;
                            end
                          end else begin
                            slave_out2_notify_r <= _GEN_1354;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              slave_out2_notify_r <= 1'h0;
                            end else begin
                              slave_out2_notify_r <= _GEN_1354;
                            end
                          end else begin
                            slave_out2_notify_r <= _GEN_1354;
                          end
                        end else begin
                          slave_out2_notify_r <= _GEN_1354;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_out2_notify_r <= 1'h0;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_out2_notify_r <= 1'h0;
                              end else begin
                                slave_out2_notify_r <= _GEN_1354;
                              end
                            end else begin
                              slave_out2_notify_r <= _GEN_1354;
                            end
                          end else begin
                            slave_out2_notify_r <= _GEN_1354;
                          end
                        end
                      end else begin
                        slave_out2_notify_r <= _GEN_1408;
                      end
                    end else begin
                      slave_out2_notify_r <= _GEN_1408;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_out2_notify_r <= 1'h0;
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_out2_notify_r <= 1'h0;
                        end else begin
                          slave_out2_notify_r <= _GEN_1408;
                        end
                      end else begin
                        slave_out2_notify_r <= _GEN_1408;
                      end
                    end else begin
                      slave_out2_notify_r <= _GEN_1408;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        slave_out2_notify_r <= 1'h0;
                      end else begin
                        slave_out2_notify_r <= _GEN_1408;
                      end
                    end else begin
                      slave_out2_notify_r <= _GEN_1408;
                    end
                  end else begin
                    slave_out2_notify_r <= _GEN_1408;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (io_slave_out3_sync) begin
                  slave_out2_notify_r <= 1'h0;
                end else begin
                  slave_out2_notify_r <= _GEN_1462;
                end
              end else begin
                slave_out2_notify_r <= _GEN_1462;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                slave_out2_notify_r <= 1'h0;
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_out2_notify_r <= 1'h0;
                  end else begin
                    slave_out2_notify_r <= _GEN_1462;
                  end
                end else begin
                  slave_out2_notify_r <= _GEN_1462;
                end
              end
            end else begin
              slave_out2_notify_r <= _GEN_1494;
            end
          end else begin
            slave_out2_notify_r <= _GEN_1494;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              slave_out2_notify_r <= 1'h0;
            end else begin
              slave_out2_notify_r <= _GEN_1494;
            end
          end else begin
            slave_out2_notify_r <= _GEN_1494;
          end
        end else begin
          slave_out2_notify_r <= _GEN_1494;
        end
      end
    end
    if (reset) begin
      slave_out3_notify_r <= 1'h0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            slave_out3_notify_r <= 1'h0;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  slave_out3_notify_r <= 1'h0;
                end else begin
                  if (_T_518) begin
                    if (io_slave_out3_sync) begin
                      slave_out3_notify_r <= 1'h0;
                    end else begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            slave_out3_notify_r <= 1'h0;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  slave_out3_notify_r <= 1'h0;
                                end else begin
                                  if (_T_479) begin
                                    if (io_slave_out2_sync) begin
                                      slave_out3_notify_r <= 1'h0;
                                    end else begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            slave_out3_notify_r <= 1'h0;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  slave_out3_notify_r <= 1'h0;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (io_slave_out1_sync) begin
                                                      slave_out3_notify_r <= 1'h0;
                                                    end else begin
                                                      if (_T_429) begin
                                                        if (io_master_out_sync) begin
                                                          slave_out3_notify_r <= 1'h0;
                                                        end else begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                slave_out3_notify_r <= 1'h0;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      slave_out3_notify_r <= 1'h0;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (io_slave_out0_sync) begin
                                                                          slave_out3_notify_r <= 1'h0;
                                                                        end else begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    slave_out3_notify_r <= 1'h1;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              slave_out3_notify_r <= 1'h1;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        slave_out3_notify_r <= 1'h0;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  slave_out3_notify_r <= 1'h0;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            slave_out3_notify_r <= 1'h0;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      slave_out3_notify_r <= 1'h0;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    slave_out3_notify_r <= 1'h0;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  slave_out3_notify_r <= 1'h0;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            slave_out3_notify_r <= 1'h0;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      slave_out3_notify_r <= 1'h0;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    slave_out3_notify_r <= 1'h0;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  slave_out3_notify_r <= 1'h0;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                slave_out3_notify_r <= 1'h0;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          slave_out3_notify_r <= 1'h0;
                                                                                                                                                                        end else begin
                                                                                                                                                                          slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        slave_out3_notify_r <= 1'h0;
                                                                                                                                                                      end else begin
                                                                                                                                                                        slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_out3_notify_r <= _GEN_94;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      slave_out3_notify_r <= 1'h0;
                                                                                                                                                                    end else begin
                                                                                                                                                                      slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  slave_out3_notify_r <= _GEN_94;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                slave_out3_notify_r <= _GEN_94;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_out3_notify_r <= _GEN_94;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out3_notify_r <= _GEN_189;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out3_notify_r <= _GEN_189;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out3_notify_r <= _GEN_189;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                slave_out3_notify_r <= 1'h0;
                                                                                                                                                              end else begin
                                                                                                                                                                slave_out3_notify_r <= _GEN_189;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              slave_out3_notify_r <= _GEN_189;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_out3_notify_r <= _GEN_189;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out3_notify_r <= _GEN_189;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out3_notify_r <= _GEN_189;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out3_notify_r <= _GEN_189;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_out3_notify_r <= _GEN_189;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              slave_out3_notify_r <= 1'h0;
                                                                                                                                                            end else begin
                                                                                                                                                              slave_out3_notify_r <= _GEN_189;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            slave_out3_notify_r <= _GEN_189;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out3_notify_r <= _GEN_189;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out3_notify_r <= _GEN_189;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out3_notify_r <= _GEN_189;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_out3_notify_r <= _GEN_189;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_out3_notify_r <= _GEN_189;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            slave_out3_notify_r <= 1'h0;
                                                                                                                                                          end else begin
                                                                                                                                                            slave_out3_notify_r <= _GEN_189;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          slave_out3_notify_r <= _GEN_189;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        slave_out3_notify_r <= _GEN_189;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      slave_out3_notify_r <= _GEN_189;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    slave_out3_notify_r <= _GEN_189;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  slave_out3_notify_r <= _GEN_189;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_out3_notify_r <= _GEN_189;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out3_notify_r <= _GEN_315;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out3_notify_r <= _GEN_315;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out3_notify_r <= _GEN_315;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  slave_out3_notify_r <= 1'h0;
                                                                                                                                                end else begin
                                                                                                                                                  slave_out3_notify_r <= _GEN_315;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                slave_out3_notify_r <= _GEN_315;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_out3_notify_r <= _GEN_315;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out3_notify_r <= _GEN_315;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out3_notify_r <= _GEN_315;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out3_notify_r <= _GEN_315;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_out3_notify_r <= _GEN_315;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                slave_out3_notify_r <= 1'h0;
                                                                                                                                              end else begin
                                                                                                                                                slave_out3_notify_r <= _GEN_315;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              slave_out3_notify_r <= _GEN_315;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out3_notify_r <= _GEN_315;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out3_notify_r <= _GEN_315;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out3_notify_r <= _GEN_315;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_out3_notify_r <= _GEN_315;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_out3_notify_r <= _GEN_315;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              slave_out3_notify_r <= 1'h0;
                                                                                                                                            end else begin
                                                                                                                                              slave_out3_notify_r <= _GEN_315;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            slave_out3_notify_r <= _GEN_315;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          slave_out3_notify_r <= _GEN_315;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        slave_out3_notify_r <= _GEN_315;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      slave_out3_notify_r <= _GEN_315;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    slave_out3_notify_r <= _GEN_315;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_out3_notify_r <= _GEN_315;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out3_notify_r <= _GEN_441;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    slave_out3_notify_r <= 1'h0;
                                                                                                                                  end else begin
                                                                                                                                    slave_out3_notify_r <= _GEN_441;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  slave_out3_notify_r <= _GEN_441;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_out3_notify_r <= _GEN_441;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out3_notify_r <= _GEN_441;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_out3_notify_r <= _GEN_441;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  slave_out3_notify_r <= 1'h0;
                                                                                                                                end else begin
                                                                                                                                  slave_out3_notify_r <= _GEN_441;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                slave_out3_notify_r <= _GEN_441;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out3_notify_r <= _GEN_441;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_out3_notify_r <= _GEN_441;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_out3_notify_r <= _GEN_441;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                slave_out3_notify_r <= 1'h0;
                                                                                                                              end else begin
                                                                                                                                slave_out3_notify_r <= _GEN_441;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              slave_out3_notify_r <= _GEN_441;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            slave_out3_notify_r <= _GEN_441;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          slave_out3_notify_r <= _GEN_441;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_out3_notify_r <= _GEN_441;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out3_notify_r <= _GEN_536;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          slave_out3_notify_r <= 1'h0;
                                                                                                                        end else begin
                                                                                                                          slave_out3_notify_r <= _GEN_536;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        slave_out3_notify_r <= _GEN_536;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_out3_notify_r <= _GEN_536;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out3_notify_r <= _GEN_536;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_out3_notify_r <= _GEN_536;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        slave_out3_notify_r <= 1'h0;
                                                                                                                      end else begin
                                                                                                                        slave_out3_notify_r <= _GEN_536;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      slave_out3_notify_r <= _GEN_536;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out3_notify_r <= _GEN_536;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_out3_notify_r <= _GEN_536;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_out3_notify_r <= _GEN_536;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      slave_out3_notify_r <= 1'h0;
                                                                                                                    end else begin
                                                                                                                      slave_out3_notify_r <= _GEN_536;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    slave_out3_notify_r <= _GEN_536;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  slave_out3_notify_r <= _GEN_536;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                slave_out3_notify_r <= _GEN_536;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_out3_notify_r <= _GEN_536;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out3_notify_r <= _GEN_631;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                slave_out3_notify_r <= 1'h0;
                                                                                                              end else begin
                                                                                                                slave_out3_notify_r <= _GEN_631;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              slave_out3_notify_r <= _GEN_631;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_out3_notify_r <= _GEN_631;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out3_notify_r <= _GEN_631;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_out3_notify_r <= _GEN_631;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              slave_out3_notify_r <= 1'h0;
                                                                                                            end else begin
                                                                                                              slave_out3_notify_r <= _GEN_631;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            slave_out3_notify_r <= _GEN_631;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out3_notify_r <= _GEN_631;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_out3_notify_r <= _GEN_631;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_out3_notify_r <= _GEN_631;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            slave_out3_notify_r <= 1'h0;
                                                                                                          end else begin
                                                                                                            slave_out3_notify_r <= _GEN_631;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          slave_out3_notify_r <= _GEN_631;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        slave_out3_notify_r <= _GEN_631;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      slave_out3_notify_r <= _GEN_631;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_out3_notify_r <= _GEN_631;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out3_notify_r <= _GEN_726;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      slave_out3_notify_r <= 1'h0;
                                                                                                    end else begin
                                                                                                      slave_out3_notify_r <= _GEN_726;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    slave_out3_notify_r <= _GEN_726;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_out3_notify_r <= _GEN_726;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out3_notify_r <= _GEN_726;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_out3_notify_r <= _GEN_726;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    slave_out3_notify_r <= 1'h0;
                                                                                                  end else begin
                                                                                                    slave_out3_notify_r <= _GEN_726;
                                                                                                  end
                                                                                                end else begin
                                                                                                  slave_out3_notify_r <= _GEN_726;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out3_notify_r <= _GEN_726;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_out3_notify_r <= _GEN_726;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_out3_notify_r <= _GEN_726;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  slave_out3_notify_r <= 1'h0;
                                                                                                end else begin
                                                                                                  slave_out3_notify_r <= _GEN_726;
                                                                                                end
                                                                                              end else begin
                                                                                                slave_out3_notify_r <= _GEN_726;
                                                                                              end
                                                                                            end else begin
                                                                                              slave_out3_notify_r <= _GEN_726;
                                                                                            end
                                                                                          end else begin
                                                                                            slave_out3_notify_r <= _GEN_726;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_out3_notify_r <= _GEN_726;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out3_notify_r <= _GEN_821;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            slave_out3_notify_r <= 1'h1;
                                                                                          end else begin
                                                                                            slave_out3_notify_r <= _GEN_821;
                                                                                          end
                                                                                        end else begin
                                                                                          slave_out3_notify_r <= _GEN_821;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_out3_notify_r <= _GEN_821;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out3_notify_r <= _GEN_821;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_out3_notify_r <= _GEN_821;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          slave_out3_notify_r <= 1'h1;
                                                                                        end else begin
                                                                                          slave_out3_notify_r <= _GEN_821;
                                                                                        end
                                                                                      end else begin
                                                                                        slave_out3_notify_r <= _GEN_821;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out3_notify_r <= _GEN_821;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_out3_notify_r <= _GEN_821;
                                                                                  end
                                                                                end else begin
                                                                                  slave_out3_notify_r <= _GEN_821;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        slave_out3_notify_r <= 1'h1;
                                                                                      end else begin
                                                                                        slave_out3_notify_r <= _GEN_821;
                                                                                      end
                                                                                    end else begin
                                                                                      slave_out3_notify_r <= _GEN_821;
                                                                                    end
                                                                                  end else begin
                                                                                    slave_out3_notify_r <= _GEN_821;
                                                                                  end
                                                                                end else begin
                                                                                  slave_out3_notify_r <= _GEN_821;
                                                                                end
                                                                              end else begin
                                                                                slave_out3_notify_r <= _GEN_821;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            slave_out3_notify_r <= _GEN_916;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_out3_notify_r <= 1'h1;
                                                                                end else begin
                                                                                  slave_out3_notify_r <= _GEN_916;
                                                                                end
                                                                              end else begin
                                                                                slave_out3_notify_r <= _GEN_916;
                                                                              end
                                                                            end else begin
                                                                              slave_out3_notify_r <= _GEN_916;
                                                                            end
                                                                          end else begin
                                                                            slave_out3_notify_r <= _GEN_916;
                                                                          end
                                                                        end else begin
                                                                          slave_out3_notify_r <= _GEN_916;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_out3_notify_r <= 1'h0;
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  slave_out3_notify_r <= 1'h1;
                                                                                end else begin
                                                                                  slave_out3_notify_r <= _GEN_916;
                                                                                end
                                                                              end else begin
                                                                                slave_out3_notify_r <= _GEN_916;
                                                                              end
                                                                            end else begin
                                                                              slave_out3_notify_r <= _GEN_916;
                                                                            end
                                                                          end else begin
                                                                            slave_out3_notify_r <= _GEN_916;
                                                                          end
                                                                        end else begin
                                                                          slave_out3_notify_r <= _GEN_916;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                slave_out3_notify_r <= 1'h1;
                                                                              end else begin
                                                                                slave_out3_notify_r <= _GEN_916;
                                                                              end
                                                                            end else begin
                                                                              slave_out3_notify_r <= _GEN_916;
                                                                            end
                                                                          end else begin
                                                                            slave_out3_notify_r <= _GEN_916;
                                                                          end
                                                                        end else begin
                                                                          slave_out3_notify_r <= _GEN_916;
                                                                        end
                                                                      end else begin
                                                                        slave_out3_notify_r <= _GEN_916;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (io_slave_out0_sync) begin
                                                                      slave_out3_notify_r <= 1'h0;
                                                                    end else begin
                                                                      slave_out3_notify_r <= _GEN_1011;
                                                                    end
                                                                  end else begin
                                                                    slave_out3_notify_r <= _GEN_1011;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_out3_notify_r <= 1'h0;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        slave_out3_notify_r <= 1'h0;
                                                                      end else begin
                                                                        slave_out3_notify_r <= _GEN_1011;
                                                                      end
                                                                    end else begin
                                                                      slave_out3_notify_r <= _GEN_1011;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  slave_out3_notify_r <= _GEN_1043;
                                                                end
                                                              end else begin
                                                                slave_out3_notify_r <= _GEN_1043;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  slave_out3_notify_r <= 1'h0;
                                                                end else begin
                                                                  slave_out3_notify_r <= _GEN_1043;
                                                                end
                                                              end else begin
                                                                slave_out3_notify_r <= _GEN_1043;
                                                              end
                                                            end else begin
                                                              slave_out3_notify_r <= _GEN_1043;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_out3_notify_r <= 1'h0;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    slave_out3_notify_r <= 1'h0;
                                                                  end else begin
                                                                    slave_out3_notify_r <= _GEN_1043;
                                                                  end
                                                                end else begin
                                                                  slave_out3_notify_r <= _GEN_1043;
                                                                end
                                                              end else begin
                                                                slave_out3_notify_r <= _GEN_1043;
                                                              end
                                                            end
                                                          end else begin
                                                            slave_out3_notify_r <= _GEN_1097;
                                                          end
                                                        end else begin
                                                          slave_out3_notify_r <= _GEN_1097;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_out3_notify_r <= 1'h0;
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              slave_out3_notify_r <= 1'h0;
                                                            end else begin
                                                              slave_out3_notify_r <= _GEN_1097;
                                                            end
                                                          end else begin
                                                            slave_out3_notify_r <= _GEN_1097;
                                                          end
                                                        end else begin
                                                          slave_out3_notify_r <= _GEN_1097;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            slave_out3_notify_r <= 1'h0;
                                                          end else begin
                                                            slave_out3_notify_r <= _GEN_1097;
                                                          end
                                                        end else begin
                                                          slave_out3_notify_r <= _GEN_1097;
                                                        end
                                                      end else begin
                                                        slave_out3_notify_r <= _GEN_1097;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_out3_notify_r <= 1'h0;
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        slave_out3_notify_r <= 1'h0;
                                                      end else begin
                                                        slave_out3_notify_r <= _GEN_1151;
                                                      end
                                                    end else begin
                                                      slave_out3_notify_r <= _GEN_1151;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (io_master_out_sync) begin
                                                      slave_out3_notify_r <= 1'h0;
                                                    end else begin
                                                      slave_out3_notify_r <= _GEN_1151;
                                                    end
                                                  end else begin
                                                    slave_out3_notify_r <= _GEN_1151;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (io_slave_out1_sync) begin
                                                  slave_out3_notify_r <= 1'h0;
                                                end else begin
                                                  slave_out3_notify_r <= _GEN_1183;
                                                end
                                              end else begin
                                                slave_out3_notify_r <= _GEN_1183;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_out3_notify_r <= 1'h0;
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    slave_out3_notify_r <= 1'h0;
                                                  end else begin
                                                    slave_out3_notify_r <= _GEN_1183;
                                                  end
                                                end else begin
                                                  slave_out3_notify_r <= _GEN_1183;
                                                end
                                              end
                                            end else begin
                                              slave_out3_notify_r <= _GEN_1215;
                                            end
                                          end else begin
                                            slave_out3_notify_r <= _GEN_1215;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              slave_out3_notify_r <= 1'h0;
                                            end else begin
                                              slave_out3_notify_r <= _GEN_1215;
                                            end
                                          end else begin
                                            slave_out3_notify_r <= _GEN_1215;
                                          end
                                        end else begin
                                          slave_out3_notify_r <= _GEN_1215;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_out3_notify_r <= 1'h0;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                slave_out3_notify_r <= 1'h0;
                                              end else begin
                                                slave_out3_notify_r <= _GEN_1215;
                                              end
                                            end else begin
                                              slave_out3_notify_r <= _GEN_1215;
                                            end
                                          end else begin
                                            slave_out3_notify_r <= _GEN_1215;
                                          end
                                        end
                                      end else begin
                                        slave_out3_notify_r <= _GEN_1269;
                                      end
                                    end else begin
                                      slave_out3_notify_r <= _GEN_1269;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_out3_notify_r <= 1'h0;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          slave_out3_notify_r <= 1'h0;
                                        end else begin
                                          slave_out3_notify_r <= _GEN_1269;
                                        end
                                      end else begin
                                        slave_out3_notify_r <= _GEN_1269;
                                      end
                                    end else begin
                                      slave_out3_notify_r <= _GEN_1269;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        slave_out3_notify_r <= 1'h0;
                                      end else begin
                                        slave_out3_notify_r <= _GEN_1269;
                                      end
                                    end else begin
                                      slave_out3_notify_r <= _GEN_1269;
                                    end
                                  end else begin
                                    slave_out3_notify_r <= _GEN_1269;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (io_slave_out2_sync) begin
                                  slave_out3_notify_r <= 1'h0;
                                end else begin
                                  slave_out3_notify_r <= _GEN_1323;
                                end
                              end else begin
                                slave_out3_notify_r <= _GEN_1323;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_out3_notify_r <= 1'h0;
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    slave_out3_notify_r <= 1'h0;
                                  end else begin
                                    slave_out3_notify_r <= _GEN_1323;
                                  end
                                end else begin
                                  slave_out3_notify_r <= _GEN_1323;
                                end
                              end
                            end else begin
                              slave_out3_notify_r <= _GEN_1355;
                            end
                          end else begin
                            slave_out3_notify_r <= _GEN_1355;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              slave_out3_notify_r <= 1'h0;
                            end else begin
                              slave_out3_notify_r <= _GEN_1355;
                            end
                          end else begin
                            slave_out3_notify_r <= _GEN_1355;
                          end
                        end else begin
                          slave_out3_notify_r <= _GEN_1355;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_out3_notify_r <= 1'h0;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                slave_out3_notify_r <= 1'h0;
                              end else begin
                                slave_out3_notify_r <= _GEN_1355;
                              end
                            end else begin
                              slave_out3_notify_r <= _GEN_1355;
                            end
                          end else begin
                            slave_out3_notify_r <= _GEN_1355;
                          end
                        end
                      end else begin
                        slave_out3_notify_r <= _GEN_1409;
                      end
                    end else begin
                      slave_out3_notify_r <= _GEN_1409;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_out3_notify_r <= 1'h0;
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          slave_out3_notify_r <= 1'h0;
                        end else begin
                          slave_out3_notify_r <= _GEN_1409;
                        end
                      end else begin
                        slave_out3_notify_r <= _GEN_1409;
                      end
                    end else begin
                      slave_out3_notify_r <= _GEN_1409;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        slave_out3_notify_r <= 1'h0;
                      end else begin
                        slave_out3_notify_r <= _GEN_1409;
                      end
                    end else begin
                      slave_out3_notify_r <= _GEN_1409;
                    end
                  end else begin
                    slave_out3_notify_r <= _GEN_1409;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (io_slave_out3_sync) begin
                  slave_out3_notify_r <= 1'h0;
                end else begin
                  slave_out3_notify_r <= _GEN_1463;
                end
              end else begin
                slave_out3_notify_r <= _GEN_1463;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                slave_out3_notify_r <= 1'h0;
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    slave_out3_notify_r <= 1'h0;
                  end else begin
                    slave_out3_notify_r <= _GEN_1463;
                  end
                end else begin
                  slave_out3_notify_r <= _GEN_1463;
                end
              end
            end else begin
              slave_out3_notify_r <= _GEN_1495;
            end
          end else begin
            slave_out3_notify_r <= _GEN_1495;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              slave_out3_notify_r <= 1'h0;
            end else begin
              slave_out3_notify_r <= _GEN_1495;
            end
          end else begin
            slave_out3_notify_r <= _GEN_1495;
          end
        end else begin
          slave_out3_notify_r <= _GEN_1495;
        end
      end
    end
    if (!(reset)) begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            master_out_r_ack <= io_slave_in3_ack;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  master_out_r_ack <= io_slave_in3_ack;
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        master_out_r_ack <= io_slave_in2_ack;
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              master_out_r_ack <= io_slave_in2_ack;
                            end else begin
                              if (_T_451) begin
                                if (_T_402) begin
                                  if (io_slave_in1_sync) begin
                                    master_out_r_ack <= io_slave_in1_ack;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_404) begin
                                        if (io_slave_in1_sync) begin
                                          master_out_r_ack <= io_slave_in1_ack;
                                        end else begin
                                          if (_T_401) begin
                                            if (_T_402) begin
                                              if (io_slave_in0_sync) begin
                                                master_out_r_ack <= io_slave_in0_ack;
                                              end else begin
                                                if (_T_401) begin
                                                  if (_T_404) begin
                                                    if (io_slave_in0_sync) begin
                                                      master_out_r_ack <= io_slave_in0_ack;
                                                    end else begin
                                                      if (_T_97) begin
                                                        if (_T_143) begin
                                                          if (_T_152) begin
                                                            if (_T_161) begin
                                                              if (_T_170) begin
                                                                if (_T_221) begin
                                                                  if (io_master_in_sync) begin
                                                                    master_out_r_ack <= 32'h0;
                                                                  end else begin
                                                                    if (_T_97) begin
                                                                      if (_T_98) begin
                                                                        if (_T_143) begin
                                                                          if (_T_152) begin
                                                                            if (_T_161) begin
                                                                              if (_T_170) begin
                                                                                if (io_master_in_sync) begin
                                                                                  master_out_r_ack <= 32'h0;
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_97) begin
                                                                    if (_T_98) begin
                                                                      if (_T_143) begin
                                                                        if (_T_152) begin
                                                                          if (_T_161) begin
                                                                            if (_T_170) begin
                                                                              if (io_master_in_sync) begin
                                                                                master_out_r_ack <= 32'h0;
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end else begin
                                                                if (_T_97) begin
                                                                  if (_T_98) begin
                                                                    if (_T_143) begin
                                                                      if (_T_152) begin
                                                                        if (_T_161) begin
                                                                          if (_T_170) begin
                                                                            if (io_master_in_sync) begin
                                                                              master_out_r_ack <= 32'h0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_97) begin
                                                                if (_T_98) begin
                                                                  if (_T_143) begin
                                                                    if (_T_152) begin
                                                                      if (_T_161) begin
                                                                        if (_T_170) begin
                                                                          if (io_master_in_sync) begin
                                                                            master_out_r_ack <= 32'h0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end else begin
                                                            master_out_r_ack <= _GEN_299;
                                                          end
                                                        end else begin
                                                          master_out_r_ack <= _GEN_299;
                                                        end
                                                      end else begin
                                                        master_out_r_ack <= _GEN_299;
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_97) begin
                                                      if (_T_143) begin
                                                        if (_T_152) begin
                                                          if (_T_161) begin
                                                            if (_T_170) begin
                                                              if (_T_221) begin
                                                                if (io_master_in_sync) begin
                                                                  master_out_r_ack <= 32'h0;
                                                                end else begin
                                                                  master_out_r_ack <= _GEN_299;
                                                                end
                                                              end else begin
                                                                master_out_r_ack <= _GEN_299;
                                                              end
                                                            end else begin
                                                              master_out_r_ack <= _GEN_299;
                                                            end
                                                          end else begin
                                                            master_out_r_ack <= _GEN_299;
                                                          end
                                                        end else begin
                                                          master_out_r_ack <= _GEN_299;
                                                        end
                                                      end else begin
                                                        master_out_r_ack <= _GEN_299;
                                                      end
                                                    end else begin
                                                      master_out_r_ack <= _GEN_299;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_97) begin
                                                    if (_T_143) begin
                                                      if (_T_152) begin
                                                        if (_T_161) begin
                                                          if (_T_170) begin
                                                            if (_T_221) begin
                                                              if (io_master_in_sync) begin
                                                                master_out_r_ack <= 32'h0;
                                                              end else begin
                                                                master_out_r_ack <= _GEN_299;
                                                              end
                                                            end else begin
                                                              master_out_r_ack <= _GEN_299;
                                                            end
                                                          end else begin
                                                            master_out_r_ack <= _GEN_299;
                                                          end
                                                        end else begin
                                                          master_out_r_ack <= _GEN_299;
                                                        end
                                                      end else begin
                                                        master_out_r_ack <= _GEN_299;
                                                      end
                                                    end else begin
                                                      master_out_r_ack <= _GEN_299;
                                                    end
                                                  end else begin
                                                    master_out_r_ack <= _GEN_299;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_401) begin
                                                if (_T_404) begin
                                                  if (io_slave_in0_sync) begin
                                                    master_out_r_ack <= io_slave_in0_ack;
                                                  end else begin
                                                    if (_T_97) begin
                                                      if (_T_143) begin
                                                        if (_T_152) begin
                                                          if (_T_161) begin
                                                            if (_T_170) begin
                                                              if (_T_221) begin
                                                                if (io_master_in_sync) begin
                                                                  master_out_r_ack <= 32'h0;
                                                                end else begin
                                                                  master_out_r_ack <= _GEN_299;
                                                                end
                                                              end else begin
                                                                master_out_r_ack <= _GEN_299;
                                                              end
                                                            end else begin
                                                              master_out_r_ack <= _GEN_299;
                                                            end
                                                          end else begin
                                                            master_out_r_ack <= _GEN_299;
                                                          end
                                                        end else begin
                                                          master_out_r_ack <= _GEN_299;
                                                        end
                                                      end else begin
                                                        master_out_r_ack <= _GEN_299;
                                                      end
                                                    end else begin
                                                      master_out_r_ack <= _GEN_299;
                                                    end
                                                  end
                                                end else begin
                                                  master_out_r_ack <= _GEN_425;
                                                end
                                              end else begin
                                                master_out_r_ack <= _GEN_425;
                                              end
                                            end
                                          end else begin
                                            if (_T_401) begin
                                              if (_T_404) begin
                                                if (io_slave_in0_sync) begin
                                                  master_out_r_ack <= io_slave_in0_ack;
                                                end else begin
                                                  master_out_r_ack <= _GEN_425;
                                                end
                                              end else begin
                                                master_out_r_ack <= _GEN_425;
                                              end
                                            end else begin
                                              master_out_r_ack <= _GEN_425;
                                            end
                                          end
                                        end
                                      end else begin
                                        if (_T_401) begin
                                          if (_T_402) begin
                                            if (io_slave_in0_sync) begin
                                              master_out_r_ack <= io_slave_in0_ack;
                                            end else begin
                                              if (_T_401) begin
                                                if (_T_404) begin
                                                  if (io_slave_in0_sync) begin
                                                    master_out_r_ack <= io_slave_in0_ack;
                                                  end else begin
                                                    master_out_r_ack <= _GEN_425;
                                                  end
                                                end else begin
                                                  master_out_r_ack <= _GEN_425;
                                                end
                                              end else begin
                                                master_out_r_ack <= _GEN_425;
                                              end
                                            end
                                          end else begin
                                            master_out_r_ack <= _GEN_1081;
                                          end
                                        end else begin
                                          master_out_r_ack <= _GEN_1081;
                                        end
                                      end
                                    end else begin
                                      if (_T_401) begin
                                        if (_T_402) begin
                                          if (io_slave_in0_sync) begin
                                            master_out_r_ack <= io_slave_in0_ack;
                                          end else begin
                                            master_out_r_ack <= _GEN_1081;
                                          end
                                        end else begin
                                          master_out_r_ack <= _GEN_1081;
                                        end
                                      end else begin
                                        master_out_r_ack <= _GEN_1081;
                                      end
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_404) begin
                                      if (io_slave_in1_sync) begin
                                        master_out_r_ack <= io_slave_in1_ack;
                                      end else begin
                                        if (_T_401) begin
                                          if (_T_402) begin
                                            if (io_slave_in0_sync) begin
                                              master_out_r_ack <= io_slave_in0_ack;
                                            end else begin
                                              master_out_r_ack <= _GEN_1081;
                                            end
                                          end else begin
                                            master_out_r_ack <= _GEN_1081;
                                          end
                                        end else begin
                                          master_out_r_ack <= _GEN_1081;
                                        end
                                      end
                                    end else begin
                                      master_out_r_ack <= _GEN_1135;
                                    end
                                  end else begin
                                    master_out_r_ack <= _GEN_1135;
                                  end
                                end
                              end else begin
                                if (_T_451) begin
                                  if (_T_404) begin
                                    if (io_slave_in1_sync) begin
                                      master_out_r_ack <= io_slave_in1_ack;
                                    end else begin
                                      master_out_r_ack <= _GEN_1135;
                                    end
                                  end else begin
                                    master_out_r_ack <= _GEN_1135;
                                  end
                                end else begin
                                  master_out_r_ack <= _GEN_1135;
                                end
                              end
                            end
                          end else begin
                            if (_T_451) begin
                              if (_T_402) begin
                                if (io_slave_in1_sync) begin
                                  master_out_r_ack <= io_slave_in1_ack;
                                end else begin
                                  if (_T_451) begin
                                    if (_T_404) begin
                                      if (io_slave_in1_sync) begin
                                        master_out_r_ack <= io_slave_in1_ack;
                                      end else begin
                                        master_out_r_ack <= _GEN_1135;
                                      end
                                    end else begin
                                      master_out_r_ack <= _GEN_1135;
                                    end
                                  end else begin
                                    master_out_r_ack <= _GEN_1135;
                                  end
                                end
                              end else begin
                                master_out_r_ack <= _GEN_1253;
                              end
                            end else begin
                              master_out_r_ack <= _GEN_1253;
                            end
                          end
                        end else begin
                          if (_T_451) begin
                            if (_T_402) begin
                              if (io_slave_in1_sync) begin
                                master_out_r_ack <= io_slave_in1_ack;
                              end else begin
                                master_out_r_ack <= _GEN_1253;
                              end
                            end else begin
                              master_out_r_ack <= _GEN_1253;
                            end
                          end else begin
                            master_out_r_ack <= _GEN_1253;
                          end
                        end
                      end
                    end else begin
                      if (_T_490) begin
                        if (_T_404) begin
                          if (io_slave_in2_sync) begin
                            master_out_r_ack <= io_slave_in2_ack;
                          end else begin
                            if (_T_451) begin
                              if (_T_402) begin
                                if (io_slave_in1_sync) begin
                                  master_out_r_ack <= io_slave_in1_ack;
                                end else begin
                                  master_out_r_ack <= _GEN_1253;
                                end
                              end else begin
                                master_out_r_ack <= _GEN_1253;
                              end
                            end else begin
                              master_out_r_ack <= _GEN_1253;
                            end
                          end
                        end else begin
                          master_out_r_ack <= _GEN_1307;
                        end
                      end else begin
                        master_out_r_ack <= _GEN_1307;
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_404) begin
                        if (io_slave_in2_sync) begin
                          master_out_r_ack <= io_slave_in2_ack;
                        end else begin
                          master_out_r_ack <= _GEN_1307;
                        end
                      end else begin
                        master_out_r_ack <= _GEN_1307;
                      end
                    end else begin
                      master_out_r_ack <= _GEN_1307;
                    end
                  end
                end
              end else begin
                if (_T_490) begin
                  if (_T_402) begin
                    if (io_slave_in2_sync) begin
                      master_out_r_ack <= io_slave_in2_ack;
                    end else begin
                      if (_T_490) begin
                        if (_T_404) begin
                          if (io_slave_in2_sync) begin
                            master_out_r_ack <= io_slave_in2_ack;
                          end else begin
                            master_out_r_ack <= _GEN_1307;
                          end
                        end else begin
                          master_out_r_ack <= _GEN_1307;
                        end
                      end else begin
                        master_out_r_ack <= _GEN_1307;
                      end
                    end
                  end else begin
                    master_out_r_ack <= _GEN_1393;
                  end
                end else begin
                  master_out_r_ack <= _GEN_1393;
                end
              end
            end else begin
              if (_T_490) begin
                if (_T_402) begin
                  if (io_slave_in2_sync) begin
                    master_out_r_ack <= io_slave_in2_ack;
                  end else begin
                    master_out_r_ack <= _GEN_1393;
                  end
                end else begin
                  master_out_r_ack <= _GEN_1393;
                end
              end else begin
                master_out_r_ack <= _GEN_1393;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                master_out_r_ack <= io_slave_in3_ack;
              end else begin
                if (_T_490) begin
                  if (_T_402) begin
                    if (io_slave_in2_sync) begin
                      master_out_r_ack <= io_slave_in2_ack;
                    end else begin
                      master_out_r_ack <= _GEN_1393;
                    end
                  end else begin
                    master_out_r_ack <= _GEN_1393;
                  end
                end else begin
                  master_out_r_ack <= _GEN_1393;
                end
              end
            end else begin
              master_out_r_ack <= _GEN_1447;
            end
          end else begin
            master_out_r_ack <= _GEN_1447;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              master_out_r_ack <= io_slave_in3_ack;
            end else begin
              master_out_r_ack <= _GEN_1447;
            end
          end else begin
            master_out_r_ack <= _GEN_1447;
          end
        end else begin
          master_out_r_ack <= _GEN_1447;
        end
      end
    end
    if (!(reset)) begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            master_out_r_data <= 32'sh0;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  master_out_r_data <= io_slave_in3_data;
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        master_out_r_data <= 32'sh0;
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              master_out_r_data <= io_slave_in2_data;
                            end else begin
                              if (_T_451) begin
                                if (_T_402) begin
                                  if (io_slave_in1_sync) begin
                                    master_out_r_data <= 32'sh0;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_404) begin
                                        if (io_slave_in1_sync) begin
                                          master_out_r_data <= io_slave_in1_data;
                                        end else begin
                                          if (_T_401) begin
                                            if (_T_402) begin
                                              if (io_slave_in0_sync) begin
                                                master_out_r_data <= 32'sh0;
                                              end else begin
                                                if (_T_401) begin
                                                  if (_T_404) begin
                                                    if (io_slave_in0_sync) begin
                                                      master_out_r_data <= io_slave_in0_data;
                                                    end else begin
                                                      if (_T_97) begin
                                                        if (_T_143) begin
                                                          if (_T_152) begin
                                                            if (_T_161) begin
                                                              if (_T_170) begin
                                                                if (_T_221) begin
                                                                  if (io_master_in_sync) begin
                                                                    master_out_r_data <= 32'sh0;
                                                                  end else begin
                                                                    if (_T_97) begin
                                                                      if (_T_98) begin
                                                                        if (_T_143) begin
                                                                          if (_T_152) begin
                                                                            if (_T_161) begin
                                                                              if (_T_170) begin
                                                                                if (io_master_in_sync) begin
                                                                                  master_out_r_data <= 32'sh0;
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_97) begin
                                                                    if (_T_98) begin
                                                                      if (_T_143) begin
                                                                        if (_T_152) begin
                                                                          if (_T_161) begin
                                                                            if (_T_170) begin
                                                                              if (io_master_in_sync) begin
                                                                                master_out_r_data <= 32'sh0;
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end else begin
                                                                if (_T_97) begin
                                                                  if (_T_98) begin
                                                                    if (_T_143) begin
                                                                      if (_T_152) begin
                                                                        if (_T_161) begin
                                                                          if (_T_170) begin
                                                                            if (io_master_in_sync) begin
                                                                              master_out_r_data <= 32'sh0;
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_97) begin
                                                                if (_T_98) begin
                                                                  if (_T_143) begin
                                                                    if (_T_152) begin
                                                                      if (_T_161) begin
                                                                        if (_T_170) begin
                                                                          if (io_master_in_sync) begin
                                                                            master_out_r_data <= 32'sh0;
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end else begin
                                                            master_out_r_data <= _GEN_300;
                                                          end
                                                        end else begin
                                                          master_out_r_data <= _GEN_300;
                                                        end
                                                      end else begin
                                                        master_out_r_data <= _GEN_300;
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_97) begin
                                                      if (_T_143) begin
                                                        if (_T_152) begin
                                                          if (_T_161) begin
                                                            if (_T_170) begin
                                                              if (_T_221) begin
                                                                if (io_master_in_sync) begin
                                                                  master_out_r_data <= 32'sh0;
                                                                end else begin
                                                                  master_out_r_data <= _GEN_300;
                                                                end
                                                              end else begin
                                                                master_out_r_data <= _GEN_300;
                                                              end
                                                            end else begin
                                                              master_out_r_data <= _GEN_300;
                                                            end
                                                          end else begin
                                                            master_out_r_data <= _GEN_300;
                                                          end
                                                        end else begin
                                                          master_out_r_data <= _GEN_300;
                                                        end
                                                      end else begin
                                                        master_out_r_data <= _GEN_300;
                                                      end
                                                    end else begin
                                                      master_out_r_data <= _GEN_300;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_97) begin
                                                    if (_T_143) begin
                                                      if (_T_152) begin
                                                        if (_T_161) begin
                                                          if (_T_170) begin
                                                            if (_T_221) begin
                                                              if (io_master_in_sync) begin
                                                                master_out_r_data <= 32'sh0;
                                                              end else begin
                                                                master_out_r_data <= _GEN_300;
                                                              end
                                                            end else begin
                                                              master_out_r_data <= _GEN_300;
                                                            end
                                                          end else begin
                                                            master_out_r_data <= _GEN_300;
                                                          end
                                                        end else begin
                                                          master_out_r_data <= _GEN_300;
                                                        end
                                                      end else begin
                                                        master_out_r_data <= _GEN_300;
                                                      end
                                                    end else begin
                                                      master_out_r_data <= _GEN_300;
                                                    end
                                                  end else begin
                                                    master_out_r_data <= _GEN_300;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_401) begin
                                                if (_T_404) begin
                                                  if (io_slave_in0_sync) begin
                                                    master_out_r_data <= io_slave_in0_data;
                                                  end else begin
                                                    if (_T_97) begin
                                                      if (_T_143) begin
                                                        if (_T_152) begin
                                                          if (_T_161) begin
                                                            if (_T_170) begin
                                                              if (_T_221) begin
                                                                if (io_master_in_sync) begin
                                                                  master_out_r_data <= 32'sh0;
                                                                end else begin
                                                                  master_out_r_data <= _GEN_300;
                                                                end
                                                              end else begin
                                                                master_out_r_data <= _GEN_300;
                                                              end
                                                            end else begin
                                                              master_out_r_data <= _GEN_300;
                                                            end
                                                          end else begin
                                                            master_out_r_data <= _GEN_300;
                                                          end
                                                        end else begin
                                                          master_out_r_data <= _GEN_300;
                                                        end
                                                      end else begin
                                                        master_out_r_data <= _GEN_300;
                                                      end
                                                    end else begin
                                                      master_out_r_data <= _GEN_300;
                                                    end
                                                  end
                                                end else begin
                                                  master_out_r_data <= _GEN_426;
                                                end
                                              end else begin
                                                master_out_r_data <= _GEN_426;
                                              end
                                            end
                                          end else begin
                                            if (_T_401) begin
                                              if (_T_404) begin
                                                if (io_slave_in0_sync) begin
                                                  master_out_r_data <= io_slave_in0_data;
                                                end else begin
                                                  master_out_r_data <= _GEN_426;
                                                end
                                              end else begin
                                                master_out_r_data <= _GEN_426;
                                              end
                                            end else begin
                                              master_out_r_data <= _GEN_426;
                                            end
                                          end
                                        end
                                      end else begin
                                        if (_T_401) begin
                                          if (_T_402) begin
                                            if (io_slave_in0_sync) begin
                                              master_out_r_data <= 32'sh0;
                                            end else begin
                                              if (_T_401) begin
                                                if (_T_404) begin
                                                  if (io_slave_in0_sync) begin
                                                    master_out_r_data <= io_slave_in0_data;
                                                  end else begin
                                                    master_out_r_data <= _GEN_426;
                                                  end
                                                end else begin
                                                  master_out_r_data <= _GEN_426;
                                                end
                                              end else begin
                                                master_out_r_data <= _GEN_426;
                                              end
                                            end
                                          end else begin
                                            master_out_r_data <= _GEN_1082;
                                          end
                                        end else begin
                                          master_out_r_data <= _GEN_1082;
                                        end
                                      end
                                    end else begin
                                      if (_T_401) begin
                                        if (_T_402) begin
                                          if (io_slave_in0_sync) begin
                                            master_out_r_data <= 32'sh0;
                                          end else begin
                                            master_out_r_data <= _GEN_1082;
                                          end
                                        end else begin
                                          master_out_r_data <= _GEN_1082;
                                        end
                                      end else begin
                                        master_out_r_data <= _GEN_1082;
                                      end
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_404) begin
                                      if (io_slave_in1_sync) begin
                                        master_out_r_data <= io_slave_in1_data;
                                      end else begin
                                        if (_T_401) begin
                                          if (_T_402) begin
                                            if (io_slave_in0_sync) begin
                                              master_out_r_data <= 32'sh0;
                                            end else begin
                                              master_out_r_data <= _GEN_1082;
                                            end
                                          end else begin
                                            master_out_r_data <= _GEN_1082;
                                          end
                                        end else begin
                                          master_out_r_data <= _GEN_1082;
                                        end
                                      end
                                    end else begin
                                      master_out_r_data <= _GEN_1136;
                                    end
                                  end else begin
                                    master_out_r_data <= _GEN_1136;
                                  end
                                end
                              end else begin
                                if (_T_451) begin
                                  if (_T_404) begin
                                    if (io_slave_in1_sync) begin
                                      master_out_r_data <= io_slave_in1_data;
                                    end else begin
                                      master_out_r_data <= _GEN_1136;
                                    end
                                  end else begin
                                    master_out_r_data <= _GEN_1136;
                                  end
                                end else begin
                                  master_out_r_data <= _GEN_1136;
                                end
                              end
                            end
                          end else begin
                            if (_T_451) begin
                              if (_T_402) begin
                                if (io_slave_in1_sync) begin
                                  master_out_r_data <= 32'sh0;
                                end else begin
                                  if (_T_451) begin
                                    if (_T_404) begin
                                      if (io_slave_in1_sync) begin
                                        master_out_r_data <= io_slave_in1_data;
                                      end else begin
                                        master_out_r_data <= _GEN_1136;
                                      end
                                    end else begin
                                      master_out_r_data <= _GEN_1136;
                                    end
                                  end else begin
                                    master_out_r_data <= _GEN_1136;
                                  end
                                end
                              end else begin
                                master_out_r_data <= _GEN_1254;
                              end
                            end else begin
                              master_out_r_data <= _GEN_1254;
                            end
                          end
                        end else begin
                          if (_T_451) begin
                            if (_T_402) begin
                              if (io_slave_in1_sync) begin
                                master_out_r_data <= 32'sh0;
                              end else begin
                                master_out_r_data <= _GEN_1254;
                              end
                            end else begin
                              master_out_r_data <= _GEN_1254;
                            end
                          end else begin
                            master_out_r_data <= _GEN_1254;
                          end
                        end
                      end
                    end else begin
                      if (_T_490) begin
                        if (_T_404) begin
                          if (io_slave_in2_sync) begin
                            master_out_r_data <= io_slave_in2_data;
                          end else begin
                            if (_T_451) begin
                              if (_T_402) begin
                                if (io_slave_in1_sync) begin
                                  master_out_r_data <= 32'sh0;
                                end else begin
                                  master_out_r_data <= _GEN_1254;
                                end
                              end else begin
                                master_out_r_data <= _GEN_1254;
                              end
                            end else begin
                              master_out_r_data <= _GEN_1254;
                            end
                          end
                        end else begin
                          master_out_r_data <= _GEN_1308;
                        end
                      end else begin
                        master_out_r_data <= _GEN_1308;
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_404) begin
                        if (io_slave_in2_sync) begin
                          master_out_r_data <= io_slave_in2_data;
                        end else begin
                          master_out_r_data <= _GEN_1308;
                        end
                      end else begin
                        master_out_r_data <= _GEN_1308;
                      end
                    end else begin
                      master_out_r_data <= _GEN_1308;
                    end
                  end
                end
              end else begin
                if (_T_490) begin
                  if (_T_402) begin
                    if (io_slave_in2_sync) begin
                      master_out_r_data <= 32'sh0;
                    end else begin
                      if (_T_490) begin
                        if (_T_404) begin
                          if (io_slave_in2_sync) begin
                            master_out_r_data <= io_slave_in2_data;
                          end else begin
                            master_out_r_data <= _GEN_1308;
                          end
                        end else begin
                          master_out_r_data <= _GEN_1308;
                        end
                      end else begin
                        master_out_r_data <= _GEN_1308;
                      end
                    end
                  end else begin
                    master_out_r_data <= _GEN_1394;
                  end
                end else begin
                  master_out_r_data <= _GEN_1394;
                end
              end
            end else begin
              if (_T_490) begin
                if (_T_402) begin
                  if (io_slave_in2_sync) begin
                    master_out_r_data <= 32'sh0;
                  end else begin
                    master_out_r_data <= _GEN_1394;
                  end
                end else begin
                  master_out_r_data <= _GEN_1394;
                end
              end else begin
                master_out_r_data <= _GEN_1394;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                master_out_r_data <= io_slave_in3_data;
              end else begin
                if (_T_490) begin
                  if (_T_402) begin
                    if (io_slave_in2_sync) begin
                      master_out_r_data <= 32'sh0;
                    end else begin
                      master_out_r_data <= _GEN_1394;
                    end
                  end else begin
                    master_out_r_data <= _GEN_1394;
                  end
                end else begin
                  master_out_r_data <= _GEN_1394;
                end
              end
            end else begin
              master_out_r_data <= _GEN_1448;
            end
          end else begin
            master_out_r_data <= _GEN_1448;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              master_out_r_data <= io_slave_in3_data;
            end else begin
              master_out_r_data <= _GEN_1448;
            end
          end else begin
            master_out_r_data <= _GEN_1448;
          end
        end else begin
          master_out_r_data <= _GEN_1448;
        end
      end
    end
    if (!(reset)) begin
      if (_T_97) begin
        if (_T_98) begin
          if (_T_102) begin
            if (_T_104) begin
              if (io_master_in_sync) begin
                slave_out0_r_addr <= io_master_in_addr;
              end else begin
                if (_T_97) begin
                  if (_T_100) begin
                    if (_T_102) begin
                      if (_T_104) begin
                        if (io_master_in_sync) begin
                          slave_out0_r_addr <= io_master_in_addr;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_97) begin
                if (_T_100) begin
                  if (_T_102) begin
                    if (_T_104) begin
                      if (io_master_in_sync) begin
                        slave_out0_r_addr <= io_master_in_addr;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_97) begin
              if (_T_100) begin
                if (_T_102) begin
                  if (_T_104) begin
                    if (io_master_in_sync) begin
                      slave_out0_r_addr <= io_master_in_addr;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_97) begin
            if (_T_100) begin
              if (_T_102) begin
                if (_T_104) begin
                  if (io_master_in_sync) begin
                    slave_out0_r_addr <= io_master_in_addr;
                  end
                end
              end
            end
          end
        end
      end else begin
        slave_out0_r_addr <= _GEN_82;
      end
    end
    if (!(reset)) begin
      if (_T_97) begin
        if (_T_98) begin
          if (_T_102) begin
            if (_T_104) begin
              if (io_master_in_sync) begin
                slave_out0_r_data <= 32'sh0;
              end else begin
                if (_T_97) begin
                  if (_T_100) begin
                    if (_T_102) begin
                      if (_T_104) begin
                        if (io_master_in_sync) begin
                          slave_out0_r_data <= io_master_in_data;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_97) begin
                if (_T_100) begin
                  if (_T_102) begin
                    if (_T_104) begin
                      if (io_master_in_sync) begin
                        slave_out0_r_data <= io_master_in_data;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_97) begin
              if (_T_100) begin
                if (_T_102) begin
                  if (_T_104) begin
                    if (io_master_in_sync) begin
                      slave_out0_r_data <= io_master_in_data;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_97) begin
            if (_T_100) begin
              if (_T_102) begin
                if (_T_104) begin
                  if (io_master_in_sync) begin
                    slave_out0_r_data <= io_master_in_data;
                  end
                end
              end
            end
          end
        end
      end else begin
        slave_out0_r_data <= _GEN_83;
      end
    end
    if (!(reset)) begin
      if (_T_97) begin
        if (_T_98) begin
          if (_T_102) begin
            if (_T_104) begin
              if (io_master_in_sync) begin
                slave_out0_r_trans_type <= io_master_in_trans_type;
              end else begin
                if (_T_97) begin
                  if (_T_100) begin
                    if (_T_102) begin
                      if (_T_104) begin
                        if (io_master_in_sync) begin
                          slave_out0_r_trans_type <= io_master_in_trans_type;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_97) begin
                if (_T_100) begin
                  if (_T_102) begin
                    if (_T_104) begin
                      if (io_master_in_sync) begin
                        slave_out0_r_trans_type <= io_master_in_trans_type;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_97) begin
              if (_T_100) begin
                if (_T_102) begin
                  if (_T_104) begin
                    if (io_master_in_sync) begin
                      slave_out0_r_trans_type <= io_master_in_trans_type;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_97) begin
            if (_T_100) begin
              if (_T_102) begin
                if (_T_104) begin
                  if (io_master_in_sync) begin
                    slave_out0_r_trans_type <= io_master_in_trans_type;
                  end
                end
              end
            end
          end
        end
      end else begin
        slave_out0_r_trans_type <= _GEN_84;
      end
    end
    if (!(reset)) begin
      if (_T_97) begin
        if (_T_98) begin
          if (_T_145) begin
            if (_T_241) begin
              if (io_master_in_sync) begin
                slave_out1_r_addr <= _T_245;
              end else begin
                if (_T_97) begin
                  if (_T_100) begin
                    if (_T_145) begin
                      if (_T_241) begin
                        if (io_master_in_sync) begin
                          slave_out1_r_addr <= _T_245;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_97) begin
                if (_T_100) begin
                  if (_T_145) begin
                    if (_T_241) begin
                      if (io_master_in_sync) begin
                        slave_out1_r_addr <= _T_245;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_97) begin
              if (_T_100) begin
                if (_T_145) begin
                  if (_T_241) begin
                    if (io_master_in_sync) begin
                      slave_out1_r_addr <= _T_245;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_97) begin
            if (_T_100) begin
              if (_T_145) begin
                if (_T_241) begin
                  if (io_master_in_sync) begin
                    slave_out1_r_addr <= _T_245;
                  end
                end
              end
            end
          end
        end
      end else begin
        slave_out1_r_addr <= _GEN_524;
      end
    end
    if (!(reset)) begin
      if (_T_97) begin
        if (_T_98) begin
          if (_T_145) begin
            if (_T_241) begin
              if (io_master_in_sync) begin
                slave_out1_r_data <= 32'sh0;
              end else begin
                if (_T_97) begin
                  if (_T_100) begin
                    if (_T_145) begin
                      if (_T_241) begin
                        if (io_master_in_sync) begin
                          slave_out1_r_data <= io_master_in_data;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_97) begin
                if (_T_100) begin
                  if (_T_145) begin
                    if (_T_241) begin
                      if (io_master_in_sync) begin
                        slave_out1_r_data <= io_master_in_data;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_97) begin
              if (_T_100) begin
                if (_T_145) begin
                  if (_T_241) begin
                    if (io_master_in_sync) begin
                      slave_out1_r_data <= io_master_in_data;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_97) begin
            if (_T_100) begin
              if (_T_145) begin
                if (_T_241) begin
                  if (io_master_in_sync) begin
                    slave_out1_r_data <= io_master_in_data;
                  end
                end
              end
            end
          end
        end
      end else begin
        slave_out1_r_data <= _GEN_525;
      end
    end
    if (!(reset)) begin
      if (_T_97) begin
        if (_T_98) begin
          if (_T_145) begin
            if (_T_241) begin
              if (io_master_in_sync) begin
                slave_out1_r_trans_type <= io_master_in_trans_type;
              end else begin
                if (_T_97) begin
                  if (_T_100) begin
                    if (_T_145) begin
                      if (_T_241) begin
                        if (io_master_in_sync) begin
                          slave_out1_r_trans_type <= io_master_in_trans_type;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_97) begin
                if (_T_100) begin
                  if (_T_145) begin
                    if (_T_241) begin
                      if (io_master_in_sync) begin
                        slave_out1_r_trans_type <= io_master_in_trans_type;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_97) begin
              if (_T_100) begin
                if (_T_145) begin
                  if (_T_241) begin
                    if (io_master_in_sync) begin
                      slave_out1_r_trans_type <= io_master_in_trans_type;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_97) begin
            if (_T_100) begin
              if (_T_145) begin
                if (_T_241) begin
                  if (io_master_in_sync) begin
                    slave_out1_r_trans_type <= io_master_in_trans_type;
                  end
                end
              end
            end
          end
        end
      end else begin
        slave_out1_r_trans_type <= _GEN_526;
      end
    end
    if (!(reset)) begin
      if (_T_97) begin
        if (_T_98) begin
          if (_T_154) begin
            if (_T_293) begin
              if (io_master_in_sync) begin
                slave_out2_r_addr <= _T_297;
              end else begin
                if (_T_97) begin
                  if (_T_100) begin
                    if (_T_154) begin
                      if (_T_293) begin
                        if (io_master_in_sync) begin
                          slave_out2_r_addr <= _T_297;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_97) begin
                if (_T_100) begin
                  if (_T_154) begin
                    if (_T_293) begin
                      if (io_master_in_sync) begin
                        slave_out2_r_addr <= _T_297;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_97) begin
              if (_T_100) begin
                if (_T_154) begin
                  if (_T_293) begin
                    if (io_master_in_sync) begin
                      slave_out2_r_addr <= _T_297;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_97) begin
            if (_T_100) begin
              if (_T_154) begin
                if (_T_293) begin
                  if (io_master_in_sync) begin
                    slave_out2_r_addr <= _T_297;
                  end
                end
              end
            end
          end
        end
      end else begin
        slave_out2_r_addr <= _GEN_714;
      end
    end
    if (!(reset)) begin
      if (_T_97) begin
        if (_T_98) begin
          if (_T_154) begin
            if (_T_293) begin
              if (io_master_in_sync) begin
                slave_out2_r_data <= 32'sh0;
              end else begin
                if (_T_97) begin
                  if (_T_100) begin
                    if (_T_154) begin
                      if (_T_293) begin
                        if (io_master_in_sync) begin
                          slave_out2_r_data <= io_master_in_data;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_97) begin
                if (_T_100) begin
                  if (_T_154) begin
                    if (_T_293) begin
                      if (io_master_in_sync) begin
                        slave_out2_r_data <= io_master_in_data;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_97) begin
              if (_T_100) begin
                if (_T_154) begin
                  if (_T_293) begin
                    if (io_master_in_sync) begin
                      slave_out2_r_data <= io_master_in_data;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_97) begin
            if (_T_100) begin
              if (_T_154) begin
                if (_T_293) begin
                  if (io_master_in_sync) begin
                    slave_out2_r_data <= io_master_in_data;
                  end
                end
              end
            end
          end
        end
      end else begin
        slave_out2_r_data <= _GEN_715;
      end
    end
    if (!(reset)) begin
      if (_T_97) begin
        if (_T_98) begin
          if (_T_154) begin
            if (_T_293) begin
              if (io_master_in_sync) begin
                slave_out2_r_trans_type <= io_master_in_trans_type;
              end else begin
                if (_T_97) begin
                  if (_T_100) begin
                    if (_T_154) begin
                      if (_T_293) begin
                        if (io_master_in_sync) begin
                          slave_out2_r_trans_type <= io_master_in_trans_type;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_97) begin
                if (_T_100) begin
                  if (_T_154) begin
                    if (_T_293) begin
                      if (io_master_in_sync) begin
                        slave_out2_r_trans_type <= io_master_in_trans_type;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_97) begin
              if (_T_100) begin
                if (_T_154) begin
                  if (_T_293) begin
                    if (io_master_in_sync) begin
                      slave_out2_r_trans_type <= io_master_in_trans_type;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_97) begin
            if (_T_100) begin
              if (_T_154) begin
                if (_T_293) begin
                  if (io_master_in_sync) begin
                    slave_out2_r_trans_type <= io_master_in_trans_type;
                  end
                end
              end
            end
          end
        end
      end else begin
        slave_out2_r_trans_type <= _GEN_716;
      end
    end
    if (!(reset)) begin
      if (_T_97) begin
        if (_T_98) begin
          if (_T_163) begin
            if (_T_345) begin
              if (io_master_in_sync) begin
                slave_out3_r_addr <= _T_349;
              end else begin
                if (_T_97) begin
                  if (_T_100) begin
                    if (_T_163) begin
                      if (_T_345) begin
                        if (io_master_in_sync) begin
                          slave_out3_r_addr <= _T_349;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_97) begin
                if (_T_100) begin
                  if (_T_163) begin
                    if (_T_345) begin
                      if (io_master_in_sync) begin
                        slave_out3_r_addr <= _T_349;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_97) begin
              if (_T_100) begin
                if (_T_163) begin
                  if (_T_345) begin
                    if (io_master_in_sync) begin
                      slave_out3_r_addr <= _T_349;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_97) begin
            if (_T_100) begin
              if (_T_163) begin
                if (_T_345) begin
                  if (io_master_in_sync) begin
                    slave_out3_r_addr <= _T_349;
                  end
                end
              end
            end
          end
        end
      end else begin
        slave_out3_r_addr <= _GEN_904;
      end
    end
    if (!(reset)) begin
      if (_T_97) begin
        if (_T_98) begin
          if (_T_163) begin
            if (_T_345) begin
              if (io_master_in_sync) begin
                slave_out3_r_data <= 32'sh0;
              end else begin
                if (_T_97) begin
                  if (_T_100) begin
                    if (_T_163) begin
                      if (_T_345) begin
                        if (io_master_in_sync) begin
                          slave_out3_r_data <= io_master_in_data;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_97) begin
                if (_T_100) begin
                  if (_T_163) begin
                    if (_T_345) begin
                      if (io_master_in_sync) begin
                        slave_out3_r_data <= io_master_in_data;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_97) begin
              if (_T_100) begin
                if (_T_163) begin
                  if (_T_345) begin
                    if (io_master_in_sync) begin
                      slave_out3_r_data <= io_master_in_data;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_97) begin
            if (_T_100) begin
              if (_T_163) begin
                if (_T_345) begin
                  if (io_master_in_sync) begin
                    slave_out3_r_data <= io_master_in_data;
                  end
                end
              end
            end
          end
        end
      end else begin
        slave_out3_r_data <= _GEN_905;
      end
    end
    if (!(reset)) begin
      if (_T_97) begin
        if (_T_98) begin
          if (_T_163) begin
            if (_T_345) begin
              if (io_master_in_sync) begin
                slave_out3_r_trans_type <= io_master_in_trans_type;
              end else begin
                if (_T_97) begin
                  if (_T_100) begin
                    if (_T_163) begin
                      if (_T_345) begin
                        if (io_master_in_sync) begin
                          slave_out3_r_trans_type <= io_master_in_trans_type;
                        end
                      end
                    end
                  end
                end
              end
            end else begin
              if (_T_97) begin
                if (_T_100) begin
                  if (_T_163) begin
                    if (_T_345) begin
                      if (io_master_in_sync) begin
                        slave_out3_r_trans_type <= io_master_in_trans_type;
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_97) begin
              if (_T_100) begin
                if (_T_163) begin
                  if (_T_345) begin
                    if (io_master_in_sync) begin
                      slave_out3_r_trans_type <= io_master_in_trans_type;
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_97) begin
            if (_T_100) begin
              if (_T_163) begin
                if (_T_345) begin
                  if (io_master_in_sync) begin
                    slave_out3_r_trans_type <= io_master_in_trans_type;
                  end
                end
              end
            end
          end
        end
      end else begin
        slave_out3_r_trans_type <= _GEN_906;
      end
    end
    if (reset) begin
      req_signal_r_addr <= 32'sh0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (!(io_slave_in3_sync)) begin
            if (_T_529) begin
              if (_T_404) begin
                if (!(io_slave_in3_sync)) begin
                  if (_T_518) begin
                    if (!(io_slave_out3_sync)) begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (!(io_slave_in2_sync)) begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (!(io_slave_in2_sync)) begin
                                  if (_T_479) begin
                                    if (!(io_slave_out2_sync)) begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (!(io_slave_in1_sync)) begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (!(io_slave_in1_sync)) begin
                                                  if (_T_440) begin
                                                    if (!(io_slave_out1_sync)) begin
                                                      if (_T_429) begin
                                                        if (!(io_master_out_sync)) begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (!(io_slave_in0_sync)) begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (!(io_slave_in0_sync)) begin
                                                                      if (_T_390) begin
                                                                        if (!(io_slave_out0_sync)) begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    req_signal_r_addr <= _T_349;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              req_signal_r_addr <= _T_349;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        req_signal_r_addr <= _T_297;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  req_signal_r_addr <= _T_297;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            req_signal_r_addr <= _T_245;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      req_signal_r_addr <= _T_245;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    req_signal_r_addr <= _GEN_77;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                                        end else begin
                                                                                                                                                                          req_signal_r_addr <= _GEN_77;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        req_signal_r_addr <= _GEN_77;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      req_signal_r_addr <= _GEN_77;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    req_signal_r_addr <= _GEN_77;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  req_signal_r_addr <= _GEN_77;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                                      end else begin
                                                                                                                                                                        req_signal_r_addr <= _GEN_77;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      req_signal_r_addr <= _GEN_77;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    req_signal_r_addr <= _GEN_77;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  req_signal_r_addr <= _GEN_77;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                req_signal_r_addr <= _GEN_77;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                                    end else begin
                                                                                                                                                                      req_signal_r_addr <= _GEN_77;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    req_signal_r_addr <= _GEN_77;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  req_signal_r_addr <= _GEN_77;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                req_signal_r_addr <= _GEN_77;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              req_signal_r_addr <= _GEN_77;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          req_signal_r_addr <= _GEN_172;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        req_signal_r_addr <= _GEN_172;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      req_signal_r_addr <= _GEN_172;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                              end else begin
                                                                                                                                                                req_signal_r_addr <= _GEN_172;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              req_signal_r_addr <= _GEN_172;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            req_signal_r_addr <= _GEN_172;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          req_signal_r_addr <= _GEN_172;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        req_signal_r_addr <= _GEN_172;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      req_signal_r_addr <= _GEN_172;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    req_signal_r_addr <= _GEN_172;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                            end else begin
                                                                                                                                                              req_signal_r_addr <= _GEN_172;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            req_signal_r_addr <= _GEN_172;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          req_signal_r_addr <= _GEN_172;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        req_signal_r_addr <= _GEN_172;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      req_signal_r_addr <= _GEN_172;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    req_signal_r_addr <= _GEN_172;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  req_signal_r_addr <= _GEN_172;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                          end else begin
                                                                                                                                                            req_signal_r_addr <= _GEN_172;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          req_signal_r_addr <= _GEN_172;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        req_signal_r_addr <= _GEN_172;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      req_signal_r_addr <= _GEN_172;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    req_signal_r_addr <= _GEN_172;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  req_signal_r_addr <= _GEN_172;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                req_signal_r_addr <= _GEN_172;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            req_signal_r_addr <= _GEN_301;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          req_signal_r_addr <= _GEN_301;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        req_signal_r_addr <= _GEN_301;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  req_signal_r_addr <= io_master_in_addr;
                                                                                                                                                end else begin
                                                                                                                                                  req_signal_r_addr <= _GEN_301;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                req_signal_r_addr <= _GEN_301;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              req_signal_r_addr <= _GEN_301;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            req_signal_r_addr <= _GEN_301;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          req_signal_r_addr <= _GEN_301;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        req_signal_r_addr <= _GEN_301;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      req_signal_r_addr <= _GEN_301;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                req_signal_r_addr <= io_master_in_addr;
                                                                                                                                              end else begin
                                                                                                                                                req_signal_r_addr <= _GEN_301;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              req_signal_r_addr <= _GEN_301;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            req_signal_r_addr <= _GEN_301;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          req_signal_r_addr <= _GEN_301;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        req_signal_r_addr <= _GEN_301;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      req_signal_r_addr <= _GEN_301;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    req_signal_r_addr <= _GEN_301;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              req_signal_r_addr <= io_master_in_addr;
                                                                                                                                            end else begin
                                                                                                                                              req_signal_r_addr <= _GEN_301;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            req_signal_r_addr <= _GEN_301;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          req_signal_r_addr <= _GEN_301;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        req_signal_r_addr <= _GEN_301;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      req_signal_r_addr <= _GEN_301;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    req_signal_r_addr <= _GEN_301;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  req_signal_r_addr <= _GEN_301;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              req_signal_r_addr <= _GEN_427;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    req_signal_r_addr <= _T_245;
                                                                                                                                  end else begin
                                                                                                                                    req_signal_r_addr <= _GEN_427;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  req_signal_r_addr <= _GEN_427;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                req_signal_r_addr <= _GEN_427;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              req_signal_r_addr <= _GEN_427;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            req_signal_r_addr <= _GEN_427;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  req_signal_r_addr <= _T_245;
                                                                                                                                end else begin
                                                                                                                                  req_signal_r_addr <= _GEN_427;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                req_signal_r_addr <= _GEN_427;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              req_signal_r_addr <= _GEN_427;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            req_signal_r_addr <= _GEN_427;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          req_signal_r_addr <= _GEN_427;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                req_signal_r_addr <= _T_245;
                                                                                                                              end else begin
                                                                                                                                req_signal_r_addr <= _GEN_427;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              req_signal_r_addr <= _GEN_427;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            req_signal_r_addr <= _GEN_427;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          req_signal_r_addr <= _GEN_427;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        req_signal_r_addr <= _GEN_427;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    req_signal_r_addr <= _GEN_519;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          req_signal_r_addr <= _T_245;
                                                                                                                        end else begin
                                                                                                                          req_signal_r_addr <= _GEN_519;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        req_signal_r_addr <= _GEN_519;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      req_signal_r_addr <= _GEN_519;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    req_signal_r_addr <= _GEN_519;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  req_signal_r_addr <= _GEN_519;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        req_signal_r_addr <= _T_245;
                                                                                                                      end else begin
                                                                                                                        req_signal_r_addr <= _GEN_519;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      req_signal_r_addr <= _GEN_519;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    req_signal_r_addr <= _GEN_519;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  req_signal_r_addr <= _GEN_519;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                req_signal_r_addr <= _GEN_519;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      req_signal_r_addr <= _T_245;
                                                                                                                    end else begin
                                                                                                                      req_signal_r_addr <= _GEN_519;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    req_signal_r_addr <= _GEN_519;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  req_signal_r_addr <= _GEN_519;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                req_signal_r_addr <= _GEN_519;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              req_signal_r_addr <= _GEN_519;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          req_signal_r_addr <= _GEN_614;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                req_signal_r_addr <= _T_297;
                                                                                                              end else begin
                                                                                                                req_signal_r_addr <= _GEN_614;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              req_signal_r_addr <= _GEN_614;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            req_signal_r_addr <= _GEN_614;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          req_signal_r_addr <= _GEN_614;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        req_signal_r_addr <= _GEN_614;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              req_signal_r_addr <= _T_297;
                                                                                                            end else begin
                                                                                                              req_signal_r_addr <= _GEN_614;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            req_signal_r_addr <= _GEN_614;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          req_signal_r_addr <= _GEN_614;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        req_signal_r_addr <= _GEN_614;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      req_signal_r_addr <= _GEN_614;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            req_signal_r_addr <= _T_297;
                                                                                                          end else begin
                                                                                                            req_signal_r_addr <= _GEN_614;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          req_signal_r_addr <= _GEN_614;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        req_signal_r_addr <= _GEN_614;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      req_signal_r_addr <= _GEN_614;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    req_signal_r_addr <= _GEN_614;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                req_signal_r_addr <= _GEN_709;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      req_signal_r_addr <= _T_297;
                                                                                                    end else begin
                                                                                                      req_signal_r_addr <= _GEN_709;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    req_signal_r_addr <= _GEN_709;
                                                                                                  end
                                                                                                end else begin
                                                                                                  req_signal_r_addr <= _GEN_709;
                                                                                                end
                                                                                              end else begin
                                                                                                req_signal_r_addr <= _GEN_709;
                                                                                              end
                                                                                            end else begin
                                                                                              req_signal_r_addr <= _GEN_709;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    req_signal_r_addr <= _T_297;
                                                                                                  end else begin
                                                                                                    req_signal_r_addr <= _GEN_709;
                                                                                                  end
                                                                                                end else begin
                                                                                                  req_signal_r_addr <= _GEN_709;
                                                                                                end
                                                                                              end else begin
                                                                                                req_signal_r_addr <= _GEN_709;
                                                                                              end
                                                                                            end else begin
                                                                                              req_signal_r_addr <= _GEN_709;
                                                                                            end
                                                                                          end else begin
                                                                                            req_signal_r_addr <= _GEN_709;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  req_signal_r_addr <= _T_297;
                                                                                                end else begin
                                                                                                  req_signal_r_addr <= _GEN_709;
                                                                                                end
                                                                                              end else begin
                                                                                                req_signal_r_addr <= _GEN_709;
                                                                                              end
                                                                                            end else begin
                                                                                              req_signal_r_addr <= _GEN_709;
                                                                                            end
                                                                                          end else begin
                                                                                            req_signal_r_addr <= _GEN_709;
                                                                                          end
                                                                                        end else begin
                                                                                          req_signal_r_addr <= _GEN_709;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      req_signal_r_addr <= _GEN_804;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            req_signal_r_addr <= _T_349;
                                                                                          end else begin
                                                                                            req_signal_r_addr <= _GEN_804;
                                                                                          end
                                                                                        end else begin
                                                                                          req_signal_r_addr <= _GEN_804;
                                                                                        end
                                                                                      end else begin
                                                                                        req_signal_r_addr <= _GEN_804;
                                                                                      end
                                                                                    end else begin
                                                                                      req_signal_r_addr <= _GEN_804;
                                                                                    end
                                                                                  end else begin
                                                                                    req_signal_r_addr <= _GEN_804;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          req_signal_r_addr <= _T_349;
                                                                                        end else begin
                                                                                          req_signal_r_addr <= _GEN_804;
                                                                                        end
                                                                                      end else begin
                                                                                        req_signal_r_addr <= _GEN_804;
                                                                                      end
                                                                                    end else begin
                                                                                      req_signal_r_addr <= _GEN_804;
                                                                                    end
                                                                                  end else begin
                                                                                    req_signal_r_addr <= _GEN_804;
                                                                                  end
                                                                                end else begin
                                                                                  req_signal_r_addr <= _GEN_804;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        req_signal_r_addr <= _T_349;
                                                                                      end else begin
                                                                                        req_signal_r_addr <= _GEN_804;
                                                                                      end
                                                                                    end else begin
                                                                                      req_signal_r_addr <= _GEN_804;
                                                                                    end
                                                                                  end else begin
                                                                                    req_signal_r_addr <= _GEN_804;
                                                                                  end
                                                                                end else begin
                                                                                  req_signal_r_addr <= _GEN_804;
                                                                                end
                                                                              end else begin
                                                                                req_signal_r_addr <= _GEN_804;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            req_signal_r_addr <= _GEN_899;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  req_signal_r_addr <= _T_349;
                                                                                end else begin
                                                                                  req_signal_r_addr <= _GEN_899;
                                                                                end
                                                                              end else begin
                                                                                req_signal_r_addr <= _GEN_899;
                                                                              end
                                                                            end else begin
                                                                              req_signal_r_addr <= _GEN_899;
                                                                            end
                                                                          end else begin
                                                                            req_signal_r_addr <= _GEN_899;
                                                                          end
                                                                        end else begin
                                                                          req_signal_r_addr <= _GEN_899;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (!(io_slave_out0_sync)) begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  req_signal_r_addr <= _T_349;
                                                                                end else begin
                                                                                  req_signal_r_addr <= _GEN_899;
                                                                                end
                                                                              end else begin
                                                                                req_signal_r_addr <= _GEN_899;
                                                                              end
                                                                            end else begin
                                                                              req_signal_r_addr <= _GEN_899;
                                                                            end
                                                                          end else begin
                                                                            req_signal_r_addr <= _GEN_899;
                                                                          end
                                                                        end else begin
                                                                          req_signal_r_addr <= _GEN_899;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                req_signal_r_addr <= _T_349;
                                                                              end else begin
                                                                                req_signal_r_addr <= _GEN_899;
                                                                              end
                                                                            end else begin
                                                                              req_signal_r_addr <= _GEN_899;
                                                                            end
                                                                          end else begin
                                                                            req_signal_r_addr <= _GEN_899;
                                                                          end
                                                                        end else begin
                                                                          req_signal_r_addr <= _GEN_899;
                                                                        end
                                                                      end else begin
                                                                        req_signal_r_addr <= _GEN_899;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (!(io_slave_out0_sync)) begin
                                                                      req_signal_r_addr <= _GEN_994;
                                                                    end
                                                                  end else begin
                                                                    req_signal_r_addr <= _GEN_994;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (!(io_slave_in0_sync)) begin
                                                                    if (_T_390) begin
                                                                      if (!(io_slave_out0_sync)) begin
                                                                        req_signal_r_addr <= _GEN_994;
                                                                      end
                                                                    end else begin
                                                                      req_signal_r_addr <= _GEN_994;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  req_signal_r_addr <= _GEN_1029;
                                                                end
                                                              end else begin
                                                                req_signal_r_addr <= _GEN_1029;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (!(io_slave_in0_sync)) begin
                                                                  req_signal_r_addr <= _GEN_1029;
                                                                end
                                                              end else begin
                                                                req_signal_r_addr <= _GEN_1029;
                                                              end
                                                            end else begin
                                                              req_signal_r_addr <= _GEN_1029;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (!(io_slave_in0_sync)) begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (!(io_slave_in0_sync)) begin
                                                                    req_signal_r_addr <= _GEN_1029;
                                                                  end
                                                                end else begin
                                                                  req_signal_r_addr <= _GEN_1029;
                                                                end
                                                              end else begin
                                                                req_signal_r_addr <= _GEN_1029;
                                                              end
                                                            end
                                                          end else begin
                                                            req_signal_r_addr <= _GEN_1083;
                                                          end
                                                        end else begin
                                                          req_signal_r_addr <= _GEN_1083;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (!(io_master_out_sync)) begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (!(io_slave_in0_sync)) begin
                                                              req_signal_r_addr <= _GEN_1083;
                                                            end
                                                          end else begin
                                                            req_signal_r_addr <= _GEN_1083;
                                                          end
                                                        end else begin
                                                          req_signal_r_addr <= _GEN_1083;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (!(io_slave_in0_sync)) begin
                                                            req_signal_r_addr <= _GEN_1083;
                                                          end
                                                        end else begin
                                                          req_signal_r_addr <= _GEN_1083;
                                                        end
                                                      end else begin
                                                        req_signal_r_addr <= _GEN_1083;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (!(io_slave_out1_sync)) begin
                                                    if (_T_429) begin
                                                      if (!(io_master_out_sync)) begin
                                                        req_signal_r_addr <= _GEN_1137;
                                                      end
                                                    end else begin
                                                      req_signal_r_addr <= _GEN_1137;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (!(io_master_out_sync)) begin
                                                      req_signal_r_addr <= _GEN_1137;
                                                    end
                                                  end else begin
                                                    req_signal_r_addr <= _GEN_1137;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (!(io_slave_out1_sync)) begin
                                                  req_signal_r_addr <= _GEN_1169;
                                                end
                                              end else begin
                                                req_signal_r_addr <= _GEN_1169;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (!(io_slave_in1_sync)) begin
                                                if (_T_440) begin
                                                  if (!(io_slave_out1_sync)) begin
                                                    req_signal_r_addr <= _GEN_1169;
                                                  end
                                                end else begin
                                                  req_signal_r_addr <= _GEN_1169;
                                                end
                                              end
                                            end else begin
                                              req_signal_r_addr <= _GEN_1201;
                                            end
                                          end else begin
                                            req_signal_r_addr <= _GEN_1201;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (!(io_slave_in1_sync)) begin
                                              req_signal_r_addr <= _GEN_1201;
                                            end
                                          end else begin
                                            req_signal_r_addr <= _GEN_1201;
                                          end
                                        end else begin
                                          req_signal_r_addr <= _GEN_1201;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (!(io_slave_in1_sync)) begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (!(io_slave_in1_sync)) begin
                                                req_signal_r_addr <= _GEN_1201;
                                              end
                                            end else begin
                                              req_signal_r_addr <= _GEN_1201;
                                            end
                                          end else begin
                                            req_signal_r_addr <= _GEN_1201;
                                          end
                                        end
                                      end else begin
                                        req_signal_r_addr <= _GEN_1255;
                                      end
                                    end else begin
                                      req_signal_r_addr <= _GEN_1255;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (!(io_slave_out2_sync)) begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (!(io_slave_in1_sync)) begin
                                          req_signal_r_addr <= _GEN_1255;
                                        end
                                      end else begin
                                        req_signal_r_addr <= _GEN_1255;
                                      end
                                    end else begin
                                      req_signal_r_addr <= _GEN_1255;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (!(io_slave_in1_sync)) begin
                                        req_signal_r_addr <= _GEN_1255;
                                      end
                                    end else begin
                                      req_signal_r_addr <= _GEN_1255;
                                    end
                                  end else begin
                                    req_signal_r_addr <= _GEN_1255;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (!(io_slave_out2_sync)) begin
                                  req_signal_r_addr <= _GEN_1309;
                                end
                              end else begin
                                req_signal_r_addr <= _GEN_1309;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (!(io_slave_in2_sync)) begin
                                if (_T_479) begin
                                  if (!(io_slave_out2_sync)) begin
                                    req_signal_r_addr <= _GEN_1309;
                                  end
                                end else begin
                                  req_signal_r_addr <= _GEN_1309;
                                end
                              end
                            end else begin
                              req_signal_r_addr <= _GEN_1341;
                            end
                          end else begin
                            req_signal_r_addr <= _GEN_1341;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (!(io_slave_in2_sync)) begin
                              req_signal_r_addr <= _GEN_1341;
                            end
                          end else begin
                            req_signal_r_addr <= _GEN_1341;
                          end
                        end else begin
                          req_signal_r_addr <= _GEN_1341;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (!(io_slave_in2_sync)) begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (!(io_slave_in2_sync)) begin
                                req_signal_r_addr <= _GEN_1341;
                              end
                            end else begin
                              req_signal_r_addr <= _GEN_1341;
                            end
                          end else begin
                            req_signal_r_addr <= _GEN_1341;
                          end
                        end
                      end else begin
                        req_signal_r_addr <= _GEN_1395;
                      end
                    end else begin
                      req_signal_r_addr <= _GEN_1395;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (!(io_slave_out3_sync)) begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (!(io_slave_in2_sync)) begin
                          req_signal_r_addr <= _GEN_1395;
                        end
                      end else begin
                        req_signal_r_addr <= _GEN_1395;
                      end
                    end else begin
                      req_signal_r_addr <= _GEN_1395;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (!(io_slave_in2_sync)) begin
                        req_signal_r_addr <= _GEN_1395;
                      end
                    end else begin
                      req_signal_r_addr <= _GEN_1395;
                    end
                  end else begin
                    req_signal_r_addr <= _GEN_1395;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (!(io_slave_out3_sync)) begin
                  req_signal_r_addr <= _GEN_1449;
                end
              end else begin
                req_signal_r_addr <= _GEN_1449;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (!(io_slave_in3_sync)) begin
                if (_T_518) begin
                  if (!(io_slave_out3_sync)) begin
                    req_signal_r_addr <= _GEN_1449;
                  end
                end else begin
                  req_signal_r_addr <= _GEN_1449;
                end
              end
            end else begin
              req_signal_r_addr <= _GEN_1481;
            end
          end else begin
            req_signal_r_addr <= _GEN_1481;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (!(io_slave_in3_sync)) begin
              req_signal_r_addr <= _GEN_1481;
            end
          end else begin
            req_signal_r_addr <= _GEN_1481;
          end
        end else begin
          req_signal_r_addr <= _GEN_1481;
        end
      end
    end
    if (reset) begin
      req_signal_r_data <= 32'sh0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (!(io_slave_in3_sync)) begin
            if (_T_529) begin
              if (_T_404) begin
                if (!(io_slave_in3_sync)) begin
                  if (_T_518) begin
                    if (!(io_slave_out3_sync)) begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (!(io_slave_in2_sync)) begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (!(io_slave_in2_sync)) begin
                                  if (_T_479) begin
                                    if (!(io_slave_out2_sync)) begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (!(io_slave_in1_sync)) begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (!(io_slave_in1_sync)) begin
                                                  if (_T_440) begin
                                                    if (!(io_slave_out1_sync)) begin
                                                      if (_T_429) begin
                                                        if (!(io_master_out_sync)) begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (!(io_slave_in0_sync)) begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (!(io_slave_in0_sync)) begin
                                                                      if (_T_390) begin
                                                                        if (!(io_slave_out0_sync)) begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    req_signal_r_data <= 32'sh0;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              req_signal_r_data <= io_master_in_data;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        req_signal_r_data <= 32'sh0;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  req_signal_r_data <= io_master_in_data;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            req_signal_r_data <= 32'sh0;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      req_signal_r_data <= io_master_in_data;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    req_signal_r_data <= io_master_in_data;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  req_signal_r_data <= 32'sh0;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            req_signal_r_data <= 32'sh0;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      req_signal_r_data <= io_master_in_data;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    req_signal_r_data <= io_master_in_data;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  req_signal_r_data <= io_master_in_data;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                req_signal_r_data <= io_master_in_data;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    req_signal_r_data <= _GEN_78;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          req_signal_r_data <= 32'sh0;
                                                                                                                                                                        end else begin
                                                                                                                                                                          req_signal_r_data <= _GEN_78;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        req_signal_r_data <= _GEN_78;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      req_signal_r_data <= _GEN_78;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    req_signal_r_data <= _GEN_78;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  req_signal_r_data <= _GEN_78;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        req_signal_r_data <= 32'sh0;
                                                                                                                                                                      end else begin
                                                                                                                                                                        req_signal_r_data <= _GEN_78;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      req_signal_r_data <= _GEN_78;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    req_signal_r_data <= _GEN_78;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  req_signal_r_data <= _GEN_78;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                req_signal_r_data <= _GEN_78;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      req_signal_r_data <= 32'sh0;
                                                                                                                                                                    end else begin
                                                                                                                                                                      req_signal_r_data <= _GEN_78;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    req_signal_r_data <= _GEN_78;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  req_signal_r_data <= _GEN_78;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                req_signal_r_data <= _GEN_78;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              req_signal_r_data <= _GEN_78;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          req_signal_r_data <= _GEN_173;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        req_signal_r_data <= _GEN_173;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      req_signal_r_data <= _GEN_173;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                req_signal_r_data <= 32'sh0;
                                                                                                                                                              end else begin
                                                                                                                                                                req_signal_r_data <= _GEN_173;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              req_signal_r_data <= _GEN_173;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            req_signal_r_data <= _GEN_173;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          req_signal_r_data <= _GEN_173;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        req_signal_r_data <= _GEN_173;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      req_signal_r_data <= _GEN_173;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    req_signal_r_data <= _GEN_173;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              req_signal_r_data <= 32'sh0;
                                                                                                                                                            end else begin
                                                                                                                                                              req_signal_r_data <= _GEN_173;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            req_signal_r_data <= _GEN_173;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          req_signal_r_data <= _GEN_173;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        req_signal_r_data <= _GEN_173;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      req_signal_r_data <= _GEN_173;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    req_signal_r_data <= _GEN_173;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  req_signal_r_data <= _GEN_173;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            req_signal_r_data <= 32'sh0;
                                                                                                                                                          end else begin
                                                                                                                                                            req_signal_r_data <= _GEN_173;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          req_signal_r_data <= _GEN_173;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        req_signal_r_data <= _GEN_173;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      req_signal_r_data <= _GEN_173;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    req_signal_r_data <= _GEN_173;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  req_signal_r_data <= _GEN_173;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                req_signal_r_data <= _GEN_173;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            req_signal_r_data <= _GEN_302;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          req_signal_r_data <= _GEN_302;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        req_signal_r_data <= _GEN_302;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  req_signal_r_data <= io_master_in_data;
                                                                                                                                                end else begin
                                                                                                                                                  req_signal_r_data <= _GEN_302;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                req_signal_r_data <= _GEN_302;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              req_signal_r_data <= _GEN_302;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            req_signal_r_data <= _GEN_302;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          req_signal_r_data <= _GEN_302;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        req_signal_r_data <= _GEN_302;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      req_signal_r_data <= _GEN_302;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                req_signal_r_data <= io_master_in_data;
                                                                                                                                              end else begin
                                                                                                                                                req_signal_r_data <= _GEN_302;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              req_signal_r_data <= _GEN_302;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            req_signal_r_data <= _GEN_302;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          req_signal_r_data <= _GEN_302;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        req_signal_r_data <= _GEN_302;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      req_signal_r_data <= _GEN_302;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    req_signal_r_data <= _GEN_302;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              req_signal_r_data <= io_master_in_data;
                                                                                                                                            end else begin
                                                                                                                                              req_signal_r_data <= _GEN_302;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            req_signal_r_data <= _GEN_302;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          req_signal_r_data <= _GEN_302;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        req_signal_r_data <= _GEN_302;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      req_signal_r_data <= _GEN_302;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    req_signal_r_data <= _GEN_302;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  req_signal_r_data <= _GEN_302;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              req_signal_r_data <= _GEN_428;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    req_signal_r_data <= io_master_in_data;
                                                                                                                                  end else begin
                                                                                                                                    req_signal_r_data <= _GEN_428;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  req_signal_r_data <= _GEN_428;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                req_signal_r_data <= _GEN_428;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              req_signal_r_data <= _GEN_428;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            req_signal_r_data <= _GEN_428;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  req_signal_r_data <= io_master_in_data;
                                                                                                                                end else begin
                                                                                                                                  req_signal_r_data <= _GEN_428;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                req_signal_r_data <= _GEN_428;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              req_signal_r_data <= _GEN_428;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            req_signal_r_data <= _GEN_428;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          req_signal_r_data <= _GEN_428;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                req_signal_r_data <= io_master_in_data;
                                                                                                                              end else begin
                                                                                                                                req_signal_r_data <= _GEN_428;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              req_signal_r_data <= _GEN_428;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            req_signal_r_data <= _GEN_428;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          req_signal_r_data <= _GEN_428;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        req_signal_r_data <= _GEN_428;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    req_signal_r_data <= _GEN_520;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          req_signal_r_data <= 32'sh0;
                                                                                                                        end else begin
                                                                                                                          req_signal_r_data <= _GEN_520;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        req_signal_r_data <= _GEN_520;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      req_signal_r_data <= _GEN_520;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    req_signal_r_data <= _GEN_520;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  req_signal_r_data <= _GEN_520;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        req_signal_r_data <= 32'sh0;
                                                                                                                      end else begin
                                                                                                                        req_signal_r_data <= _GEN_520;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      req_signal_r_data <= _GEN_520;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    req_signal_r_data <= _GEN_520;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  req_signal_r_data <= _GEN_520;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                req_signal_r_data <= _GEN_520;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      req_signal_r_data <= 32'sh0;
                                                                                                                    end else begin
                                                                                                                      req_signal_r_data <= _GEN_520;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    req_signal_r_data <= _GEN_520;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  req_signal_r_data <= _GEN_520;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                req_signal_r_data <= _GEN_520;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              req_signal_r_data <= _GEN_520;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          req_signal_r_data <= _GEN_615;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                req_signal_r_data <= io_master_in_data;
                                                                                                              end else begin
                                                                                                                req_signal_r_data <= _GEN_615;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              req_signal_r_data <= _GEN_615;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            req_signal_r_data <= _GEN_615;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          req_signal_r_data <= _GEN_615;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        req_signal_r_data <= _GEN_615;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              req_signal_r_data <= io_master_in_data;
                                                                                                            end else begin
                                                                                                              req_signal_r_data <= _GEN_615;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            req_signal_r_data <= _GEN_615;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          req_signal_r_data <= _GEN_615;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        req_signal_r_data <= _GEN_615;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      req_signal_r_data <= _GEN_615;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            req_signal_r_data <= io_master_in_data;
                                                                                                          end else begin
                                                                                                            req_signal_r_data <= _GEN_615;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          req_signal_r_data <= _GEN_615;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        req_signal_r_data <= _GEN_615;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      req_signal_r_data <= _GEN_615;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    req_signal_r_data <= _GEN_615;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                req_signal_r_data <= _GEN_710;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      req_signal_r_data <= 32'sh0;
                                                                                                    end else begin
                                                                                                      req_signal_r_data <= _GEN_710;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    req_signal_r_data <= _GEN_710;
                                                                                                  end
                                                                                                end else begin
                                                                                                  req_signal_r_data <= _GEN_710;
                                                                                                end
                                                                                              end else begin
                                                                                                req_signal_r_data <= _GEN_710;
                                                                                              end
                                                                                            end else begin
                                                                                              req_signal_r_data <= _GEN_710;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    req_signal_r_data <= 32'sh0;
                                                                                                  end else begin
                                                                                                    req_signal_r_data <= _GEN_710;
                                                                                                  end
                                                                                                end else begin
                                                                                                  req_signal_r_data <= _GEN_710;
                                                                                                end
                                                                                              end else begin
                                                                                                req_signal_r_data <= _GEN_710;
                                                                                              end
                                                                                            end else begin
                                                                                              req_signal_r_data <= _GEN_710;
                                                                                            end
                                                                                          end else begin
                                                                                            req_signal_r_data <= _GEN_710;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  req_signal_r_data <= 32'sh0;
                                                                                                end else begin
                                                                                                  req_signal_r_data <= _GEN_710;
                                                                                                end
                                                                                              end else begin
                                                                                                req_signal_r_data <= _GEN_710;
                                                                                              end
                                                                                            end else begin
                                                                                              req_signal_r_data <= _GEN_710;
                                                                                            end
                                                                                          end else begin
                                                                                            req_signal_r_data <= _GEN_710;
                                                                                          end
                                                                                        end else begin
                                                                                          req_signal_r_data <= _GEN_710;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      req_signal_r_data <= _GEN_805;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            req_signal_r_data <= io_master_in_data;
                                                                                          end else begin
                                                                                            req_signal_r_data <= _GEN_805;
                                                                                          end
                                                                                        end else begin
                                                                                          req_signal_r_data <= _GEN_805;
                                                                                        end
                                                                                      end else begin
                                                                                        req_signal_r_data <= _GEN_805;
                                                                                      end
                                                                                    end else begin
                                                                                      req_signal_r_data <= _GEN_805;
                                                                                    end
                                                                                  end else begin
                                                                                    req_signal_r_data <= _GEN_805;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          req_signal_r_data <= io_master_in_data;
                                                                                        end else begin
                                                                                          req_signal_r_data <= _GEN_805;
                                                                                        end
                                                                                      end else begin
                                                                                        req_signal_r_data <= _GEN_805;
                                                                                      end
                                                                                    end else begin
                                                                                      req_signal_r_data <= _GEN_805;
                                                                                    end
                                                                                  end else begin
                                                                                    req_signal_r_data <= _GEN_805;
                                                                                  end
                                                                                end else begin
                                                                                  req_signal_r_data <= _GEN_805;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        req_signal_r_data <= io_master_in_data;
                                                                                      end else begin
                                                                                        req_signal_r_data <= _GEN_805;
                                                                                      end
                                                                                    end else begin
                                                                                      req_signal_r_data <= _GEN_805;
                                                                                    end
                                                                                  end else begin
                                                                                    req_signal_r_data <= _GEN_805;
                                                                                  end
                                                                                end else begin
                                                                                  req_signal_r_data <= _GEN_805;
                                                                                end
                                                                              end else begin
                                                                                req_signal_r_data <= _GEN_805;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            req_signal_r_data <= _GEN_900;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  req_signal_r_data <= 32'sh0;
                                                                                end else begin
                                                                                  req_signal_r_data <= _GEN_900;
                                                                                end
                                                                              end else begin
                                                                                req_signal_r_data <= _GEN_900;
                                                                              end
                                                                            end else begin
                                                                              req_signal_r_data <= _GEN_900;
                                                                            end
                                                                          end else begin
                                                                            req_signal_r_data <= _GEN_900;
                                                                          end
                                                                        end else begin
                                                                          req_signal_r_data <= _GEN_900;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (!(io_slave_out0_sync)) begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  req_signal_r_data <= 32'sh0;
                                                                                end else begin
                                                                                  req_signal_r_data <= _GEN_900;
                                                                                end
                                                                              end else begin
                                                                                req_signal_r_data <= _GEN_900;
                                                                              end
                                                                            end else begin
                                                                              req_signal_r_data <= _GEN_900;
                                                                            end
                                                                          end else begin
                                                                            req_signal_r_data <= _GEN_900;
                                                                          end
                                                                        end else begin
                                                                          req_signal_r_data <= _GEN_900;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                req_signal_r_data <= 32'sh0;
                                                                              end else begin
                                                                                req_signal_r_data <= _GEN_900;
                                                                              end
                                                                            end else begin
                                                                              req_signal_r_data <= _GEN_900;
                                                                            end
                                                                          end else begin
                                                                            req_signal_r_data <= _GEN_900;
                                                                          end
                                                                        end else begin
                                                                          req_signal_r_data <= _GEN_900;
                                                                        end
                                                                      end else begin
                                                                        req_signal_r_data <= _GEN_900;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (!(io_slave_out0_sync)) begin
                                                                      req_signal_r_data <= _GEN_995;
                                                                    end
                                                                  end else begin
                                                                    req_signal_r_data <= _GEN_995;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (!(io_slave_in0_sync)) begin
                                                                    if (_T_390) begin
                                                                      if (!(io_slave_out0_sync)) begin
                                                                        req_signal_r_data <= _GEN_995;
                                                                      end
                                                                    end else begin
                                                                      req_signal_r_data <= _GEN_995;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  req_signal_r_data <= _GEN_1030;
                                                                end
                                                              end else begin
                                                                req_signal_r_data <= _GEN_1030;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (!(io_slave_in0_sync)) begin
                                                                  req_signal_r_data <= _GEN_1030;
                                                                end
                                                              end else begin
                                                                req_signal_r_data <= _GEN_1030;
                                                              end
                                                            end else begin
                                                              req_signal_r_data <= _GEN_1030;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (!(io_slave_in0_sync)) begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (!(io_slave_in0_sync)) begin
                                                                    req_signal_r_data <= _GEN_1030;
                                                                  end
                                                                end else begin
                                                                  req_signal_r_data <= _GEN_1030;
                                                                end
                                                              end else begin
                                                                req_signal_r_data <= _GEN_1030;
                                                              end
                                                            end
                                                          end else begin
                                                            req_signal_r_data <= _GEN_1084;
                                                          end
                                                        end else begin
                                                          req_signal_r_data <= _GEN_1084;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (!(io_master_out_sync)) begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (!(io_slave_in0_sync)) begin
                                                              req_signal_r_data <= _GEN_1084;
                                                            end
                                                          end else begin
                                                            req_signal_r_data <= _GEN_1084;
                                                          end
                                                        end else begin
                                                          req_signal_r_data <= _GEN_1084;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (!(io_slave_in0_sync)) begin
                                                            req_signal_r_data <= _GEN_1084;
                                                          end
                                                        end else begin
                                                          req_signal_r_data <= _GEN_1084;
                                                        end
                                                      end else begin
                                                        req_signal_r_data <= _GEN_1084;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (!(io_slave_out1_sync)) begin
                                                    if (_T_429) begin
                                                      if (!(io_master_out_sync)) begin
                                                        req_signal_r_data <= _GEN_1138;
                                                      end
                                                    end else begin
                                                      req_signal_r_data <= _GEN_1138;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (!(io_master_out_sync)) begin
                                                      req_signal_r_data <= _GEN_1138;
                                                    end
                                                  end else begin
                                                    req_signal_r_data <= _GEN_1138;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (!(io_slave_out1_sync)) begin
                                                  req_signal_r_data <= _GEN_1170;
                                                end
                                              end else begin
                                                req_signal_r_data <= _GEN_1170;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (!(io_slave_in1_sync)) begin
                                                if (_T_440) begin
                                                  if (!(io_slave_out1_sync)) begin
                                                    req_signal_r_data <= _GEN_1170;
                                                  end
                                                end else begin
                                                  req_signal_r_data <= _GEN_1170;
                                                end
                                              end
                                            end else begin
                                              req_signal_r_data <= _GEN_1202;
                                            end
                                          end else begin
                                            req_signal_r_data <= _GEN_1202;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (!(io_slave_in1_sync)) begin
                                              req_signal_r_data <= _GEN_1202;
                                            end
                                          end else begin
                                            req_signal_r_data <= _GEN_1202;
                                          end
                                        end else begin
                                          req_signal_r_data <= _GEN_1202;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (!(io_slave_in1_sync)) begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (!(io_slave_in1_sync)) begin
                                                req_signal_r_data <= _GEN_1202;
                                              end
                                            end else begin
                                              req_signal_r_data <= _GEN_1202;
                                            end
                                          end else begin
                                            req_signal_r_data <= _GEN_1202;
                                          end
                                        end
                                      end else begin
                                        req_signal_r_data <= _GEN_1256;
                                      end
                                    end else begin
                                      req_signal_r_data <= _GEN_1256;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (!(io_slave_out2_sync)) begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (!(io_slave_in1_sync)) begin
                                          req_signal_r_data <= _GEN_1256;
                                        end
                                      end else begin
                                        req_signal_r_data <= _GEN_1256;
                                      end
                                    end else begin
                                      req_signal_r_data <= _GEN_1256;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (!(io_slave_in1_sync)) begin
                                        req_signal_r_data <= _GEN_1256;
                                      end
                                    end else begin
                                      req_signal_r_data <= _GEN_1256;
                                    end
                                  end else begin
                                    req_signal_r_data <= _GEN_1256;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (!(io_slave_out2_sync)) begin
                                  req_signal_r_data <= _GEN_1310;
                                end
                              end else begin
                                req_signal_r_data <= _GEN_1310;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (!(io_slave_in2_sync)) begin
                                if (_T_479) begin
                                  if (!(io_slave_out2_sync)) begin
                                    req_signal_r_data <= _GEN_1310;
                                  end
                                end else begin
                                  req_signal_r_data <= _GEN_1310;
                                end
                              end
                            end else begin
                              req_signal_r_data <= _GEN_1342;
                            end
                          end else begin
                            req_signal_r_data <= _GEN_1342;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (!(io_slave_in2_sync)) begin
                              req_signal_r_data <= _GEN_1342;
                            end
                          end else begin
                            req_signal_r_data <= _GEN_1342;
                          end
                        end else begin
                          req_signal_r_data <= _GEN_1342;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (!(io_slave_in2_sync)) begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (!(io_slave_in2_sync)) begin
                                req_signal_r_data <= _GEN_1342;
                              end
                            end else begin
                              req_signal_r_data <= _GEN_1342;
                            end
                          end else begin
                            req_signal_r_data <= _GEN_1342;
                          end
                        end
                      end else begin
                        req_signal_r_data <= _GEN_1396;
                      end
                    end else begin
                      req_signal_r_data <= _GEN_1396;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (!(io_slave_out3_sync)) begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (!(io_slave_in2_sync)) begin
                          req_signal_r_data <= _GEN_1396;
                        end
                      end else begin
                        req_signal_r_data <= _GEN_1396;
                      end
                    end else begin
                      req_signal_r_data <= _GEN_1396;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (!(io_slave_in2_sync)) begin
                        req_signal_r_data <= _GEN_1396;
                      end
                    end else begin
                      req_signal_r_data <= _GEN_1396;
                    end
                  end else begin
                    req_signal_r_data <= _GEN_1396;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (!(io_slave_out3_sync)) begin
                  req_signal_r_data <= _GEN_1450;
                end
              end else begin
                req_signal_r_data <= _GEN_1450;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (!(io_slave_in3_sync)) begin
                if (_T_518) begin
                  if (!(io_slave_out3_sync)) begin
                    req_signal_r_data <= _GEN_1450;
                  end
                end else begin
                  req_signal_r_data <= _GEN_1450;
                end
              end
            end else begin
              req_signal_r_data <= _GEN_1482;
            end
          end else begin
            req_signal_r_data <= _GEN_1482;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (!(io_slave_in3_sync)) begin
              req_signal_r_data <= _GEN_1482;
            end
          end else begin
            req_signal_r_data <= _GEN_1482;
          end
        end else begin
          req_signal_r_data <= _GEN_1482;
        end
      end
    end
    if (reset) begin
      req_signal_r_trans_type <= 32'h0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (!(io_slave_in3_sync)) begin
            if (_T_529) begin
              if (_T_404) begin
                if (!(io_slave_in3_sync)) begin
                  if (_T_518) begin
                    if (!(io_slave_out3_sync)) begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (!(io_slave_in2_sync)) begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (!(io_slave_in2_sync)) begin
                                  if (_T_479) begin
                                    if (!(io_slave_out2_sync)) begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (!(io_slave_in1_sync)) begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (!(io_slave_in1_sync)) begin
                                                  if (_T_440) begin
                                                    if (!(io_slave_out1_sync)) begin
                                                      if (_T_429) begin
                                                        if (!(io_master_out_sync)) begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (!(io_slave_in0_sync)) begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (!(io_slave_in0_sync)) begin
                                                                      if (_T_390) begin
                                                                        if (!(io_slave_out0_sync)) begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                                        end else begin
                                                                                                                                                                          req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                                      end else begin
                                                                                                                                                                        req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                                    end else begin
                                                                                                                                                                      req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              req_signal_r_trans_type <= _GEN_79;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                              end else begin
                                                                                                                                                                req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                            end else begin
                                                                                                                                                              req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                          end else begin
                                                                                                                                                            req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  req_signal_r_trans_type <= _GEN_174;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                req_signal_r_trans_type <= _GEN_174;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            req_signal_r_trans_type <= _GEN_303;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          req_signal_r_trans_type <= _GEN_303;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        req_signal_r_trans_type <= _GEN_303;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                                end else begin
                                                                                                                                                  req_signal_r_trans_type <= _GEN_303;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                req_signal_r_trans_type <= _GEN_303;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              req_signal_r_trans_type <= _GEN_303;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            req_signal_r_trans_type <= _GEN_303;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          req_signal_r_trans_type <= _GEN_303;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        req_signal_r_trans_type <= _GEN_303;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      req_signal_r_trans_type <= _GEN_303;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                              end else begin
                                                                                                                                                req_signal_r_trans_type <= _GEN_303;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              req_signal_r_trans_type <= _GEN_303;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            req_signal_r_trans_type <= _GEN_303;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          req_signal_r_trans_type <= _GEN_303;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        req_signal_r_trans_type <= _GEN_303;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      req_signal_r_trans_type <= _GEN_303;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    req_signal_r_trans_type <= _GEN_303;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                            end else begin
                                                                                                                                              req_signal_r_trans_type <= _GEN_303;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            req_signal_r_trans_type <= _GEN_303;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          req_signal_r_trans_type <= _GEN_303;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        req_signal_r_trans_type <= _GEN_303;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      req_signal_r_trans_type <= _GEN_303;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    req_signal_r_trans_type <= _GEN_303;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  req_signal_r_trans_type <= _GEN_303;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              req_signal_r_trans_type <= _GEN_429;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                  end else begin
                                                                                                                                    req_signal_r_trans_type <= _GEN_429;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  req_signal_r_trans_type <= _GEN_429;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                req_signal_r_trans_type <= _GEN_429;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              req_signal_r_trans_type <= _GEN_429;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            req_signal_r_trans_type <= _GEN_429;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                                end else begin
                                                                                                                                  req_signal_r_trans_type <= _GEN_429;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                req_signal_r_trans_type <= _GEN_429;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              req_signal_r_trans_type <= _GEN_429;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            req_signal_r_trans_type <= _GEN_429;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          req_signal_r_trans_type <= _GEN_429;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                              end else begin
                                                                                                                                req_signal_r_trans_type <= _GEN_429;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              req_signal_r_trans_type <= _GEN_429;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            req_signal_r_trans_type <= _GEN_429;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          req_signal_r_trans_type <= _GEN_429;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        req_signal_r_trans_type <= _GEN_429;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    req_signal_r_trans_type <= _GEN_521;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                        end else begin
                                                                                                                          req_signal_r_trans_type <= _GEN_521;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        req_signal_r_trans_type <= _GEN_521;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      req_signal_r_trans_type <= _GEN_521;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    req_signal_r_trans_type <= _GEN_521;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  req_signal_r_trans_type <= _GEN_521;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                      end else begin
                                                                                                                        req_signal_r_trans_type <= _GEN_521;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      req_signal_r_trans_type <= _GEN_521;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    req_signal_r_trans_type <= _GEN_521;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  req_signal_r_trans_type <= _GEN_521;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                req_signal_r_trans_type <= _GEN_521;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                                    end else begin
                                                                                                                      req_signal_r_trans_type <= _GEN_521;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    req_signal_r_trans_type <= _GEN_521;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  req_signal_r_trans_type <= _GEN_521;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                req_signal_r_trans_type <= _GEN_521;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              req_signal_r_trans_type <= _GEN_521;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          req_signal_r_trans_type <= _GEN_616;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                              end else begin
                                                                                                                req_signal_r_trans_type <= _GEN_616;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              req_signal_r_trans_type <= _GEN_616;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            req_signal_r_trans_type <= _GEN_616;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          req_signal_r_trans_type <= _GEN_616;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        req_signal_r_trans_type <= _GEN_616;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                            end else begin
                                                                                                              req_signal_r_trans_type <= _GEN_616;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            req_signal_r_trans_type <= _GEN_616;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          req_signal_r_trans_type <= _GEN_616;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        req_signal_r_trans_type <= _GEN_616;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      req_signal_r_trans_type <= _GEN_616;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                          end else begin
                                                                                                            req_signal_r_trans_type <= _GEN_616;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          req_signal_r_trans_type <= _GEN_616;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        req_signal_r_trans_type <= _GEN_616;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      req_signal_r_trans_type <= _GEN_616;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    req_signal_r_trans_type <= _GEN_616;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                req_signal_r_trans_type <= _GEN_711;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                    end else begin
                                                                                                      req_signal_r_trans_type <= _GEN_711;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    req_signal_r_trans_type <= _GEN_711;
                                                                                                  end
                                                                                                end else begin
                                                                                                  req_signal_r_trans_type <= _GEN_711;
                                                                                                end
                                                                                              end else begin
                                                                                                req_signal_r_trans_type <= _GEN_711;
                                                                                              end
                                                                                            end else begin
                                                                                              req_signal_r_trans_type <= _GEN_711;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                  end else begin
                                                                                                    req_signal_r_trans_type <= _GEN_711;
                                                                                                  end
                                                                                                end else begin
                                                                                                  req_signal_r_trans_type <= _GEN_711;
                                                                                                end
                                                                                              end else begin
                                                                                                req_signal_r_trans_type <= _GEN_711;
                                                                                              end
                                                                                            end else begin
                                                                                              req_signal_r_trans_type <= _GEN_711;
                                                                                            end
                                                                                          end else begin
                                                                                            req_signal_r_trans_type <= _GEN_711;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                                end else begin
                                                                                                  req_signal_r_trans_type <= _GEN_711;
                                                                                                end
                                                                                              end else begin
                                                                                                req_signal_r_trans_type <= _GEN_711;
                                                                                              end
                                                                                            end else begin
                                                                                              req_signal_r_trans_type <= _GEN_711;
                                                                                            end
                                                                                          end else begin
                                                                                            req_signal_r_trans_type <= _GEN_711;
                                                                                          end
                                                                                        end else begin
                                                                                          req_signal_r_trans_type <= _GEN_711;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      req_signal_r_trans_type <= _GEN_806;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                          end else begin
                                                                                            req_signal_r_trans_type <= _GEN_806;
                                                                                          end
                                                                                        end else begin
                                                                                          req_signal_r_trans_type <= _GEN_806;
                                                                                        end
                                                                                      end else begin
                                                                                        req_signal_r_trans_type <= _GEN_806;
                                                                                      end
                                                                                    end else begin
                                                                                      req_signal_r_trans_type <= _GEN_806;
                                                                                    end
                                                                                  end else begin
                                                                                    req_signal_r_trans_type <= _GEN_806;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                        end else begin
                                                                                          req_signal_r_trans_type <= _GEN_806;
                                                                                        end
                                                                                      end else begin
                                                                                        req_signal_r_trans_type <= _GEN_806;
                                                                                      end
                                                                                    end else begin
                                                                                      req_signal_r_trans_type <= _GEN_806;
                                                                                    end
                                                                                  end else begin
                                                                                    req_signal_r_trans_type <= _GEN_806;
                                                                                  end
                                                                                end else begin
                                                                                  req_signal_r_trans_type <= _GEN_806;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                      end else begin
                                                                                        req_signal_r_trans_type <= _GEN_806;
                                                                                      end
                                                                                    end else begin
                                                                                      req_signal_r_trans_type <= _GEN_806;
                                                                                    end
                                                                                  end else begin
                                                                                    req_signal_r_trans_type <= _GEN_806;
                                                                                  end
                                                                                end else begin
                                                                                  req_signal_r_trans_type <= _GEN_806;
                                                                                end
                                                                              end else begin
                                                                                req_signal_r_trans_type <= _GEN_806;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            req_signal_r_trans_type <= _GEN_901;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                end else begin
                                                                                  req_signal_r_trans_type <= _GEN_901;
                                                                                end
                                                                              end else begin
                                                                                req_signal_r_trans_type <= _GEN_901;
                                                                              end
                                                                            end else begin
                                                                              req_signal_r_trans_type <= _GEN_901;
                                                                            end
                                                                          end else begin
                                                                            req_signal_r_trans_type <= _GEN_901;
                                                                          end
                                                                        end else begin
                                                                          req_signal_r_trans_type <= _GEN_901;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (!(io_slave_out0_sync)) begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  req_signal_r_trans_type <= io_master_in_trans_type;
                                                                                end else begin
                                                                                  req_signal_r_trans_type <= _GEN_901;
                                                                                end
                                                                              end else begin
                                                                                req_signal_r_trans_type <= _GEN_901;
                                                                              end
                                                                            end else begin
                                                                              req_signal_r_trans_type <= _GEN_901;
                                                                            end
                                                                          end else begin
                                                                            req_signal_r_trans_type <= _GEN_901;
                                                                          end
                                                                        end else begin
                                                                          req_signal_r_trans_type <= _GEN_901;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                req_signal_r_trans_type <= io_master_in_trans_type;
                                                                              end else begin
                                                                                req_signal_r_trans_type <= _GEN_901;
                                                                              end
                                                                            end else begin
                                                                              req_signal_r_trans_type <= _GEN_901;
                                                                            end
                                                                          end else begin
                                                                            req_signal_r_trans_type <= _GEN_901;
                                                                          end
                                                                        end else begin
                                                                          req_signal_r_trans_type <= _GEN_901;
                                                                        end
                                                                      end else begin
                                                                        req_signal_r_trans_type <= _GEN_901;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (!(io_slave_out0_sync)) begin
                                                                      req_signal_r_trans_type <= _GEN_996;
                                                                    end
                                                                  end else begin
                                                                    req_signal_r_trans_type <= _GEN_996;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (!(io_slave_in0_sync)) begin
                                                                    if (_T_390) begin
                                                                      if (!(io_slave_out0_sync)) begin
                                                                        req_signal_r_trans_type <= _GEN_996;
                                                                      end
                                                                    end else begin
                                                                      req_signal_r_trans_type <= _GEN_996;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  req_signal_r_trans_type <= _GEN_1031;
                                                                end
                                                              end else begin
                                                                req_signal_r_trans_type <= _GEN_1031;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (!(io_slave_in0_sync)) begin
                                                                  req_signal_r_trans_type <= _GEN_1031;
                                                                end
                                                              end else begin
                                                                req_signal_r_trans_type <= _GEN_1031;
                                                              end
                                                            end else begin
                                                              req_signal_r_trans_type <= _GEN_1031;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (!(io_slave_in0_sync)) begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (!(io_slave_in0_sync)) begin
                                                                    req_signal_r_trans_type <= _GEN_1031;
                                                                  end
                                                                end else begin
                                                                  req_signal_r_trans_type <= _GEN_1031;
                                                                end
                                                              end else begin
                                                                req_signal_r_trans_type <= _GEN_1031;
                                                              end
                                                            end
                                                          end else begin
                                                            req_signal_r_trans_type <= _GEN_1085;
                                                          end
                                                        end else begin
                                                          req_signal_r_trans_type <= _GEN_1085;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (!(io_master_out_sync)) begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (!(io_slave_in0_sync)) begin
                                                              req_signal_r_trans_type <= _GEN_1085;
                                                            end
                                                          end else begin
                                                            req_signal_r_trans_type <= _GEN_1085;
                                                          end
                                                        end else begin
                                                          req_signal_r_trans_type <= _GEN_1085;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (!(io_slave_in0_sync)) begin
                                                            req_signal_r_trans_type <= _GEN_1085;
                                                          end
                                                        end else begin
                                                          req_signal_r_trans_type <= _GEN_1085;
                                                        end
                                                      end else begin
                                                        req_signal_r_trans_type <= _GEN_1085;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (!(io_slave_out1_sync)) begin
                                                    if (_T_429) begin
                                                      if (!(io_master_out_sync)) begin
                                                        req_signal_r_trans_type <= _GEN_1139;
                                                      end
                                                    end else begin
                                                      req_signal_r_trans_type <= _GEN_1139;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (!(io_master_out_sync)) begin
                                                      req_signal_r_trans_type <= _GEN_1139;
                                                    end
                                                  end else begin
                                                    req_signal_r_trans_type <= _GEN_1139;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (!(io_slave_out1_sync)) begin
                                                  req_signal_r_trans_type <= _GEN_1171;
                                                end
                                              end else begin
                                                req_signal_r_trans_type <= _GEN_1171;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (!(io_slave_in1_sync)) begin
                                                if (_T_440) begin
                                                  if (!(io_slave_out1_sync)) begin
                                                    req_signal_r_trans_type <= _GEN_1171;
                                                  end
                                                end else begin
                                                  req_signal_r_trans_type <= _GEN_1171;
                                                end
                                              end
                                            end else begin
                                              req_signal_r_trans_type <= _GEN_1203;
                                            end
                                          end else begin
                                            req_signal_r_trans_type <= _GEN_1203;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (!(io_slave_in1_sync)) begin
                                              req_signal_r_trans_type <= _GEN_1203;
                                            end
                                          end else begin
                                            req_signal_r_trans_type <= _GEN_1203;
                                          end
                                        end else begin
                                          req_signal_r_trans_type <= _GEN_1203;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (!(io_slave_in1_sync)) begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (!(io_slave_in1_sync)) begin
                                                req_signal_r_trans_type <= _GEN_1203;
                                              end
                                            end else begin
                                              req_signal_r_trans_type <= _GEN_1203;
                                            end
                                          end else begin
                                            req_signal_r_trans_type <= _GEN_1203;
                                          end
                                        end
                                      end else begin
                                        req_signal_r_trans_type <= _GEN_1257;
                                      end
                                    end else begin
                                      req_signal_r_trans_type <= _GEN_1257;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (!(io_slave_out2_sync)) begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (!(io_slave_in1_sync)) begin
                                          req_signal_r_trans_type <= _GEN_1257;
                                        end
                                      end else begin
                                        req_signal_r_trans_type <= _GEN_1257;
                                      end
                                    end else begin
                                      req_signal_r_trans_type <= _GEN_1257;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (!(io_slave_in1_sync)) begin
                                        req_signal_r_trans_type <= _GEN_1257;
                                      end
                                    end else begin
                                      req_signal_r_trans_type <= _GEN_1257;
                                    end
                                  end else begin
                                    req_signal_r_trans_type <= _GEN_1257;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (!(io_slave_out2_sync)) begin
                                  req_signal_r_trans_type <= _GEN_1311;
                                end
                              end else begin
                                req_signal_r_trans_type <= _GEN_1311;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (!(io_slave_in2_sync)) begin
                                if (_T_479) begin
                                  if (!(io_slave_out2_sync)) begin
                                    req_signal_r_trans_type <= _GEN_1311;
                                  end
                                end else begin
                                  req_signal_r_trans_type <= _GEN_1311;
                                end
                              end
                            end else begin
                              req_signal_r_trans_type <= _GEN_1343;
                            end
                          end else begin
                            req_signal_r_trans_type <= _GEN_1343;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (!(io_slave_in2_sync)) begin
                              req_signal_r_trans_type <= _GEN_1343;
                            end
                          end else begin
                            req_signal_r_trans_type <= _GEN_1343;
                          end
                        end else begin
                          req_signal_r_trans_type <= _GEN_1343;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (!(io_slave_in2_sync)) begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (!(io_slave_in2_sync)) begin
                                req_signal_r_trans_type <= _GEN_1343;
                              end
                            end else begin
                              req_signal_r_trans_type <= _GEN_1343;
                            end
                          end else begin
                            req_signal_r_trans_type <= _GEN_1343;
                          end
                        end
                      end else begin
                        req_signal_r_trans_type <= _GEN_1397;
                      end
                    end else begin
                      req_signal_r_trans_type <= _GEN_1397;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (!(io_slave_out3_sync)) begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (!(io_slave_in2_sync)) begin
                          req_signal_r_trans_type <= _GEN_1397;
                        end
                      end else begin
                        req_signal_r_trans_type <= _GEN_1397;
                      end
                    end else begin
                      req_signal_r_trans_type <= _GEN_1397;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (!(io_slave_in2_sync)) begin
                        req_signal_r_trans_type <= _GEN_1397;
                      end
                    end else begin
                      req_signal_r_trans_type <= _GEN_1397;
                    end
                  end else begin
                    req_signal_r_trans_type <= _GEN_1397;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (!(io_slave_out3_sync)) begin
                  req_signal_r_trans_type <= _GEN_1451;
                end
              end else begin
                req_signal_r_trans_type <= _GEN_1451;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (!(io_slave_in3_sync)) begin
                if (_T_518) begin
                  if (!(io_slave_out3_sync)) begin
                    req_signal_r_trans_type <= _GEN_1451;
                  end
                end else begin
                  req_signal_r_trans_type <= _GEN_1451;
                end
              end
            end else begin
              req_signal_r_trans_type <= _GEN_1483;
            end
          end else begin
            req_signal_r_trans_type <= _GEN_1483;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (!(io_slave_in3_sync)) begin
              req_signal_r_trans_type <= _GEN_1483;
            end
          end else begin
            req_signal_r_trans_type <= _GEN_1483;
          end
        end else begin
          req_signal_r_trans_type <= _GEN_1483;
        end
      end
    end
    if (reset) begin
      resp_signal_r_ack <= 32'h2;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            resp_signal_r_ack <= io_slave_in3_ack;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  resp_signal_r_ack <= io_slave_in3_ack;
                end else begin
                  if (_T_518) begin
                    if (!(io_slave_out3_sync)) begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            resp_signal_r_ack <= io_slave_in2_ack;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  resp_signal_r_ack <= io_slave_in2_ack;
                                end else begin
                                  if (_T_479) begin
                                    if (!(io_slave_out2_sync)) begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            resp_signal_r_ack <= io_slave_in1_ack;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  resp_signal_r_ack <= io_slave_in1_ack;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (!(io_slave_out1_sync)) begin
                                                      if (_T_429) begin
                                                        if (!(io_master_out_sync)) begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                resp_signal_r_ack <= io_slave_in0_ack;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      resp_signal_r_ack <= io_slave_in0_ack;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (!(io_slave_out0_sync)) begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (!(io_master_in_sync)) begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (!(io_master_in_sync)) begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (!(io_master_in_sync)) begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (!(io_master_in_sync)) begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (!(io_master_in_sync)) begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (!(io_master_in_sync)) begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    resp_signal_r_ack <= 32'h0;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  resp_signal_r_ack <= 32'h0;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                resp_signal_r_ack <= 32'h0;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              resp_signal_r_ack <= 32'h0;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            resp_signal_r_ack <= 32'h0;
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            resp_signal_r_ack <= _GEN_304;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          resp_signal_r_ack <= _GEN_304;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        resp_signal_r_ack <= _GEN_304;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  resp_signal_r_ack <= 32'h0;
                                                                                                                                                end else begin
                                                                                                                                                  resp_signal_r_ack <= _GEN_304;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                resp_signal_r_ack <= _GEN_304;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              resp_signal_r_ack <= _GEN_304;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            resp_signal_r_ack <= _GEN_304;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          resp_signal_r_ack <= _GEN_304;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        resp_signal_r_ack <= _GEN_304;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      resp_signal_r_ack <= _GEN_304;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                resp_signal_r_ack <= 32'h0;
                                                                                                                                              end else begin
                                                                                                                                                resp_signal_r_ack <= _GEN_304;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              resp_signal_r_ack <= _GEN_304;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            resp_signal_r_ack <= _GEN_304;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          resp_signal_r_ack <= _GEN_304;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        resp_signal_r_ack <= _GEN_304;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      resp_signal_r_ack <= _GEN_304;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    resp_signal_r_ack <= _GEN_304;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              resp_signal_r_ack <= 32'h0;
                                                                                                                                            end else begin
                                                                                                                                              resp_signal_r_ack <= _GEN_304;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            resp_signal_r_ack <= _GEN_304;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          resp_signal_r_ack <= _GEN_304;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        resp_signal_r_ack <= _GEN_304;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      resp_signal_r_ack <= _GEN_304;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    resp_signal_r_ack <= _GEN_304;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  resp_signal_r_ack <= _GEN_304;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              resp_signal_r_ack <= _GEN_430;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (!(io_master_in_sync)) begin
                                                                                                                                    resp_signal_r_ack <= _GEN_430;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  resp_signal_r_ack <= _GEN_430;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                resp_signal_r_ack <= _GEN_430;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              resp_signal_r_ack <= _GEN_430;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            resp_signal_r_ack <= _GEN_430;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (!(io_master_in_sync)) begin
                                                                                                                                  resp_signal_r_ack <= _GEN_430;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                resp_signal_r_ack <= _GEN_430;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              resp_signal_r_ack <= _GEN_430;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            resp_signal_r_ack <= _GEN_430;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          resp_signal_r_ack <= _GEN_430;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (!(io_master_in_sync)) begin
                                                                                                                                resp_signal_r_ack <= _GEN_430;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              resp_signal_r_ack <= _GEN_430;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            resp_signal_r_ack <= _GEN_430;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          resp_signal_r_ack <= _GEN_430;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        resp_signal_r_ack <= _GEN_430;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    resp_signal_r_ack <= _GEN_522;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (!(io_master_in_sync)) begin
                                                                                                                          resp_signal_r_ack <= _GEN_522;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        resp_signal_r_ack <= _GEN_522;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      resp_signal_r_ack <= _GEN_522;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    resp_signal_r_ack <= _GEN_522;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  resp_signal_r_ack <= _GEN_522;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (!(io_master_in_sync)) begin
                                                                                                                        resp_signal_r_ack <= _GEN_522;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      resp_signal_r_ack <= _GEN_522;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    resp_signal_r_ack <= _GEN_522;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  resp_signal_r_ack <= _GEN_522;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                resp_signal_r_ack <= _GEN_522;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (!(io_master_in_sync)) begin
                                                                                                                      resp_signal_r_ack <= _GEN_522;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    resp_signal_r_ack <= _GEN_522;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  resp_signal_r_ack <= _GEN_522;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                resp_signal_r_ack <= _GEN_522;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              resp_signal_r_ack <= _GEN_522;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          resp_signal_r_ack <= _GEN_617;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (!(io_master_in_sync)) begin
                                                                                                                resp_signal_r_ack <= _GEN_617;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              resp_signal_r_ack <= _GEN_617;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            resp_signal_r_ack <= _GEN_617;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          resp_signal_r_ack <= _GEN_617;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        resp_signal_r_ack <= _GEN_617;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (!(io_master_in_sync)) begin
                                                                                                              resp_signal_r_ack <= _GEN_617;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            resp_signal_r_ack <= _GEN_617;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          resp_signal_r_ack <= _GEN_617;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        resp_signal_r_ack <= _GEN_617;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      resp_signal_r_ack <= _GEN_617;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (!(io_master_in_sync)) begin
                                                                                                            resp_signal_r_ack <= _GEN_617;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          resp_signal_r_ack <= _GEN_617;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        resp_signal_r_ack <= _GEN_617;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      resp_signal_r_ack <= _GEN_617;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    resp_signal_r_ack <= _GEN_617;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                resp_signal_r_ack <= _GEN_712;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (!(io_master_in_sync)) begin
                                                                                                      resp_signal_r_ack <= _GEN_712;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    resp_signal_r_ack <= _GEN_712;
                                                                                                  end
                                                                                                end else begin
                                                                                                  resp_signal_r_ack <= _GEN_712;
                                                                                                end
                                                                                              end else begin
                                                                                                resp_signal_r_ack <= _GEN_712;
                                                                                              end
                                                                                            end else begin
                                                                                              resp_signal_r_ack <= _GEN_712;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (!(io_master_in_sync)) begin
                                                                                                    resp_signal_r_ack <= _GEN_712;
                                                                                                  end
                                                                                                end else begin
                                                                                                  resp_signal_r_ack <= _GEN_712;
                                                                                                end
                                                                                              end else begin
                                                                                                resp_signal_r_ack <= _GEN_712;
                                                                                              end
                                                                                            end else begin
                                                                                              resp_signal_r_ack <= _GEN_712;
                                                                                            end
                                                                                          end else begin
                                                                                            resp_signal_r_ack <= _GEN_712;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (!(io_master_in_sync)) begin
                                                                                                  resp_signal_r_ack <= _GEN_712;
                                                                                                end
                                                                                              end else begin
                                                                                                resp_signal_r_ack <= _GEN_712;
                                                                                              end
                                                                                            end else begin
                                                                                              resp_signal_r_ack <= _GEN_712;
                                                                                            end
                                                                                          end else begin
                                                                                            resp_signal_r_ack <= _GEN_712;
                                                                                          end
                                                                                        end else begin
                                                                                          resp_signal_r_ack <= _GEN_712;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      resp_signal_r_ack <= _GEN_807;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (!(io_master_in_sync)) begin
                                                                                            resp_signal_r_ack <= _GEN_807;
                                                                                          end
                                                                                        end else begin
                                                                                          resp_signal_r_ack <= _GEN_807;
                                                                                        end
                                                                                      end else begin
                                                                                        resp_signal_r_ack <= _GEN_807;
                                                                                      end
                                                                                    end else begin
                                                                                      resp_signal_r_ack <= _GEN_807;
                                                                                    end
                                                                                  end else begin
                                                                                    resp_signal_r_ack <= _GEN_807;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (!(io_master_in_sync)) begin
                                                                                          resp_signal_r_ack <= _GEN_807;
                                                                                        end
                                                                                      end else begin
                                                                                        resp_signal_r_ack <= _GEN_807;
                                                                                      end
                                                                                    end else begin
                                                                                      resp_signal_r_ack <= _GEN_807;
                                                                                    end
                                                                                  end else begin
                                                                                    resp_signal_r_ack <= _GEN_807;
                                                                                  end
                                                                                end else begin
                                                                                  resp_signal_r_ack <= _GEN_807;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (!(io_master_in_sync)) begin
                                                                                        resp_signal_r_ack <= _GEN_807;
                                                                                      end
                                                                                    end else begin
                                                                                      resp_signal_r_ack <= _GEN_807;
                                                                                    end
                                                                                  end else begin
                                                                                    resp_signal_r_ack <= _GEN_807;
                                                                                  end
                                                                                end else begin
                                                                                  resp_signal_r_ack <= _GEN_807;
                                                                                end
                                                                              end else begin
                                                                                resp_signal_r_ack <= _GEN_807;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            resp_signal_r_ack <= _GEN_902;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (!(io_master_in_sync)) begin
                                                                                  resp_signal_r_ack <= _GEN_902;
                                                                                end
                                                                              end else begin
                                                                                resp_signal_r_ack <= _GEN_902;
                                                                              end
                                                                            end else begin
                                                                              resp_signal_r_ack <= _GEN_902;
                                                                            end
                                                                          end else begin
                                                                            resp_signal_r_ack <= _GEN_902;
                                                                          end
                                                                        end else begin
                                                                          resp_signal_r_ack <= _GEN_902;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (!(io_slave_out0_sync)) begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (!(io_master_in_sync)) begin
                                                                                  resp_signal_r_ack <= _GEN_902;
                                                                                end
                                                                              end else begin
                                                                                resp_signal_r_ack <= _GEN_902;
                                                                              end
                                                                            end else begin
                                                                              resp_signal_r_ack <= _GEN_902;
                                                                            end
                                                                          end else begin
                                                                            resp_signal_r_ack <= _GEN_902;
                                                                          end
                                                                        end else begin
                                                                          resp_signal_r_ack <= _GEN_902;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (!(io_master_in_sync)) begin
                                                                                resp_signal_r_ack <= _GEN_902;
                                                                              end
                                                                            end else begin
                                                                              resp_signal_r_ack <= _GEN_902;
                                                                            end
                                                                          end else begin
                                                                            resp_signal_r_ack <= _GEN_902;
                                                                          end
                                                                        end else begin
                                                                          resp_signal_r_ack <= _GEN_902;
                                                                        end
                                                                      end else begin
                                                                        resp_signal_r_ack <= _GEN_902;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (!(io_slave_out0_sync)) begin
                                                                      resp_signal_r_ack <= _GEN_997;
                                                                    end
                                                                  end else begin
                                                                    resp_signal_r_ack <= _GEN_997;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    resp_signal_r_ack <= io_slave_in0_ack;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (!(io_slave_out0_sync)) begin
                                                                        resp_signal_r_ack <= _GEN_997;
                                                                      end
                                                                    end else begin
                                                                      resp_signal_r_ack <= _GEN_997;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  resp_signal_r_ack <= _GEN_1032;
                                                                end
                                                              end else begin
                                                                resp_signal_r_ack <= _GEN_1032;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  resp_signal_r_ack <= io_slave_in0_ack;
                                                                end else begin
                                                                  resp_signal_r_ack <= _GEN_1032;
                                                                end
                                                              end else begin
                                                                resp_signal_r_ack <= _GEN_1032;
                                                              end
                                                            end else begin
                                                              resp_signal_r_ack <= _GEN_1032;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              resp_signal_r_ack <= io_slave_in0_ack;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    resp_signal_r_ack <= io_slave_in0_ack;
                                                                  end else begin
                                                                    resp_signal_r_ack <= _GEN_1032;
                                                                  end
                                                                end else begin
                                                                  resp_signal_r_ack <= _GEN_1032;
                                                                end
                                                              end else begin
                                                                resp_signal_r_ack <= _GEN_1032;
                                                              end
                                                            end
                                                          end else begin
                                                            resp_signal_r_ack <= _GEN_1086;
                                                          end
                                                        end else begin
                                                          resp_signal_r_ack <= _GEN_1086;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (!(io_master_out_sync)) begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              resp_signal_r_ack <= io_slave_in0_ack;
                                                            end else begin
                                                              resp_signal_r_ack <= _GEN_1086;
                                                            end
                                                          end else begin
                                                            resp_signal_r_ack <= _GEN_1086;
                                                          end
                                                        end else begin
                                                          resp_signal_r_ack <= _GEN_1086;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            resp_signal_r_ack <= io_slave_in0_ack;
                                                          end else begin
                                                            resp_signal_r_ack <= _GEN_1086;
                                                          end
                                                        end else begin
                                                          resp_signal_r_ack <= _GEN_1086;
                                                        end
                                                      end else begin
                                                        resp_signal_r_ack <= _GEN_1086;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (!(io_slave_out1_sync)) begin
                                                    if (_T_429) begin
                                                      if (!(io_master_out_sync)) begin
                                                        resp_signal_r_ack <= _GEN_1140;
                                                      end
                                                    end else begin
                                                      resp_signal_r_ack <= _GEN_1140;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (!(io_master_out_sync)) begin
                                                      resp_signal_r_ack <= _GEN_1140;
                                                    end
                                                  end else begin
                                                    resp_signal_r_ack <= _GEN_1140;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (!(io_slave_out1_sync)) begin
                                                  resp_signal_r_ack <= _GEN_1172;
                                                end
                                              end else begin
                                                resp_signal_r_ack <= _GEN_1172;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                resp_signal_r_ack <= io_slave_in1_ack;
                                              end else begin
                                                if (_T_440) begin
                                                  if (!(io_slave_out1_sync)) begin
                                                    resp_signal_r_ack <= _GEN_1172;
                                                  end
                                                end else begin
                                                  resp_signal_r_ack <= _GEN_1172;
                                                end
                                              end
                                            end else begin
                                              resp_signal_r_ack <= _GEN_1204;
                                            end
                                          end else begin
                                            resp_signal_r_ack <= _GEN_1204;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              resp_signal_r_ack <= io_slave_in1_ack;
                                            end else begin
                                              resp_signal_r_ack <= _GEN_1204;
                                            end
                                          end else begin
                                            resp_signal_r_ack <= _GEN_1204;
                                          end
                                        end else begin
                                          resp_signal_r_ack <= _GEN_1204;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          resp_signal_r_ack <= io_slave_in1_ack;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                resp_signal_r_ack <= io_slave_in1_ack;
                                              end else begin
                                                resp_signal_r_ack <= _GEN_1204;
                                              end
                                            end else begin
                                              resp_signal_r_ack <= _GEN_1204;
                                            end
                                          end else begin
                                            resp_signal_r_ack <= _GEN_1204;
                                          end
                                        end
                                      end else begin
                                        resp_signal_r_ack <= _GEN_1258;
                                      end
                                    end else begin
                                      resp_signal_r_ack <= _GEN_1258;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (!(io_slave_out2_sync)) begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          resp_signal_r_ack <= io_slave_in1_ack;
                                        end else begin
                                          resp_signal_r_ack <= _GEN_1258;
                                        end
                                      end else begin
                                        resp_signal_r_ack <= _GEN_1258;
                                      end
                                    end else begin
                                      resp_signal_r_ack <= _GEN_1258;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        resp_signal_r_ack <= io_slave_in1_ack;
                                      end else begin
                                        resp_signal_r_ack <= _GEN_1258;
                                      end
                                    end else begin
                                      resp_signal_r_ack <= _GEN_1258;
                                    end
                                  end else begin
                                    resp_signal_r_ack <= _GEN_1258;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (!(io_slave_out2_sync)) begin
                                  resp_signal_r_ack <= _GEN_1312;
                                end
                              end else begin
                                resp_signal_r_ack <= _GEN_1312;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                resp_signal_r_ack <= io_slave_in2_ack;
                              end else begin
                                if (_T_479) begin
                                  if (!(io_slave_out2_sync)) begin
                                    resp_signal_r_ack <= _GEN_1312;
                                  end
                                end else begin
                                  resp_signal_r_ack <= _GEN_1312;
                                end
                              end
                            end else begin
                              resp_signal_r_ack <= _GEN_1344;
                            end
                          end else begin
                            resp_signal_r_ack <= _GEN_1344;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              resp_signal_r_ack <= io_slave_in2_ack;
                            end else begin
                              resp_signal_r_ack <= _GEN_1344;
                            end
                          end else begin
                            resp_signal_r_ack <= _GEN_1344;
                          end
                        end else begin
                          resp_signal_r_ack <= _GEN_1344;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          resp_signal_r_ack <= io_slave_in2_ack;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                resp_signal_r_ack <= io_slave_in2_ack;
                              end else begin
                                resp_signal_r_ack <= _GEN_1344;
                              end
                            end else begin
                              resp_signal_r_ack <= _GEN_1344;
                            end
                          end else begin
                            resp_signal_r_ack <= _GEN_1344;
                          end
                        end
                      end else begin
                        resp_signal_r_ack <= _GEN_1398;
                      end
                    end else begin
                      resp_signal_r_ack <= _GEN_1398;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (!(io_slave_out3_sync)) begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          resp_signal_r_ack <= io_slave_in2_ack;
                        end else begin
                          resp_signal_r_ack <= _GEN_1398;
                        end
                      end else begin
                        resp_signal_r_ack <= _GEN_1398;
                      end
                    end else begin
                      resp_signal_r_ack <= _GEN_1398;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        resp_signal_r_ack <= io_slave_in2_ack;
                      end else begin
                        resp_signal_r_ack <= _GEN_1398;
                      end
                    end else begin
                      resp_signal_r_ack <= _GEN_1398;
                    end
                  end else begin
                    resp_signal_r_ack <= _GEN_1398;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (!(io_slave_out3_sync)) begin
                  resp_signal_r_ack <= _GEN_1452;
                end
              end else begin
                resp_signal_r_ack <= _GEN_1452;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                resp_signal_r_ack <= io_slave_in3_ack;
              end else begin
                if (_T_518) begin
                  if (!(io_slave_out3_sync)) begin
                    resp_signal_r_ack <= _GEN_1452;
                  end
                end else begin
                  resp_signal_r_ack <= _GEN_1452;
                end
              end
            end else begin
              resp_signal_r_ack <= _GEN_1484;
            end
          end else begin
            resp_signal_r_ack <= _GEN_1484;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              resp_signal_r_ack <= io_slave_in3_ack;
            end else begin
              resp_signal_r_ack <= _GEN_1484;
            end
          end else begin
            resp_signal_r_ack <= _GEN_1484;
          end
        end else begin
          resp_signal_r_ack <= _GEN_1484;
        end
      end
    end
    if (reset) begin
      resp_signal_r_data <= 32'sh0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            resp_signal_r_data <= 32'sh0;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  resp_signal_r_data <= io_slave_in3_data;
                end else begin
                  if (_T_518) begin
                    if (!(io_slave_out3_sync)) begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            resp_signal_r_data <= 32'sh0;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  resp_signal_r_data <= io_slave_in2_data;
                                end else begin
                                  if (_T_479) begin
                                    if (!(io_slave_out2_sync)) begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            resp_signal_r_data <= 32'sh0;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  resp_signal_r_data <= io_slave_in1_data;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (!(io_slave_out1_sync)) begin
                                                      if (_T_429) begin
                                                        if (!(io_master_out_sync)) begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                resp_signal_r_data <= 32'sh0;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      resp_signal_r_data <= io_slave_in0_data;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (!(io_slave_out0_sync)) begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (!(io_master_in_sync)) begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (!(io_master_in_sync)) begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (!(io_master_in_sync)) begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (!(io_master_in_sync)) begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (!(io_master_in_sync)) begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (!(io_master_in_sync)) begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    resp_signal_r_data <= 32'sh0;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  resp_signal_r_data <= 32'sh0;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                resp_signal_r_data <= 32'sh0;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              resp_signal_r_data <= 32'sh0;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            resp_signal_r_data <= 32'sh0;
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            resp_signal_r_data <= _GEN_305;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          resp_signal_r_data <= _GEN_305;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        resp_signal_r_data <= _GEN_305;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  resp_signal_r_data <= 32'sh0;
                                                                                                                                                end else begin
                                                                                                                                                  resp_signal_r_data <= _GEN_305;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                resp_signal_r_data <= _GEN_305;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              resp_signal_r_data <= _GEN_305;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            resp_signal_r_data <= _GEN_305;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          resp_signal_r_data <= _GEN_305;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        resp_signal_r_data <= _GEN_305;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      resp_signal_r_data <= _GEN_305;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                resp_signal_r_data <= 32'sh0;
                                                                                                                                              end else begin
                                                                                                                                                resp_signal_r_data <= _GEN_305;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              resp_signal_r_data <= _GEN_305;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            resp_signal_r_data <= _GEN_305;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          resp_signal_r_data <= _GEN_305;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        resp_signal_r_data <= _GEN_305;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      resp_signal_r_data <= _GEN_305;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    resp_signal_r_data <= _GEN_305;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              resp_signal_r_data <= 32'sh0;
                                                                                                                                            end else begin
                                                                                                                                              resp_signal_r_data <= _GEN_305;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            resp_signal_r_data <= _GEN_305;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          resp_signal_r_data <= _GEN_305;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        resp_signal_r_data <= _GEN_305;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      resp_signal_r_data <= _GEN_305;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    resp_signal_r_data <= _GEN_305;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  resp_signal_r_data <= _GEN_305;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              resp_signal_r_data <= _GEN_431;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (!(io_master_in_sync)) begin
                                                                                                                                    resp_signal_r_data <= _GEN_431;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  resp_signal_r_data <= _GEN_431;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                resp_signal_r_data <= _GEN_431;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              resp_signal_r_data <= _GEN_431;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            resp_signal_r_data <= _GEN_431;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (!(io_master_in_sync)) begin
                                                                                                                                  resp_signal_r_data <= _GEN_431;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                resp_signal_r_data <= _GEN_431;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              resp_signal_r_data <= _GEN_431;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            resp_signal_r_data <= _GEN_431;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          resp_signal_r_data <= _GEN_431;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (!(io_master_in_sync)) begin
                                                                                                                                resp_signal_r_data <= _GEN_431;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              resp_signal_r_data <= _GEN_431;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            resp_signal_r_data <= _GEN_431;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          resp_signal_r_data <= _GEN_431;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        resp_signal_r_data <= _GEN_431;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    resp_signal_r_data <= _GEN_523;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (!(io_master_in_sync)) begin
                                                                                                                          resp_signal_r_data <= _GEN_523;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        resp_signal_r_data <= _GEN_523;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      resp_signal_r_data <= _GEN_523;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    resp_signal_r_data <= _GEN_523;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  resp_signal_r_data <= _GEN_523;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (!(io_master_in_sync)) begin
                                                                                                                        resp_signal_r_data <= _GEN_523;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      resp_signal_r_data <= _GEN_523;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    resp_signal_r_data <= _GEN_523;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  resp_signal_r_data <= _GEN_523;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                resp_signal_r_data <= _GEN_523;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (!(io_master_in_sync)) begin
                                                                                                                      resp_signal_r_data <= _GEN_523;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    resp_signal_r_data <= _GEN_523;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  resp_signal_r_data <= _GEN_523;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                resp_signal_r_data <= _GEN_523;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              resp_signal_r_data <= _GEN_523;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          resp_signal_r_data <= _GEN_618;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (!(io_master_in_sync)) begin
                                                                                                                resp_signal_r_data <= _GEN_618;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              resp_signal_r_data <= _GEN_618;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            resp_signal_r_data <= _GEN_618;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          resp_signal_r_data <= _GEN_618;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        resp_signal_r_data <= _GEN_618;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (!(io_master_in_sync)) begin
                                                                                                              resp_signal_r_data <= _GEN_618;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            resp_signal_r_data <= _GEN_618;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          resp_signal_r_data <= _GEN_618;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        resp_signal_r_data <= _GEN_618;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      resp_signal_r_data <= _GEN_618;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (!(io_master_in_sync)) begin
                                                                                                            resp_signal_r_data <= _GEN_618;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          resp_signal_r_data <= _GEN_618;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        resp_signal_r_data <= _GEN_618;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      resp_signal_r_data <= _GEN_618;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    resp_signal_r_data <= _GEN_618;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                resp_signal_r_data <= _GEN_713;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (!(io_master_in_sync)) begin
                                                                                                      resp_signal_r_data <= _GEN_713;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    resp_signal_r_data <= _GEN_713;
                                                                                                  end
                                                                                                end else begin
                                                                                                  resp_signal_r_data <= _GEN_713;
                                                                                                end
                                                                                              end else begin
                                                                                                resp_signal_r_data <= _GEN_713;
                                                                                              end
                                                                                            end else begin
                                                                                              resp_signal_r_data <= _GEN_713;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (!(io_master_in_sync)) begin
                                                                                                    resp_signal_r_data <= _GEN_713;
                                                                                                  end
                                                                                                end else begin
                                                                                                  resp_signal_r_data <= _GEN_713;
                                                                                                end
                                                                                              end else begin
                                                                                                resp_signal_r_data <= _GEN_713;
                                                                                              end
                                                                                            end else begin
                                                                                              resp_signal_r_data <= _GEN_713;
                                                                                            end
                                                                                          end else begin
                                                                                            resp_signal_r_data <= _GEN_713;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (!(io_master_in_sync)) begin
                                                                                                  resp_signal_r_data <= _GEN_713;
                                                                                                end
                                                                                              end else begin
                                                                                                resp_signal_r_data <= _GEN_713;
                                                                                              end
                                                                                            end else begin
                                                                                              resp_signal_r_data <= _GEN_713;
                                                                                            end
                                                                                          end else begin
                                                                                            resp_signal_r_data <= _GEN_713;
                                                                                          end
                                                                                        end else begin
                                                                                          resp_signal_r_data <= _GEN_713;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      resp_signal_r_data <= _GEN_808;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (!(io_master_in_sync)) begin
                                                                                            resp_signal_r_data <= _GEN_808;
                                                                                          end
                                                                                        end else begin
                                                                                          resp_signal_r_data <= _GEN_808;
                                                                                        end
                                                                                      end else begin
                                                                                        resp_signal_r_data <= _GEN_808;
                                                                                      end
                                                                                    end else begin
                                                                                      resp_signal_r_data <= _GEN_808;
                                                                                    end
                                                                                  end else begin
                                                                                    resp_signal_r_data <= _GEN_808;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (!(io_master_in_sync)) begin
                                                                                          resp_signal_r_data <= _GEN_808;
                                                                                        end
                                                                                      end else begin
                                                                                        resp_signal_r_data <= _GEN_808;
                                                                                      end
                                                                                    end else begin
                                                                                      resp_signal_r_data <= _GEN_808;
                                                                                    end
                                                                                  end else begin
                                                                                    resp_signal_r_data <= _GEN_808;
                                                                                  end
                                                                                end else begin
                                                                                  resp_signal_r_data <= _GEN_808;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (!(io_master_in_sync)) begin
                                                                                        resp_signal_r_data <= _GEN_808;
                                                                                      end
                                                                                    end else begin
                                                                                      resp_signal_r_data <= _GEN_808;
                                                                                    end
                                                                                  end else begin
                                                                                    resp_signal_r_data <= _GEN_808;
                                                                                  end
                                                                                end else begin
                                                                                  resp_signal_r_data <= _GEN_808;
                                                                                end
                                                                              end else begin
                                                                                resp_signal_r_data <= _GEN_808;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            resp_signal_r_data <= _GEN_903;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (!(io_master_in_sync)) begin
                                                                                  resp_signal_r_data <= _GEN_903;
                                                                                end
                                                                              end else begin
                                                                                resp_signal_r_data <= _GEN_903;
                                                                              end
                                                                            end else begin
                                                                              resp_signal_r_data <= _GEN_903;
                                                                            end
                                                                          end else begin
                                                                            resp_signal_r_data <= _GEN_903;
                                                                          end
                                                                        end else begin
                                                                          resp_signal_r_data <= _GEN_903;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (!(io_slave_out0_sync)) begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (!(io_master_in_sync)) begin
                                                                                  resp_signal_r_data <= _GEN_903;
                                                                                end
                                                                              end else begin
                                                                                resp_signal_r_data <= _GEN_903;
                                                                              end
                                                                            end else begin
                                                                              resp_signal_r_data <= _GEN_903;
                                                                            end
                                                                          end else begin
                                                                            resp_signal_r_data <= _GEN_903;
                                                                          end
                                                                        end else begin
                                                                          resp_signal_r_data <= _GEN_903;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (!(io_master_in_sync)) begin
                                                                                resp_signal_r_data <= _GEN_903;
                                                                              end
                                                                            end else begin
                                                                              resp_signal_r_data <= _GEN_903;
                                                                            end
                                                                          end else begin
                                                                            resp_signal_r_data <= _GEN_903;
                                                                          end
                                                                        end else begin
                                                                          resp_signal_r_data <= _GEN_903;
                                                                        end
                                                                      end else begin
                                                                        resp_signal_r_data <= _GEN_903;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (!(io_slave_out0_sync)) begin
                                                                      resp_signal_r_data <= _GEN_998;
                                                                    end
                                                                  end else begin
                                                                    resp_signal_r_data <= _GEN_998;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    resp_signal_r_data <= io_slave_in0_data;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (!(io_slave_out0_sync)) begin
                                                                        resp_signal_r_data <= _GEN_998;
                                                                      end
                                                                    end else begin
                                                                      resp_signal_r_data <= _GEN_998;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  resp_signal_r_data <= _GEN_1033;
                                                                end
                                                              end else begin
                                                                resp_signal_r_data <= _GEN_1033;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  resp_signal_r_data <= io_slave_in0_data;
                                                                end else begin
                                                                  resp_signal_r_data <= _GEN_1033;
                                                                end
                                                              end else begin
                                                                resp_signal_r_data <= _GEN_1033;
                                                              end
                                                            end else begin
                                                              resp_signal_r_data <= _GEN_1033;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              resp_signal_r_data <= 32'sh0;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    resp_signal_r_data <= io_slave_in0_data;
                                                                  end else begin
                                                                    resp_signal_r_data <= _GEN_1033;
                                                                  end
                                                                end else begin
                                                                  resp_signal_r_data <= _GEN_1033;
                                                                end
                                                              end else begin
                                                                resp_signal_r_data <= _GEN_1033;
                                                              end
                                                            end
                                                          end else begin
                                                            resp_signal_r_data <= _GEN_1087;
                                                          end
                                                        end else begin
                                                          resp_signal_r_data <= _GEN_1087;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (!(io_master_out_sync)) begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              resp_signal_r_data <= 32'sh0;
                                                            end else begin
                                                              resp_signal_r_data <= _GEN_1087;
                                                            end
                                                          end else begin
                                                            resp_signal_r_data <= _GEN_1087;
                                                          end
                                                        end else begin
                                                          resp_signal_r_data <= _GEN_1087;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            resp_signal_r_data <= 32'sh0;
                                                          end else begin
                                                            resp_signal_r_data <= _GEN_1087;
                                                          end
                                                        end else begin
                                                          resp_signal_r_data <= _GEN_1087;
                                                        end
                                                      end else begin
                                                        resp_signal_r_data <= _GEN_1087;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (!(io_slave_out1_sync)) begin
                                                    if (_T_429) begin
                                                      if (!(io_master_out_sync)) begin
                                                        resp_signal_r_data <= _GEN_1141;
                                                      end
                                                    end else begin
                                                      resp_signal_r_data <= _GEN_1141;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (!(io_master_out_sync)) begin
                                                      resp_signal_r_data <= _GEN_1141;
                                                    end
                                                  end else begin
                                                    resp_signal_r_data <= _GEN_1141;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (!(io_slave_out1_sync)) begin
                                                  resp_signal_r_data <= _GEN_1173;
                                                end
                                              end else begin
                                                resp_signal_r_data <= _GEN_1173;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                resp_signal_r_data <= io_slave_in1_data;
                                              end else begin
                                                if (_T_440) begin
                                                  if (!(io_slave_out1_sync)) begin
                                                    resp_signal_r_data <= _GEN_1173;
                                                  end
                                                end else begin
                                                  resp_signal_r_data <= _GEN_1173;
                                                end
                                              end
                                            end else begin
                                              resp_signal_r_data <= _GEN_1205;
                                            end
                                          end else begin
                                            resp_signal_r_data <= _GEN_1205;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              resp_signal_r_data <= io_slave_in1_data;
                                            end else begin
                                              resp_signal_r_data <= _GEN_1205;
                                            end
                                          end else begin
                                            resp_signal_r_data <= _GEN_1205;
                                          end
                                        end else begin
                                          resp_signal_r_data <= _GEN_1205;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          resp_signal_r_data <= 32'sh0;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                resp_signal_r_data <= io_slave_in1_data;
                                              end else begin
                                                resp_signal_r_data <= _GEN_1205;
                                              end
                                            end else begin
                                              resp_signal_r_data <= _GEN_1205;
                                            end
                                          end else begin
                                            resp_signal_r_data <= _GEN_1205;
                                          end
                                        end
                                      end else begin
                                        resp_signal_r_data <= _GEN_1259;
                                      end
                                    end else begin
                                      resp_signal_r_data <= _GEN_1259;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (!(io_slave_out2_sync)) begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          resp_signal_r_data <= 32'sh0;
                                        end else begin
                                          resp_signal_r_data <= _GEN_1259;
                                        end
                                      end else begin
                                        resp_signal_r_data <= _GEN_1259;
                                      end
                                    end else begin
                                      resp_signal_r_data <= _GEN_1259;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        resp_signal_r_data <= 32'sh0;
                                      end else begin
                                        resp_signal_r_data <= _GEN_1259;
                                      end
                                    end else begin
                                      resp_signal_r_data <= _GEN_1259;
                                    end
                                  end else begin
                                    resp_signal_r_data <= _GEN_1259;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (!(io_slave_out2_sync)) begin
                                  resp_signal_r_data <= _GEN_1313;
                                end
                              end else begin
                                resp_signal_r_data <= _GEN_1313;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                resp_signal_r_data <= io_slave_in2_data;
                              end else begin
                                if (_T_479) begin
                                  if (!(io_slave_out2_sync)) begin
                                    resp_signal_r_data <= _GEN_1313;
                                  end
                                end else begin
                                  resp_signal_r_data <= _GEN_1313;
                                end
                              end
                            end else begin
                              resp_signal_r_data <= _GEN_1345;
                            end
                          end else begin
                            resp_signal_r_data <= _GEN_1345;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              resp_signal_r_data <= io_slave_in2_data;
                            end else begin
                              resp_signal_r_data <= _GEN_1345;
                            end
                          end else begin
                            resp_signal_r_data <= _GEN_1345;
                          end
                        end else begin
                          resp_signal_r_data <= _GEN_1345;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          resp_signal_r_data <= 32'sh0;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                resp_signal_r_data <= io_slave_in2_data;
                              end else begin
                                resp_signal_r_data <= _GEN_1345;
                              end
                            end else begin
                              resp_signal_r_data <= _GEN_1345;
                            end
                          end else begin
                            resp_signal_r_data <= _GEN_1345;
                          end
                        end
                      end else begin
                        resp_signal_r_data <= _GEN_1399;
                      end
                    end else begin
                      resp_signal_r_data <= _GEN_1399;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (!(io_slave_out3_sync)) begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          resp_signal_r_data <= 32'sh0;
                        end else begin
                          resp_signal_r_data <= _GEN_1399;
                        end
                      end else begin
                        resp_signal_r_data <= _GEN_1399;
                      end
                    end else begin
                      resp_signal_r_data <= _GEN_1399;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        resp_signal_r_data <= 32'sh0;
                      end else begin
                        resp_signal_r_data <= _GEN_1399;
                      end
                    end else begin
                      resp_signal_r_data <= _GEN_1399;
                    end
                  end else begin
                    resp_signal_r_data <= _GEN_1399;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (!(io_slave_out3_sync)) begin
                  resp_signal_r_data <= _GEN_1453;
                end
              end else begin
                resp_signal_r_data <= _GEN_1453;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                resp_signal_r_data <= io_slave_in3_data;
              end else begin
                if (_T_518) begin
                  if (!(io_slave_out3_sync)) begin
                    resp_signal_r_data <= _GEN_1453;
                  end
                end else begin
                  resp_signal_r_data <= _GEN_1453;
                end
              end
            end else begin
              resp_signal_r_data <= _GEN_1485;
            end
          end else begin
            resp_signal_r_data <= _GEN_1485;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              resp_signal_r_data <= io_slave_in3_data;
            end else begin
              resp_signal_r_data <= _GEN_1485;
            end
          end else begin
            resp_signal_r_data <= _GEN_1485;
          end
        end else begin
          resp_signal_r_data <= _GEN_1485;
        end
      end
    end
    if (reset) begin
      state_r <= 4'h0;
    end else begin
      if (_T_529) begin
        if (_T_402) begin
          if (io_slave_in3_sync) begin
            state_r <= 4'h3;
          end else begin
            if (_T_529) begin
              if (_T_404) begin
                if (io_slave_in3_sync) begin
                  state_r <= 4'h3;
                end else begin
                  if (_T_518) begin
                    if (io_slave_out3_sync) begin
                      state_r <= 4'h9;
                    end else begin
                      if (_T_490) begin
                        if (_T_402) begin
                          if (io_slave_in2_sync) begin
                            state_r <= 4'h3;
                          end else begin
                            if (_T_490) begin
                              if (_T_404) begin
                                if (io_slave_in2_sync) begin
                                  state_r <= 4'h3;
                                end else begin
                                  if (_T_479) begin
                                    if (io_slave_out2_sync) begin
                                      state_r <= 4'h7;
                                    end else begin
                                      if (_T_451) begin
                                        if (_T_402) begin
                                          if (io_slave_in1_sync) begin
                                            state_r <= 4'h3;
                                          end else begin
                                            if (_T_451) begin
                                              if (_T_404) begin
                                                if (io_slave_in1_sync) begin
                                                  state_r <= 4'h3;
                                                end else begin
                                                  if (_T_440) begin
                                                    if (io_slave_out1_sync) begin
                                                      state_r <= 4'h5;
                                                    end else begin
                                                      if (_T_429) begin
                                                        if (io_master_out_sync) begin
                                                          state_r <= 4'h0;
                                                        end else begin
                                                          if (_T_401) begin
                                                            if (_T_402) begin
                                                              if (io_slave_in0_sync) begin
                                                                state_r <= 4'h3;
                                                              end else begin
                                                                if (_T_401) begin
                                                                  if (_T_404) begin
                                                                    if (io_slave_in0_sync) begin
                                                                      state_r <= 4'h3;
                                                                    end else begin
                                                                      if (_T_390) begin
                                                                        if (io_slave_out0_sync) begin
                                                                          state_r <= 4'h2;
                                                                        end else begin
                                                                          if (_T_97) begin
                                                                            if (_T_98) begin
                                                                              if (_T_163) begin
                                                                                if (_T_345) begin
                                                                                  if (io_master_in_sync) begin
                                                                                    state_r <= 4'h8;
                                                                                  end else begin
                                                                                    if (_T_97) begin
                                                                                      if (_T_100) begin
                                                                                        if (_T_163) begin
                                                                                          if (_T_345) begin
                                                                                            if (io_master_in_sync) begin
                                                                                              state_r <= 4'h8;
                                                                                            end else begin
                                                                                              if (_T_97) begin
                                                                                                if (_T_98) begin
                                                                                                  if (_T_154) begin
                                                                                                    if (_T_293) begin
                                                                                                      if (io_master_in_sync) begin
                                                                                                        state_r <= 4'h6;
                                                                                                      end else begin
                                                                                                        if (_T_97) begin
                                                                                                          if (_T_100) begin
                                                                                                            if (_T_154) begin
                                                                                                              if (_T_293) begin
                                                                                                                if (io_master_in_sync) begin
                                                                                                                  state_r <= 4'h6;
                                                                                                                end else begin
                                                                                                                  if (_T_97) begin
                                                                                                                    if (_T_98) begin
                                                                                                                      if (_T_145) begin
                                                                                                                        if (_T_241) begin
                                                                                                                          if (io_master_in_sync) begin
                                                                                                                            state_r <= 4'h4;
                                                                                                                          end else begin
                                                                                                                            if (_T_97) begin
                                                                                                                              if (_T_100) begin
                                                                                                                                if (_T_145) begin
                                                                                                                                  if (_T_241) begin
                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                      state_r <= 4'h4;
                                                                                                                                    end else begin
                                                                                                                                      if (_T_97) begin
                                                                                                                                        if (_T_143) begin
                                                                                                                                          if (_T_152) begin
                                                                                                                                            if (_T_161) begin
                                                                                                                                              if (_T_170) begin
                                                                                                                                                if (_T_221) begin
                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                    state_r <= 4'h3;
                                                                                                                                                  end else begin
                                                                                                                                                    if (_T_97) begin
                                                                                                                                                      if (_T_98) begin
                                                                                                                                                        if (_T_143) begin
                                                                                                                                                          if (_T_152) begin
                                                                                                                                                            if (_T_161) begin
                                                                                                                                                              if (_T_170) begin
                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                  state_r <= 4'h3;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (_T_97) begin
                                                                                                                                                                    if (_T_98) begin
                                                                                                                                                                      if (_T_102) begin
                                                                                                                                                                        if (_T_104) begin
                                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                                            state_r <= 4'h1;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (_T_97) begin
                                                                                                                                                                              if (_T_100) begin
                                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                                      state_r <= 4'h1;
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (_T_97) begin
                                                                                                                                                                            if (_T_100) begin
                                                                                                                                                                              if (_T_102) begin
                                                                                                                                                                                if (_T_104) begin
                                                                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                                                                    state_r <= 4'h1;
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (_T_97) begin
                                                                                                                                                                          if (_T_100) begin
                                                                                                                                                                            if (_T_102) begin
                                                                                                                                                                              if (_T_104) begin
                                                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                                                  state_r <= 4'h1;
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (_T_97) begin
                                                                                                                                                                        if (_T_100) begin
                                                                                                                                                                          if (_T_102) begin
                                                                                                                                                                            if (_T_104) begin
                                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                                state_r <= 4'h1;
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    state_r <= _GEN_76;
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                if (_T_97) begin
                                                                                                                                                                  if (_T_98) begin
                                                                                                                                                                    if (_T_102) begin
                                                                                                                                                                      if (_T_104) begin
                                                                                                                                                                        if (io_master_in_sync) begin
                                                                                                                                                                          state_r <= 4'h1;
                                                                                                                                                                        end else begin
                                                                                                                                                                          state_r <= _GEN_76;
                                                                                                                                                                        end
                                                                                                                                                                      end else begin
                                                                                                                                                                        state_r <= _GEN_76;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      state_r <= _GEN_76;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    state_r <= _GEN_76;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  state_r <= _GEN_76;
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              if (_T_97) begin
                                                                                                                                                                if (_T_98) begin
                                                                                                                                                                  if (_T_102) begin
                                                                                                                                                                    if (_T_104) begin
                                                                                                                                                                      if (io_master_in_sync) begin
                                                                                                                                                                        state_r <= 4'h1;
                                                                                                                                                                      end else begin
                                                                                                                                                                        state_r <= _GEN_76;
                                                                                                                                                                      end
                                                                                                                                                                    end else begin
                                                                                                                                                                      state_r <= _GEN_76;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    state_r <= _GEN_76;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  state_r <= _GEN_76;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                state_r <= _GEN_76;
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            if (_T_97) begin
                                                                                                                                                              if (_T_98) begin
                                                                                                                                                                if (_T_102) begin
                                                                                                                                                                  if (_T_104) begin
                                                                                                                                                                    if (io_master_in_sync) begin
                                                                                                                                                                      state_r <= 4'h1;
                                                                                                                                                                    end else begin
                                                                                                                                                                      state_r <= _GEN_76;
                                                                                                                                                                    end
                                                                                                                                                                  end else begin
                                                                                                                                                                    state_r <= _GEN_76;
                                                                                                                                                                  end
                                                                                                                                                                end else begin
                                                                                                                                                                  state_r <= _GEN_76;
                                                                                                                                                                end
                                                                                                                                                              end else begin
                                                                                                                                                                state_r <= _GEN_76;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              state_r <= _GEN_76;
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          state_r <= _GEN_171;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        state_r <= _GEN_171;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      state_r <= _GEN_171;
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  if (_T_97) begin
                                                                                                                                                    if (_T_98) begin
                                                                                                                                                      if (_T_143) begin
                                                                                                                                                        if (_T_152) begin
                                                                                                                                                          if (_T_161) begin
                                                                                                                                                            if (_T_170) begin
                                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                                state_r <= 4'h3;
                                                                                                                                                              end else begin
                                                                                                                                                                state_r <= _GEN_171;
                                                                                                                                                              end
                                                                                                                                                            end else begin
                                                                                                                                                              state_r <= _GEN_171;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            state_r <= _GEN_171;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          state_r <= _GEN_171;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        state_r <= _GEN_171;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      state_r <= _GEN_171;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    state_r <= _GEN_171;
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                if (_T_97) begin
                                                                                                                                                  if (_T_98) begin
                                                                                                                                                    if (_T_143) begin
                                                                                                                                                      if (_T_152) begin
                                                                                                                                                        if (_T_161) begin
                                                                                                                                                          if (_T_170) begin
                                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                                              state_r <= 4'h3;
                                                                                                                                                            end else begin
                                                                                                                                                              state_r <= _GEN_171;
                                                                                                                                                            end
                                                                                                                                                          end else begin
                                                                                                                                                            state_r <= _GEN_171;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          state_r <= _GEN_171;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        state_r <= _GEN_171;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      state_r <= _GEN_171;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    state_r <= _GEN_171;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  state_r <= _GEN_171;
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              if (_T_97) begin
                                                                                                                                                if (_T_98) begin
                                                                                                                                                  if (_T_143) begin
                                                                                                                                                    if (_T_152) begin
                                                                                                                                                      if (_T_161) begin
                                                                                                                                                        if (_T_170) begin
                                                                                                                                                          if (io_master_in_sync) begin
                                                                                                                                                            state_r <= 4'h3;
                                                                                                                                                          end else begin
                                                                                                                                                            state_r <= _GEN_171;
                                                                                                                                                          end
                                                                                                                                                        end else begin
                                                                                                                                                          state_r <= _GEN_171;
                                                                                                                                                        end
                                                                                                                                                      end else begin
                                                                                                                                                        state_r <= _GEN_171;
                                                                                                                                                      end
                                                                                                                                                    end else begin
                                                                                                                                                      state_r <= _GEN_171;
                                                                                                                                                    end
                                                                                                                                                  end else begin
                                                                                                                                                    state_r <= _GEN_171;
                                                                                                                                                  end
                                                                                                                                                end else begin
                                                                                                                                                  state_r <= _GEN_171;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                state_r <= _GEN_171;
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            state_r <= _GEN_298;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          state_r <= _GEN_298;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        state_r <= _GEN_298;
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    if (_T_97) begin
                                                                                                                                      if (_T_143) begin
                                                                                                                                        if (_T_152) begin
                                                                                                                                          if (_T_161) begin
                                                                                                                                            if (_T_170) begin
                                                                                                                                              if (_T_221) begin
                                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                                  state_r <= 4'h3;
                                                                                                                                                end else begin
                                                                                                                                                  state_r <= _GEN_298;
                                                                                                                                                end
                                                                                                                                              end else begin
                                                                                                                                                state_r <= _GEN_298;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              state_r <= _GEN_298;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            state_r <= _GEN_298;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          state_r <= _GEN_298;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        state_r <= _GEN_298;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      state_r <= _GEN_298;
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  if (_T_97) begin
                                                                                                                                    if (_T_143) begin
                                                                                                                                      if (_T_152) begin
                                                                                                                                        if (_T_161) begin
                                                                                                                                          if (_T_170) begin
                                                                                                                                            if (_T_221) begin
                                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                                state_r <= 4'h3;
                                                                                                                                              end else begin
                                                                                                                                                state_r <= _GEN_298;
                                                                                                                                              end
                                                                                                                                            end else begin
                                                                                                                                              state_r <= _GEN_298;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            state_r <= _GEN_298;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          state_r <= _GEN_298;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        state_r <= _GEN_298;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      state_r <= _GEN_298;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    state_r <= _GEN_298;
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                if (_T_97) begin
                                                                                                                                  if (_T_143) begin
                                                                                                                                    if (_T_152) begin
                                                                                                                                      if (_T_161) begin
                                                                                                                                        if (_T_170) begin
                                                                                                                                          if (_T_221) begin
                                                                                                                                            if (io_master_in_sync) begin
                                                                                                                                              state_r <= 4'h3;
                                                                                                                                            end else begin
                                                                                                                                              state_r <= _GEN_298;
                                                                                                                                            end
                                                                                                                                          end else begin
                                                                                                                                            state_r <= _GEN_298;
                                                                                                                                          end
                                                                                                                                        end else begin
                                                                                                                                          state_r <= _GEN_298;
                                                                                                                                        end
                                                                                                                                      end else begin
                                                                                                                                        state_r <= _GEN_298;
                                                                                                                                      end
                                                                                                                                    end else begin
                                                                                                                                      state_r <= _GEN_298;
                                                                                                                                    end
                                                                                                                                  end else begin
                                                                                                                                    state_r <= _GEN_298;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  state_r <= _GEN_298;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              state_r <= _GEN_424;
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          if (_T_97) begin
                                                                                                                            if (_T_100) begin
                                                                                                                              if (_T_145) begin
                                                                                                                                if (_T_241) begin
                                                                                                                                  if (io_master_in_sync) begin
                                                                                                                                    state_r <= 4'h4;
                                                                                                                                  end else begin
                                                                                                                                    state_r <= _GEN_424;
                                                                                                                                  end
                                                                                                                                end else begin
                                                                                                                                  state_r <= _GEN_424;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                state_r <= _GEN_424;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              state_r <= _GEN_424;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            state_r <= _GEN_424;
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        if (_T_97) begin
                                                                                                                          if (_T_100) begin
                                                                                                                            if (_T_145) begin
                                                                                                                              if (_T_241) begin
                                                                                                                                if (io_master_in_sync) begin
                                                                                                                                  state_r <= 4'h4;
                                                                                                                                end else begin
                                                                                                                                  state_r <= _GEN_424;
                                                                                                                                end
                                                                                                                              end else begin
                                                                                                                                state_r <= _GEN_424;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              state_r <= _GEN_424;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            state_r <= _GEN_424;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          state_r <= _GEN_424;
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      if (_T_97) begin
                                                                                                                        if (_T_100) begin
                                                                                                                          if (_T_145) begin
                                                                                                                            if (_T_241) begin
                                                                                                                              if (io_master_in_sync) begin
                                                                                                                                state_r <= 4'h4;
                                                                                                                              end else begin
                                                                                                                                state_r <= _GEN_424;
                                                                                                                              end
                                                                                                                            end else begin
                                                                                                                              state_r <= _GEN_424;
                                                                                                                            end
                                                                                                                          end else begin
                                                                                                                            state_r <= _GEN_424;
                                                                                                                          end
                                                                                                                        end else begin
                                                                                                                          state_r <= _GEN_424;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        state_r <= _GEN_424;
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    state_r <= _GEN_518;
                                                                                                                  end
                                                                                                                end
                                                                                                              end else begin
                                                                                                                if (_T_97) begin
                                                                                                                  if (_T_98) begin
                                                                                                                    if (_T_145) begin
                                                                                                                      if (_T_241) begin
                                                                                                                        if (io_master_in_sync) begin
                                                                                                                          state_r <= 4'h4;
                                                                                                                        end else begin
                                                                                                                          state_r <= _GEN_518;
                                                                                                                        end
                                                                                                                      end else begin
                                                                                                                        state_r <= _GEN_518;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      state_r <= _GEN_518;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    state_r <= _GEN_518;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  state_r <= _GEN_518;
                                                                                                                end
                                                                                                              end
                                                                                                            end else begin
                                                                                                              if (_T_97) begin
                                                                                                                if (_T_98) begin
                                                                                                                  if (_T_145) begin
                                                                                                                    if (_T_241) begin
                                                                                                                      if (io_master_in_sync) begin
                                                                                                                        state_r <= 4'h4;
                                                                                                                      end else begin
                                                                                                                        state_r <= _GEN_518;
                                                                                                                      end
                                                                                                                    end else begin
                                                                                                                      state_r <= _GEN_518;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    state_r <= _GEN_518;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  state_r <= _GEN_518;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                state_r <= _GEN_518;
                                                                                                              end
                                                                                                            end
                                                                                                          end else begin
                                                                                                            if (_T_97) begin
                                                                                                              if (_T_98) begin
                                                                                                                if (_T_145) begin
                                                                                                                  if (_T_241) begin
                                                                                                                    if (io_master_in_sync) begin
                                                                                                                      state_r <= 4'h4;
                                                                                                                    end else begin
                                                                                                                      state_r <= _GEN_518;
                                                                                                                    end
                                                                                                                  end else begin
                                                                                                                    state_r <= _GEN_518;
                                                                                                                  end
                                                                                                                end else begin
                                                                                                                  state_r <= _GEN_518;
                                                                                                                end
                                                                                                              end else begin
                                                                                                                state_r <= _GEN_518;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              state_r <= _GEN_518;
                                                                                                            end
                                                                                                          end
                                                                                                        end else begin
                                                                                                          state_r <= _GEN_613;
                                                                                                        end
                                                                                                      end
                                                                                                    end else begin
                                                                                                      if (_T_97) begin
                                                                                                        if (_T_100) begin
                                                                                                          if (_T_154) begin
                                                                                                            if (_T_293) begin
                                                                                                              if (io_master_in_sync) begin
                                                                                                                state_r <= 4'h6;
                                                                                                              end else begin
                                                                                                                state_r <= _GEN_613;
                                                                                                              end
                                                                                                            end else begin
                                                                                                              state_r <= _GEN_613;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            state_r <= _GEN_613;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          state_r <= _GEN_613;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        state_r <= _GEN_613;
                                                                                                      end
                                                                                                    end
                                                                                                  end else begin
                                                                                                    if (_T_97) begin
                                                                                                      if (_T_100) begin
                                                                                                        if (_T_154) begin
                                                                                                          if (_T_293) begin
                                                                                                            if (io_master_in_sync) begin
                                                                                                              state_r <= 4'h6;
                                                                                                            end else begin
                                                                                                              state_r <= _GEN_613;
                                                                                                            end
                                                                                                          end else begin
                                                                                                            state_r <= _GEN_613;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          state_r <= _GEN_613;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        state_r <= _GEN_613;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      state_r <= _GEN_613;
                                                                                                    end
                                                                                                  end
                                                                                                end else begin
                                                                                                  if (_T_97) begin
                                                                                                    if (_T_100) begin
                                                                                                      if (_T_154) begin
                                                                                                        if (_T_293) begin
                                                                                                          if (io_master_in_sync) begin
                                                                                                            state_r <= 4'h6;
                                                                                                          end else begin
                                                                                                            state_r <= _GEN_613;
                                                                                                          end
                                                                                                        end else begin
                                                                                                          state_r <= _GEN_613;
                                                                                                        end
                                                                                                      end else begin
                                                                                                        state_r <= _GEN_613;
                                                                                                      end
                                                                                                    end else begin
                                                                                                      state_r <= _GEN_613;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    state_r <= _GEN_613;
                                                                                                  end
                                                                                                end
                                                                                              end else begin
                                                                                                state_r <= _GEN_708;
                                                                                              end
                                                                                            end
                                                                                          end else begin
                                                                                            if (_T_97) begin
                                                                                              if (_T_98) begin
                                                                                                if (_T_154) begin
                                                                                                  if (_T_293) begin
                                                                                                    if (io_master_in_sync) begin
                                                                                                      state_r <= 4'h6;
                                                                                                    end else begin
                                                                                                      state_r <= _GEN_708;
                                                                                                    end
                                                                                                  end else begin
                                                                                                    state_r <= _GEN_708;
                                                                                                  end
                                                                                                end else begin
                                                                                                  state_r <= _GEN_708;
                                                                                                end
                                                                                              end else begin
                                                                                                state_r <= _GEN_708;
                                                                                              end
                                                                                            end else begin
                                                                                              state_r <= _GEN_708;
                                                                                            end
                                                                                          end
                                                                                        end else begin
                                                                                          if (_T_97) begin
                                                                                            if (_T_98) begin
                                                                                              if (_T_154) begin
                                                                                                if (_T_293) begin
                                                                                                  if (io_master_in_sync) begin
                                                                                                    state_r <= 4'h6;
                                                                                                  end else begin
                                                                                                    state_r <= _GEN_708;
                                                                                                  end
                                                                                                end else begin
                                                                                                  state_r <= _GEN_708;
                                                                                                end
                                                                                              end else begin
                                                                                                state_r <= _GEN_708;
                                                                                              end
                                                                                            end else begin
                                                                                              state_r <= _GEN_708;
                                                                                            end
                                                                                          end else begin
                                                                                            state_r <= _GEN_708;
                                                                                          end
                                                                                        end
                                                                                      end else begin
                                                                                        if (_T_97) begin
                                                                                          if (_T_98) begin
                                                                                            if (_T_154) begin
                                                                                              if (_T_293) begin
                                                                                                if (io_master_in_sync) begin
                                                                                                  state_r <= 4'h6;
                                                                                                end else begin
                                                                                                  state_r <= _GEN_708;
                                                                                                end
                                                                                              end else begin
                                                                                                state_r <= _GEN_708;
                                                                                              end
                                                                                            end else begin
                                                                                              state_r <= _GEN_708;
                                                                                            end
                                                                                          end else begin
                                                                                            state_r <= _GEN_708;
                                                                                          end
                                                                                        end else begin
                                                                                          state_r <= _GEN_708;
                                                                                        end
                                                                                      end
                                                                                    end else begin
                                                                                      state_r <= _GEN_803;
                                                                                    end
                                                                                  end
                                                                                end else begin
                                                                                  if (_T_97) begin
                                                                                    if (_T_100) begin
                                                                                      if (_T_163) begin
                                                                                        if (_T_345) begin
                                                                                          if (io_master_in_sync) begin
                                                                                            state_r <= 4'h8;
                                                                                          end else begin
                                                                                            state_r <= _GEN_803;
                                                                                          end
                                                                                        end else begin
                                                                                          state_r <= _GEN_803;
                                                                                        end
                                                                                      end else begin
                                                                                        state_r <= _GEN_803;
                                                                                      end
                                                                                    end else begin
                                                                                      state_r <= _GEN_803;
                                                                                    end
                                                                                  end else begin
                                                                                    state_r <= _GEN_803;
                                                                                  end
                                                                                end
                                                                              end else begin
                                                                                if (_T_97) begin
                                                                                  if (_T_100) begin
                                                                                    if (_T_163) begin
                                                                                      if (_T_345) begin
                                                                                        if (io_master_in_sync) begin
                                                                                          state_r <= 4'h8;
                                                                                        end else begin
                                                                                          state_r <= _GEN_803;
                                                                                        end
                                                                                      end else begin
                                                                                        state_r <= _GEN_803;
                                                                                      end
                                                                                    end else begin
                                                                                      state_r <= _GEN_803;
                                                                                    end
                                                                                  end else begin
                                                                                    state_r <= _GEN_803;
                                                                                  end
                                                                                end else begin
                                                                                  state_r <= _GEN_803;
                                                                                end
                                                                              end
                                                                            end else begin
                                                                              if (_T_97) begin
                                                                                if (_T_100) begin
                                                                                  if (_T_163) begin
                                                                                    if (_T_345) begin
                                                                                      if (io_master_in_sync) begin
                                                                                        state_r <= 4'h8;
                                                                                      end else begin
                                                                                        state_r <= _GEN_803;
                                                                                      end
                                                                                    end else begin
                                                                                      state_r <= _GEN_803;
                                                                                    end
                                                                                  end else begin
                                                                                    state_r <= _GEN_803;
                                                                                  end
                                                                                end else begin
                                                                                  state_r <= _GEN_803;
                                                                                end
                                                                              end else begin
                                                                                state_r <= _GEN_803;
                                                                              end
                                                                            end
                                                                          end else begin
                                                                            state_r <= _GEN_898;
                                                                          end
                                                                        end
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  state_r <= 4'h8;
                                                                                end else begin
                                                                                  state_r <= _GEN_898;
                                                                                end
                                                                              end else begin
                                                                                state_r <= _GEN_898;
                                                                              end
                                                                            end else begin
                                                                              state_r <= _GEN_898;
                                                                            end
                                                                          end else begin
                                                                            state_r <= _GEN_898;
                                                                          end
                                                                        end else begin
                                                                          state_r <= _GEN_898;
                                                                        end
                                                                      end
                                                                    end
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        state_r <= 4'h2;
                                                                      end else begin
                                                                        if (_T_97) begin
                                                                          if (_T_98) begin
                                                                            if (_T_163) begin
                                                                              if (_T_345) begin
                                                                                if (io_master_in_sync) begin
                                                                                  state_r <= 4'h8;
                                                                                end else begin
                                                                                  state_r <= _GEN_898;
                                                                                end
                                                                              end else begin
                                                                                state_r <= _GEN_898;
                                                                              end
                                                                            end else begin
                                                                              state_r <= _GEN_898;
                                                                            end
                                                                          end else begin
                                                                            state_r <= _GEN_898;
                                                                          end
                                                                        end else begin
                                                                          state_r <= _GEN_898;
                                                                        end
                                                                      end
                                                                    end else begin
                                                                      if (_T_97) begin
                                                                        if (_T_98) begin
                                                                          if (_T_163) begin
                                                                            if (_T_345) begin
                                                                              if (io_master_in_sync) begin
                                                                                state_r <= 4'h8;
                                                                              end else begin
                                                                                state_r <= _GEN_898;
                                                                              end
                                                                            end else begin
                                                                              state_r <= _GEN_898;
                                                                            end
                                                                          end else begin
                                                                            state_r <= _GEN_898;
                                                                          end
                                                                        end else begin
                                                                          state_r <= _GEN_898;
                                                                        end
                                                                      end else begin
                                                                        state_r <= _GEN_898;
                                                                      end
                                                                    end
                                                                  end
                                                                end else begin
                                                                  if (_T_390) begin
                                                                    if (io_slave_out0_sync) begin
                                                                      state_r <= 4'h2;
                                                                    end else begin
                                                                      state_r <= _GEN_993;
                                                                    end
                                                                  end else begin
                                                                    state_r <= _GEN_993;
                                                                  end
                                                                end
                                                              end
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    state_r <= 4'h3;
                                                                  end else begin
                                                                    if (_T_390) begin
                                                                      if (io_slave_out0_sync) begin
                                                                        state_r <= 4'h2;
                                                                      end else begin
                                                                        state_r <= _GEN_993;
                                                                      end
                                                                    end else begin
                                                                      state_r <= _GEN_993;
                                                                    end
                                                                  end
                                                                end else begin
                                                                  state_r <= _GEN_1028;
                                                                end
                                                              end else begin
                                                                state_r <= _GEN_1028;
                                                              end
                                                            end
                                                          end else begin
                                                            if (_T_401) begin
                                                              if (_T_404) begin
                                                                if (io_slave_in0_sync) begin
                                                                  state_r <= 4'h3;
                                                                end else begin
                                                                  state_r <= _GEN_1028;
                                                                end
                                                              end else begin
                                                                state_r <= _GEN_1028;
                                                              end
                                                            end else begin
                                                              state_r <= _GEN_1028;
                                                            end
                                                          end
                                                        end
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              state_r <= 4'h3;
                                                            end else begin
                                                              if (_T_401) begin
                                                                if (_T_404) begin
                                                                  if (io_slave_in0_sync) begin
                                                                    state_r <= 4'h3;
                                                                  end else begin
                                                                    state_r <= _GEN_1028;
                                                                  end
                                                                end else begin
                                                                  state_r <= _GEN_1028;
                                                                end
                                                              end else begin
                                                                state_r <= _GEN_1028;
                                                              end
                                                            end
                                                          end else begin
                                                            state_r <= _GEN_1080;
                                                          end
                                                        end else begin
                                                          state_r <= _GEN_1080;
                                                        end
                                                      end
                                                    end
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        state_r <= 4'h0;
                                                      end else begin
                                                        if (_T_401) begin
                                                          if (_T_402) begin
                                                            if (io_slave_in0_sync) begin
                                                              state_r <= 4'h3;
                                                            end else begin
                                                              state_r <= _GEN_1080;
                                                            end
                                                          end else begin
                                                            state_r <= _GEN_1080;
                                                          end
                                                        end else begin
                                                          state_r <= _GEN_1080;
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_401) begin
                                                        if (_T_402) begin
                                                          if (io_slave_in0_sync) begin
                                                            state_r <= 4'h3;
                                                          end else begin
                                                            state_r <= _GEN_1080;
                                                          end
                                                        end else begin
                                                          state_r <= _GEN_1080;
                                                        end
                                                      end else begin
                                                        state_r <= _GEN_1080;
                                                      end
                                                    end
                                                  end
                                                end
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    state_r <= 4'h5;
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (io_master_out_sync) begin
                                                        state_r <= 4'h0;
                                                      end else begin
                                                        state_r <= _GEN_1134;
                                                      end
                                                    end else begin
                                                      state_r <= _GEN_1134;
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_429) begin
                                                    if (io_master_out_sync) begin
                                                      state_r <= 4'h0;
                                                    end else begin
                                                      state_r <= _GEN_1134;
                                                    end
                                                  end else begin
                                                    state_r <= _GEN_1134;
                                                  end
                                                end
                                              end
                                            end else begin
                                              if (_T_440) begin
                                                if (io_slave_out1_sync) begin
                                                  state_r <= 4'h5;
                                                end else begin
                                                  state_r <= _GEN_1168;
                                                end
                                              end else begin
                                                state_r <= _GEN_1168;
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                state_r <= 4'h3;
                                              end else begin
                                                if (_T_440) begin
                                                  if (io_slave_out1_sync) begin
                                                    state_r <= 4'h5;
                                                  end else begin
                                                    state_r <= _GEN_1168;
                                                  end
                                                end else begin
                                                  state_r <= _GEN_1168;
                                                end
                                              end
                                            end else begin
                                              state_r <= _GEN_1200;
                                            end
                                          end else begin
                                            state_r <= _GEN_1200;
                                          end
                                        end
                                      end else begin
                                        if (_T_451) begin
                                          if (_T_404) begin
                                            if (io_slave_in1_sync) begin
                                              state_r <= 4'h3;
                                            end else begin
                                              state_r <= _GEN_1200;
                                            end
                                          end else begin
                                            state_r <= _GEN_1200;
                                          end
                                        end else begin
                                          state_r <= _GEN_1200;
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          state_r <= 4'h3;
                                        end else begin
                                          if (_T_451) begin
                                            if (_T_404) begin
                                              if (io_slave_in1_sync) begin
                                                state_r <= 4'h3;
                                              end else begin
                                                state_r <= _GEN_1200;
                                              end
                                            end else begin
                                              state_r <= _GEN_1200;
                                            end
                                          end else begin
                                            state_r <= _GEN_1200;
                                          end
                                        end
                                      end else begin
                                        state_r <= _GEN_1252;
                                      end
                                    end else begin
                                      state_r <= _GEN_1252;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    state_r <= 4'h7;
                                  end else begin
                                    if (_T_451) begin
                                      if (_T_402) begin
                                        if (io_slave_in1_sync) begin
                                          state_r <= 4'h3;
                                        end else begin
                                          state_r <= _GEN_1252;
                                        end
                                      end else begin
                                        state_r <= _GEN_1252;
                                      end
                                    end else begin
                                      state_r <= _GEN_1252;
                                    end
                                  end
                                end else begin
                                  if (_T_451) begin
                                    if (_T_402) begin
                                      if (io_slave_in1_sync) begin
                                        state_r <= 4'h3;
                                      end else begin
                                        state_r <= _GEN_1252;
                                      end
                                    end else begin
                                      state_r <= _GEN_1252;
                                    end
                                  end else begin
                                    state_r <= _GEN_1252;
                                  end
                                end
                              end
                            end else begin
                              if (_T_479) begin
                                if (io_slave_out2_sync) begin
                                  state_r <= 4'h7;
                                end else begin
                                  state_r <= _GEN_1306;
                                end
                              end else begin
                                state_r <= _GEN_1306;
                              end
                            end
                          end
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                state_r <= 4'h3;
                              end else begin
                                if (_T_479) begin
                                  if (io_slave_out2_sync) begin
                                    state_r <= 4'h7;
                                  end else begin
                                    state_r <= _GEN_1306;
                                  end
                                end else begin
                                  state_r <= _GEN_1306;
                                end
                              end
                            end else begin
                              state_r <= _GEN_1340;
                            end
                          end else begin
                            state_r <= _GEN_1340;
                          end
                        end
                      end else begin
                        if (_T_490) begin
                          if (_T_404) begin
                            if (io_slave_in2_sync) begin
                              state_r <= 4'h3;
                            end else begin
                              state_r <= _GEN_1340;
                            end
                          end else begin
                            state_r <= _GEN_1340;
                          end
                        end else begin
                          state_r <= _GEN_1340;
                        end
                      end
                    end
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          state_r <= 4'h3;
                        end else begin
                          if (_T_490) begin
                            if (_T_404) begin
                              if (io_slave_in2_sync) begin
                                state_r <= 4'h3;
                              end else begin
                                state_r <= _GEN_1340;
                              end
                            end else begin
                              state_r <= _GEN_1340;
                            end
                          end else begin
                            state_r <= _GEN_1340;
                          end
                        end
                      end else begin
                        state_r <= _GEN_1392;
                      end
                    end else begin
                      state_r <= _GEN_1392;
                    end
                  end
                end
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    state_r <= 4'h9;
                  end else begin
                    if (_T_490) begin
                      if (_T_402) begin
                        if (io_slave_in2_sync) begin
                          state_r <= 4'h3;
                        end else begin
                          state_r <= _GEN_1392;
                        end
                      end else begin
                        state_r <= _GEN_1392;
                      end
                    end else begin
                      state_r <= _GEN_1392;
                    end
                  end
                end else begin
                  if (_T_490) begin
                    if (_T_402) begin
                      if (io_slave_in2_sync) begin
                        state_r <= 4'h3;
                      end else begin
                        state_r <= _GEN_1392;
                      end
                    end else begin
                      state_r <= _GEN_1392;
                    end
                  end else begin
                    state_r <= _GEN_1392;
                  end
                end
              end
            end else begin
              if (_T_518) begin
                if (io_slave_out3_sync) begin
                  state_r <= 4'h9;
                end else begin
                  state_r <= _GEN_1446;
                end
              end else begin
                state_r <= _GEN_1446;
              end
            end
          end
        end else begin
          if (_T_529) begin
            if (_T_404) begin
              if (io_slave_in3_sync) begin
                state_r <= 4'h3;
              end else begin
                if (_T_518) begin
                  if (io_slave_out3_sync) begin
                    state_r <= 4'h9;
                  end else begin
                    state_r <= _GEN_1446;
                  end
                end else begin
                  state_r <= _GEN_1446;
                end
              end
            end else begin
              state_r <= _GEN_1480;
            end
          end else begin
            state_r <= _GEN_1480;
          end
        end
      end else begin
        if (_T_529) begin
          if (_T_404) begin
            if (io_slave_in3_sync) begin
              state_r <= 4'h3;
            end else begin
              state_r <= _GEN_1480;
            end
          end else begin
            state_r <= _GEN_1480;
          end
        end else begin
          state_r <= _GEN_1480;
        end
      end
    end
  end
endmodule
