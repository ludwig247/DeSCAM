package testbasic2_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic2_SECTIONS;

endpackage
