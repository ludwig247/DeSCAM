library ieee;
use IEEE.numeric_std.all;

package TestFunction1_types is
type TestFunction1_SECTIONS is (run);
end package TestFunction1_types;
