library ieee;
use IEEE.numeric_std.all;

package TestBasic0_types is
type TestBasic0_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic0_types;
