library ieee;
use IEEE.numeric_std.all;

package TestFunction2_types is
type TestFunction2_SECTIONS is (run);
end package TestFunction2_types;
