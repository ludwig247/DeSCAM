library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package sc_main_types is
-- No local datatypes implemented!


end package sc_main_types;