
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_CPU is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
subtype bool is BOOLEAN range FALSE to TRUE ;
   
   -- Declarations for conversion functions.
   function std_logic_to_bool(arg : in std_logic) return bool;
   function bool_to_std_logic(arg : in bool) return std_logic;

end CONV_PACK_CPU;

package body CONV_PACK_CPU is
   
   -- std_logic to enum type function
   function std_logic_to_bool(arg : in std_logic) return bool is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when '0' => return FALSE;
         when '1' => return TRUE;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return FALSE;
      end case;
   end;
   
   -- enum type to std_logic function
   function bool_to_std_logic(arg : in bool) return std_logic is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when FALSE => return '0';
         when TRUE => return '1';
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return '0';
      end case;
   end;

end CONV_PACK_CPU;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_35 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_35;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_34 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_34;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_33 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_33;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_32 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_32;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_31 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_31;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_30 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_30;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_29 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_29;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_28 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_28;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_27 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_27;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_26 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_26;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_25 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_25;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_24 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_24;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_23 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_23;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_22 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_22;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_21 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_21;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_20 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_20;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_19 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_19;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_18 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_18;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_17 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_17;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_16 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_16;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_15 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_15;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_14 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_14;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_13 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_13;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_12 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_12;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_11 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_11;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_10 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_10;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_9 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_9;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_8 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_8;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_7 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_7;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_6 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_6;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_5 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_5;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_4 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_4;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_3 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_3;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_2 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_2;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_1 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_1;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_36 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_36;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_0;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net6517 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net6517);
   main_gate : AND2_X1 port map( A1 => net6517, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity CPU is

   port( clk, rst : in std_logic;  fromMemoryPortxLOADEDDATAx : in 
         std_logic_vector (31 downto 0);  fromMemoryPort_sync : in bool;  
         fromMemoryPort_notify : out bool;  toMemoryPort_sync : in bool;  
         toMemoryPort_notify : out bool;  toMemoryPortxADDRINxx31x, 
         toMemoryPortxADDRINxx30x, toMemoryPortxADDRINxx29x, 
         toMemoryPortxADDRINxx28x, toMemoryPortxADDRINxx27x, 
         toMemoryPortxADDRINxx26x, toMemoryPortxADDRINxx25x, 
         toMemoryPortxADDRINxx24x, toMemoryPortxADDRINxx23x, 
         toMemoryPortxADDRINxx22x, toMemoryPortxADDRINxx21x, 
         toMemoryPortxADDRINxx20x, toMemoryPortxADDRINxx19x, 
         toMemoryPortxADDRINxx18x, toMemoryPortxADDRINxx17x, 
         toMemoryPortxADDRINxx16x, toMemoryPortxADDRINxx15x, 
         toMemoryPortxADDRINxx14x, toMemoryPortxADDRINxx13x, 
         toMemoryPortxADDRINxx12x, toMemoryPortxADDRINxx11x, 
         toMemoryPortxADDRINxx10x, toMemoryPortxADDRINxx9x, 
         toMemoryPortxADDRINxx8x, toMemoryPortxADDRINxx7x, 
         toMemoryPortxADDRINxx6x, toMemoryPortxADDRINxx5x, 
         toMemoryPortxADDRINxx4x, toMemoryPortxADDRINxx3x, 
         toMemoryPortxADDRINxx2x, toMemoryPortxADDRINxx1x, 
         toMemoryPortxADDRINxx0x, toMemoryPortxDATAINxx31x, 
         toMemoryPortxDATAINxx30x, toMemoryPortxDATAINxx29x, 
         toMemoryPortxDATAINxx28x, toMemoryPortxDATAINxx27x, 
         toMemoryPortxDATAINxx26x, toMemoryPortxDATAINxx25x, 
         toMemoryPortxDATAINxx24x, toMemoryPortxDATAINxx23x, 
         toMemoryPortxDATAINxx22x, toMemoryPortxDATAINxx21x, 
         toMemoryPortxDATAINxx20x, toMemoryPortxDATAINxx19x, 
         toMemoryPortxDATAINxx18x, toMemoryPortxDATAINxx17x, 
         toMemoryPortxDATAINxx16x, toMemoryPortxDATAINxx15x, 
         toMemoryPortxDATAINxx14x, toMemoryPortxDATAINxx13x, 
         toMemoryPortxDATAINxx12x, toMemoryPortxDATAINxx11x, 
         toMemoryPortxDATAINxx10x, toMemoryPortxDATAINxx9x, 
         toMemoryPortxDATAINxx8x, toMemoryPortxDATAINxx7x, 
         toMemoryPortxDATAINxx6x, toMemoryPortxDATAINxx5x, 
         toMemoryPortxDATAINxx4x, toMemoryPortxDATAINxx3x, 
         toMemoryPortxDATAINxx2x, toMemoryPortxDATAINxx1x, 
         toMemoryPortxDATAINxx0x, toMemoryPortxMASKxx2x, toMemoryPortxMASKxx1x,
         toMemoryPortxMASKxx0x, toMemoryPortxREQxx1x, toMemoryPortxREQxx0x : 
         out std_logic_vector (0 to 0));

end CPU;

architecture SYN_CPU_arch of CPU is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_1
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_2
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_3
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_4
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_5
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_6
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_7
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_8
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_9
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_10
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_11
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_12
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_13
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_14
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_15
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_16
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_17
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_18
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_19
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_20
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_21
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_22
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_23
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_24
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_25
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_26
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_27
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_28
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_29
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_30
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_31
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_32
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_33
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_34
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_35
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_36
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal fromMemoryPort_sync_port, toMemoryPort_sync_port, 
      toMemoryPort_notify_port, toRegsPortxDSTxx4x, toRegsPortxDSTxx3x, 
      toRegsPortxDSTxx2x, toRegsPortxDSTxx1x, toRegsPortxDSTxx0x, 
      toRegsPortxDSTDATAxx31x, toRegsPortxDSTDATAxx30x, toRegsPortxDSTDATAxx29x
      , toRegsPortxDSTDATAxx28x, toRegsPortxDSTDATAxx27x, 
      toRegsPortxDSTDATAxx26x, toRegsPortxDSTDATAxx25x, toRegsPortxDSTDATAxx24x
      , toRegsPortxDSTDATAxx23x, toRegsPortxDSTDATAxx22x, 
      toRegsPortxDSTDATAxx21x, toRegsPortxDSTDATAxx20x, toRegsPortxDSTDATAxx19x
      , toRegsPortxDSTDATAxx18x, toRegsPortxDSTDATAxx17x, 
      toRegsPortxDSTDATAxx16x, toRegsPortxDSTDATAxx15x, toRegsPortxDSTDATAxx14x
      , toRegsPortxDSTDATAxx13x, toRegsPortxDSTDATAxx12x, 
      toRegsPortxDSTDATAxx11x, toRegsPortxDSTDATAxx10x, toRegsPortxDSTDATAxx9x,
      toRegsPortxDSTDATAxx8x, toRegsPortxDSTDATAxx7x, toRegsPortxDSTDATAxx6x, 
      toRegsPortxDSTDATAxx5x, toRegsPortxDSTDATAxx4x, toRegsPortxDSTDATAxx3x, 
      toRegsPortxDSTDATAxx2x, toRegsPortxDSTDATAxx1x, toRegsPortxDSTDATAxx0x, 
      toRegsPort_notify, fromRegsPortxREG_FILE_01xx31x, 
      fromRegsPortxREG_FILE_01xx30x, fromRegsPortxREG_FILE_01xx29x, 
      fromRegsPortxREG_FILE_01xx28x, fromRegsPortxREG_FILE_01xx27x, 
      fromRegsPortxREG_FILE_01xx26x, fromRegsPortxREG_FILE_01xx25x, 
      fromRegsPortxREG_FILE_01xx24x, fromRegsPortxREG_FILE_01xx23x, 
      fromRegsPortxREG_FILE_01xx22x, fromRegsPortxREG_FILE_01xx21x, 
      fromRegsPortxREG_FILE_01xx20x, fromRegsPortxREG_FILE_01xx19x, 
      fromRegsPortxREG_FILE_01xx18x, fromRegsPortxREG_FILE_01xx17x, 
      fromRegsPortxREG_FILE_01xx16x, fromRegsPortxREG_FILE_01xx15x, 
      fromRegsPortxREG_FILE_01xx14x, fromRegsPortxREG_FILE_01xx13x, 
      fromRegsPortxREG_FILE_01xx12x, fromRegsPortxREG_FILE_01xx11x, 
      fromRegsPortxREG_FILE_01xx10x, fromRegsPortxREG_FILE_01xx9x, 
      fromRegsPortxREG_FILE_01xx8x, fromRegsPortxREG_FILE_01xx7x, 
      fromRegsPortxREG_FILE_01xx6x, fromRegsPortxREG_FILE_01xx5x, 
      fromRegsPortxREG_FILE_01xx4x, fromRegsPortxREG_FILE_01xx3x, 
      fromRegsPortxREG_FILE_01xx2x, fromRegsPortxREG_FILE_01xx1x, 
      fromRegsPortxREG_FILE_01xx0x, fromRegsPortxREG_FILE_02xx31x, 
      fromRegsPortxREG_FILE_02xx30x, fromRegsPortxREG_FILE_02xx29x, 
      fromRegsPortxREG_FILE_02xx28x, fromRegsPortxREG_FILE_02xx27x, 
      fromRegsPortxREG_FILE_02xx26x, fromRegsPortxREG_FILE_02xx25x, 
      fromRegsPortxREG_FILE_02xx24x, fromRegsPortxREG_FILE_02xx23x, 
      fromRegsPortxREG_FILE_02xx22x, fromRegsPortxREG_FILE_02xx21x, 
      fromRegsPortxREG_FILE_02xx20x, fromRegsPortxREG_FILE_02xx19x, 
      fromRegsPortxREG_FILE_02xx18x, fromRegsPortxREG_FILE_02xx17x, 
      fromRegsPortxREG_FILE_02xx16x, fromRegsPortxREG_FILE_02xx15x, 
      fromRegsPortxREG_FILE_02xx14x, fromRegsPortxREG_FILE_02xx13x, 
      fromRegsPortxREG_FILE_02xx12x, fromRegsPortxREG_FILE_02xx11x, 
      fromRegsPortxREG_FILE_02xx10x, fromRegsPortxREG_FILE_02xx9x, 
      fromRegsPortxREG_FILE_02xx8x, fromRegsPortxREG_FILE_02xx7x, 
      fromRegsPortxREG_FILE_02xx6x, fromRegsPortxREG_FILE_02xx5x, 
      fromRegsPortxREG_FILE_02xx4x, fromRegsPortxREG_FILE_02xx3x, 
      fromRegsPortxREG_FILE_02xx2x, fromRegsPortxREG_FILE_02xx1x, 
      fromRegsPortxREG_FILE_02xx0x, fromRegsPortxREG_FILE_03xx31x, 
      fromRegsPortxREG_FILE_03xx30x, fromRegsPortxREG_FILE_03xx29x, 
      fromRegsPortxREG_FILE_03xx28x, fromRegsPortxREG_FILE_03xx27x, 
      fromRegsPortxREG_FILE_03xx26x, fromRegsPortxREG_FILE_03xx25x, 
      fromRegsPortxREG_FILE_03xx24x, fromRegsPortxREG_FILE_03xx23x, 
      fromRegsPortxREG_FILE_03xx22x, fromRegsPortxREG_FILE_03xx21x, 
      fromRegsPortxREG_FILE_03xx20x, fromRegsPortxREG_FILE_03xx19x, 
      fromRegsPortxREG_FILE_03xx18x, fromRegsPortxREG_FILE_03xx17x, 
      fromRegsPortxREG_FILE_03xx16x, fromRegsPortxREG_FILE_03xx15x, 
      fromRegsPortxREG_FILE_03xx14x, fromRegsPortxREG_FILE_03xx13x, 
      fromRegsPortxREG_FILE_03xx12x, fromRegsPortxREG_FILE_03xx11x, 
      fromRegsPortxREG_FILE_03xx10x, fromRegsPortxREG_FILE_03xx9x, 
      fromRegsPortxREG_FILE_03xx8x, fromRegsPortxREG_FILE_03xx7x, 
      fromRegsPortxREG_FILE_03xx6x, fromRegsPortxREG_FILE_03xx5x, 
      fromRegsPortxREG_FILE_03xx4x, fromRegsPortxREG_FILE_03xx3x, 
      fromRegsPortxREG_FILE_03xx2x, fromRegsPortxREG_FILE_03xx1x, 
      fromRegsPortxREG_FILE_03xx0x, fromRegsPortxREG_FILE_04xx31x, 
      fromRegsPortxREG_FILE_04xx30x, fromRegsPortxREG_FILE_04xx29x, 
      fromRegsPortxREG_FILE_04xx28x, fromRegsPortxREG_FILE_04xx27x, 
      fromRegsPortxREG_FILE_04xx26x, fromRegsPortxREG_FILE_04xx25x, 
      fromRegsPortxREG_FILE_04xx24x, fromRegsPortxREG_FILE_04xx23x, 
      fromRegsPortxREG_FILE_04xx22x, fromRegsPortxREG_FILE_04xx21x, 
      fromRegsPortxREG_FILE_04xx20x, fromRegsPortxREG_FILE_04xx19x, 
      fromRegsPortxREG_FILE_04xx18x, fromRegsPortxREG_FILE_04xx17x, 
      fromRegsPortxREG_FILE_04xx16x, fromRegsPortxREG_FILE_04xx15x, 
      fromRegsPortxREG_FILE_04xx14x, fromRegsPortxREG_FILE_04xx13x, 
      fromRegsPortxREG_FILE_04xx12x, fromRegsPortxREG_FILE_04xx11x, 
      fromRegsPortxREG_FILE_04xx10x, fromRegsPortxREG_FILE_04xx9x, 
      fromRegsPortxREG_FILE_04xx8x, fromRegsPortxREG_FILE_04xx7x, 
      fromRegsPortxREG_FILE_04xx6x, fromRegsPortxREG_FILE_04xx5x, 
      fromRegsPortxREG_FILE_04xx4x, fromRegsPortxREG_FILE_04xx3x, 
      fromRegsPortxREG_FILE_04xx2x, fromRegsPortxREG_FILE_04xx1x, 
      fromRegsPortxREG_FILE_04xx0x, fromRegsPortxREG_FILE_05xx31x, 
      fromRegsPortxREG_FILE_05xx30x, fromRegsPortxREG_FILE_05xx29x, 
      fromRegsPortxREG_FILE_05xx28x, fromRegsPortxREG_FILE_05xx27x, 
      fromRegsPortxREG_FILE_05xx26x, fromRegsPortxREG_FILE_05xx25x, 
      fromRegsPortxREG_FILE_05xx24x, fromRegsPortxREG_FILE_05xx23x, 
      fromRegsPortxREG_FILE_05xx22x, fromRegsPortxREG_FILE_05xx21x, 
      fromRegsPortxREG_FILE_05xx20x, fromRegsPortxREG_FILE_05xx19x, 
      fromRegsPortxREG_FILE_05xx18x, fromRegsPortxREG_FILE_05xx17x, 
      fromRegsPortxREG_FILE_05xx16x, fromRegsPortxREG_FILE_05xx15x, 
      fromRegsPortxREG_FILE_05xx14x, fromRegsPortxREG_FILE_05xx13x, 
      fromRegsPortxREG_FILE_05xx12x, fromRegsPortxREG_FILE_05xx11x, 
      fromRegsPortxREG_FILE_05xx10x, fromRegsPortxREG_FILE_05xx9x, 
      fromRegsPortxREG_FILE_05xx8x, fromRegsPortxREG_FILE_05xx7x, 
      fromRegsPortxREG_FILE_05xx6x, fromRegsPortxREG_FILE_05xx5x, 
      fromRegsPortxREG_FILE_05xx4x, fromRegsPortxREG_FILE_05xx3x, 
      fromRegsPortxREG_FILE_05xx2x, fromRegsPortxREG_FILE_05xx1x, 
      fromRegsPortxREG_FILE_05xx0x, fromRegsPortxREG_FILE_06xx31x, 
      fromRegsPortxREG_FILE_06xx30x, fromRegsPortxREG_FILE_06xx29x, 
      fromRegsPortxREG_FILE_06xx28x, fromRegsPortxREG_FILE_06xx27x, 
      fromRegsPortxREG_FILE_06xx26x, fromRegsPortxREG_FILE_06xx25x, 
      fromRegsPortxREG_FILE_06xx24x, fromRegsPortxREG_FILE_06xx23x, 
      fromRegsPortxREG_FILE_06xx22x, fromRegsPortxREG_FILE_06xx21x, 
      fromRegsPortxREG_FILE_06xx20x, fromRegsPortxREG_FILE_06xx19x, 
      fromRegsPortxREG_FILE_06xx18x, fromRegsPortxREG_FILE_06xx17x, 
      fromRegsPortxREG_FILE_06xx16x, fromRegsPortxREG_FILE_06xx15x, 
      fromRegsPortxREG_FILE_06xx14x, fromRegsPortxREG_FILE_06xx13x, 
      fromRegsPortxREG_FILE_06xx12x, fromRegsPortxREG_FILE_06xx11x, 
      fromRegsPortxREG_FILE_06xx10x, fromRegsPortxREG_FILE_06xx9x, 
      fromRegsPortxREG_FILE_06xx8x, fromRegsPortxREG_FILE_06xx7x, 
      fromRegsPortxREG_FILE_06xx6x, fromRegsPortxREG_FILE_06xx5x, 
      fromRegsPortxREG_FILE_06xx4x, fromRegsPortxREG_FILE_06xx3x, 
      fromRegsPortxREG_FILE_06xx2x, fromRegsPortxREG_FILE_06xx1x, 
      fromRegsPortxREG_FILE_06xx0x, fromRegsPortxREG_FILE_07xx31x, 
      fromRegsPortxREG_FILE_07xx30x, fromRegsPortxREG_FILE_07xx29x, 
      fromRegsPortxREG_FILE_07xx28x, fromRegsPortxREG_FILE_07xx27x, 
      fromRegsPortxREG_FILE_07xx26x, fromRegsPortxREG_FILE_07xx25x, 
      fromRegsPortxREG_FILE_07xx24x, fromRegsPortxREG_FILE_07xx23x, 
      fromRegsPortxREG_FILE_07xx22x, fromRegsPortxREG_FILE_07xx21x, 
      fromRegsPortxREG_FILE_07xx20x, fromRegsPortxREG_FILE_07xx19x, 
      fromRegsPortxREG_FILE_07xx18x, fromRegsPortxREG_FILE_07xx17x, 
      fromRegsPortxREG_FILE_07xx16x, fromRegsPortxREG_FILE_07xx15x, 
      fromRegsPortxREG_FILE_07xx14x, fromRegsPortxREG_FILE_07xx13x, 
      fromRegsPortxREG_FILE_07xx12x, fromRegsPortxREG_FILE_07xx11x, 
      fromRegsPortxREG_FILE_07xx10x, fromRegsPortxREG_FILE_07xx9x, 
      fromRegsPortxREG_FILE_07xx8x, fromRegsPortxREG_FILE_07xx7x, 
      fromRegsPortxREG_FILE_07xx6x, fromRegsPortxREG_FILE_07xx5x, 
      fromRegsPortxREG_FILE_07xx4x, fromRegsPortxREG_FILE_07xx3x, 
      fromRegsPortxREG_FILE_07xx2x, fromRegsPortxREG_FILE_07xx1x, 
      fromRegsPortxREG_FILE_07xx0x, fromRegsPortxREG_FILE_08xx31x, 
      fromRegsPortxREG_FILE_08xx30x, fromRegsPortxREG_FILE_08xx29x, 
      fromRegsPortxREG_FILE_08xx28x, fromRegsPortxREG_FILE_08xx27x, 
      fromRegsPortxREG_FILE_08xx26x, fromRegsPortxREG_FILE_08xx25x, 
      fromRegsPortxREG_FILE_08xx24x, fromRegsPortxREG_FILE_08xx23x, 
      fromRegsPortxREG_FILE_08xx22x, fromRegsPortxREG_FILE_08xx21x, 
      fromRegsPortxREG_FILE_08xx20x, fromRegsPortxREG_FILE_08xx19x, 
      fromRegsPortxREG_FILE_08xx18x, fromRegsPortxREG_FILE_08xx17x, 
      fromRegsPortxREG_FILE_08xx16x, fromRegsPortxREG_FILE_08xx15x, 
      fromRegsPortxREG_FILE_08xx14x, fromRegsPortxREG_FILE_08xx13x, 
      fromRegsPortxREG_FILE_08xx12x, fromRegsPortxREG_FILE_08xx11x, 
      fromRegsPortxREG_FILE_08xx10x, fromRegsPortxREG_FILE_08xx9x, 
      fromRegsPortxREG_FILE_08xx8x, fromRegsPortxREG_FILE_08xx7x, 
      fromRegsPortxREG_FILE_08xx6x, fromRegsPortxREG_FILE_08xx5x, 
      fromRegsPortxREG_FILE_08xx4x, fromRegsPortxREG_FILE_08xx3x, 
      fromRegsPortxREG_FILE_08xx2x, fromRegsPortxREG_FILE_08xx1x, 
      fromRegsPortxREG_FILE_08xx0x, fromRegsPortxREG_FILE_09xx31x, 
      fromRegsPortxREG_FILE_09xx30x, fromRegsPortxREG_FILE_09xx29x, 
      fromRegsPortxREG_FILE_09xx28x, fromRegsPortxREG_FILE_09xx27x, 
      fromRegsPortxREG_FILE_09xx26x, fromRegsPortxREG_FILE_09xx25x, 
      fromRegsPortxREG_FILE_09xx24x, fromRegsPortxREG_FILE_09xx23x, 
      fromRegsPortxREG_FILE_09xx22x, fromRegsPortxREG_FILE_09xx21x, 
      fromRegsPortxREG_FILE_09xx20x, fromRegsPortxREG_FILE_09xx19x, 
      fromRegsPortxREG_FILE_09xx18x, fromRegsPortxREG_FILE_09xx17x, 
      fromRegsPortxREG_FILE_09xx16x, fromRegsPortxREG_FILE_09xx15x, 
      fromRegsPortxREG_FILE_09xx14x, fromRegsPortxREG_FILE_09xx13x, 
      fromRegsPortxREG_FILE_09xx12x, fromRegsPortxREG_FILE_09xx11x, 
      fromRegsPortxREG_FILE_09xx10x, fromRegsPortxREG_FILE_09xx9x, 
      fromRegsPortxREG_FILE_09xx8x, fromRegsPortxREG_FILE_09xx7x, 
      fromRegsPortxREG_FILE_09xx6x, fromRegsPortxREG_FILE_09xx5x, 
      fromRegsPortxREG_FILE_09xx4x, fromRegsPortxREG_FILE_09xx3x, 
      fromRegsPortxREG_FILE_09xx2x, fromRegsPortxREG_FILE_09xx1x, 
      fromRegsPortxREG_FILE_09xx0x, fromRegsPortxREG_FILE_10xx31x, 
      fromRegsPortxREG_FILE_10xx30x, fromRegsPortxREG_FILE_10xx29x, 
      fromRegsPortxREG_FILE_10xx28x, fromRegsPortxREG_FILE_10xx27x, 
      fromRegsPortxREG_FILE_10xx26x, fromRegsPortxREG_FILE_10xx25x, 
      fromRegsPortxREG_FILE_10xx24x, fromRegsPortxREG_FILE_10xx23x, 
      fromRegsPortxREG_FILE_10xx22x, fromRegsPortxREG_FILE_10xx21x, 
      fromRegsPortxREG_FILE_10xx20x, fromRegsPortxREG_FILE_10xx19x, 
      fromRegsPortxREG_FILE_10xx18x, fromRegsPortxREG_FILE_10xx17x, 
      fromRegsPortxREG_FILE_10xx16x, fromRegsPortxREG_FILE_10xx15x, 
      fromRegsPortxREG_FILE_10xx14x, fromRegsPortxREG_FILE_10xx13x, 
      fromRegsPortxREG_FILE_10xx12x, fromRegsPortxREG_FILE_10xx11x, 
      fromRegsPortxREG_FILE_10xx10x, fromRegsPortxREG_FILE_10xx9x, 
      fromRegsPortxREG_FILE_10xx8x, fromRegsPortxREG_FILE_10xx7x, 
      fromRegsPortxREG_FILE_10xx6x, fromRegsPortxREG_FILE_10xx5x, 
      fromRegsPortxREG_FILE_10xx4x, fromRegsPortxREG_FILE_10xx3x, 
      fromRegsPortxREG_FILE_10xx2x, fromRegsPortxREG_FILE_10xx1x, 
      fromRegsPortxREG_FILE_10xx0x, fromRegsPortxREG_FILE_11xx31x, 
      fromRegsPortxREG_FILE_11xx30x, fromRegsPortxREG_FILE_11xx29x, 
      fromRegsPortxREG_FILE_11xx28x, fromRegsPortxREG_FILE_11xx27x, 
      fromRegsPortxREG_FILE_11xx26x, fromRegsPortxREG_FILE_11xx25x, 
      fromRegsPortxREG_FILE_11xx24x, fromRegsPortxREG_FILE_11xx23x, 
      fromRegsPortxREG_FILE_11xx22x, fromRegsPortxREG_FILE_11xx21x, 
      fromRegsPortxREG_FILE_11xx20x, fromRegsPortxREG_FILE_11xx19x, 
      fromRegsPortxREG_FILE_11xx18x, fromRegsPortxREG_FILE_11xx17x, 
      fromRegsPortxREG_FILE_11xx16x, fromRegsPortxREG_FILE_11xx15x, 
      fromRegsPortxREG_FILE_11xx14x, fromRegsPortxREG_FILE_11xx13x, 
      fromRegsPortxREG_FILE_11xx12x, fromRegsPortxREG_FILE_11xx11x, 
      fromRegsPortxREG_FILE_11xx10x, fromRegsPortxREG_FILE_11xx9x, 
      fromRegsPortxREG_FILE_11xx8x, fromRegsPortxREG_FILE_11xx7x, 
      fromRegsPortxREG_FILE_11xx6x, fromRegsPortxREG_FILE_11xx5x, 
      fromRegsPortxREG_FILE_11xx4x, fromRegsPortxREG_FILE_11xx3x, 
      fromRegsPortxREG_FILE_11xx2x, fromRegsPortxREG_FILE_11xx1x, 
      fromRegsPortxREG_FILE_11xx0x, fromRegsPortxREG_FILE_12xx31x, 
      fromRegsPortxREG_FILE_12xx30x, fromRegsPortxREG_FILE_12xx29x, 
      fromRegsPortxREG_FILE_12xx28x, fromRegsPortxREG_FILE_12xx27x, 
      fromRegsPortxREG_FILE_12xx26x, fromRegsPortxREG_FILE_12xx25x, 
      fromRegsPortxREG_FILE_12xx24x, fromRegsPortxREG_FILE_12xx23x, 
      fromRegsPortxREG_FILE_12xx22x, fromRegsPortxREG_FILE_12xx21x, 
      fromRegsPortxREG_FILE_12xx20x, fromRegsPortxREG_FILE_12xx19x, 
      fromRegsPortxREG_FILE_12xx18x, fromRegsPortxREG_FILE_12xx17x, 
      fromRegsPortxREG_FILE_12xx16x, fromRegsPortxREG_FILE_12xx15x, 
      fromRegsPortxREG_FILE_12xx14x, fromRegsPortxREG_FILE_12xx13x, 
      fromRegsPortxREG_FILE_12xx12x, fromRegsPortxREG_FILE_12xx11x, 
      fromRegsPortxREG_FILE_12xx10x, fromRegsPortxREG_FILE_12xx9x, 
      fromRegsPortxREG_FILE_12xx8x, fromRegsPortxREG_FILE_12xx7x, 
      fromRegsPortxREG_FILE_12xx6x, fromRegsPortxREG_FILE_12xx5x, 
      fromRegsPortxREG_FILE_12xx4x, fromRegsPortxREG_FILE_12xx3x, 
      fromRegsPortxREG_FILE_12xx2x, fromRegsPortxREG_FILE_12xx1x, 
      fromRegsPortxREG_FILE_12xx0x, fromRegsPortxREG_FILE_13xx31x, 
      fromRegsPortxREG_FILE_13xx30x, fromRegsPortxREG_FILE_13xx29x, 
      fromRegsPortxREG_FILE_13xx28x, fromRegsPortxREG_FILE_13xx27x, 
      fromRegsPortxREG_FILE_13xx26x, fromRegsPortxREG_FILE_13xx25x, 
      fromRegsPortxREG_FILE_13xx24x, fromRegsPortxREG_FILE_13xx23x, 
      fromRegsPortxREG_FILE_13xx22x, fromRegsPortxREG_FILE_13xx21x, 
      fromRegsPortxREG_FILE_13xx20x, fromRegsPortxREG_FILE_13xx19x, 
      fromRegsPortxREG_FILE_13xx18x, fromRegsPortxREG_FILE_13xx17x, 
      fromRegsPortxREG_FILE_13xx16x, fromRegsPortxREG_FILE_13xx15x, 
      fromRegsPortxREG_FILE_13xx14x, fromRegsPortxREG_FILE_13xx13x, 
      fromRegsPortxREG_FILE_13xx12x, fromRegsPortxREG_FILE_13xx11x, 
      fromRegsPortxREG_FILE_13xx10x, fromRegsPortxREG_FILE_13xx9x, 
      fromRegsPortxREG_FILE_13xx8x, fromRegsPortxREG_FILE_13xx7x, 
      fromRegsPortxREG_FILE_13xx6x, fromRegsPortxREG_FILE_13xx5x, 
      fromRegsPortxREG_FILE_13xx4x, fromRegsPortxREG_FILE_13xx3x, 
      fromRegsPortxREG_FILE_13xx2x, fromRegsPortxREG_FILE_13xx1x, 
      fromRegsPortxREG_FILE_13xx0x, fromRegsPortxREG_FILE_14xx31x, 
      fromRegsPortxREG_FILE_14xx30x, fromRegsPortxREG_FILE_14xx29x, 
      fromRegsPortxREG_FILE_14xx28x, fromRegsPortxREG_FILE_14xx27x, 
      fromRegsPortxREG_FILE_14xx26x, fromRegsPortxREG_FILE_14xx25x, 
      fromRegsPortxREG_FILE_14xx24x, fromRegsPortxREG_FILE_14xx23x, 
      fromRegsPortxREG_FILE_14xx22x, fromRegsPortxREG_FILE_14xx21x, 
      fromRegsPortxREG_FILE_14xx20x, fromRegsPortxREG_FILE_14xx19x, 
      fromRegsPortxREG_FILE_14xx18x, fromRegsPortxREG_FILE_14xx17x, 
      fromRegsPortxREG_FILE_14xx16x, fromRegsPortxREG_FILE_14xx15x, 
      fromRegsPortxREG_FILE_14xx14x, fromRegsPortxREG_FILE_14xx13x, 
      fromRegsPortxREG_FILE_14xx12x, fromRegsPortxREG_FILE_14xx11x, 
      fromRegsPortxREG_FILE_14xx10x, fromRegsPortxREG_FILE_14xx9x, 
      fromRegsPortxREG_FILE_14xx8x, fromRegsPortxREG_FILE_14xx7x, 
      fromRegsPortxREG_FILE_14xx6x, fromRegsPortxREG_FILE_14xx5x, 
      fromRegsPortxREG_FILE_14xx4x, fromRegsPortxREG_FILE_14xx3x, 
      fromRegsPortxREG_FILE_14xx2x, fromRegsPortxREG_FILE_14xx1x, 
      fromRegsPortxREG_FILE_14xx0x, fromRegsPortxREG_FILE_15xx31x, 
      fromRegsPortxREG_FILE_15xx30x, fromRegsPortxREG_FILE_15xx29x, 
      fromRegsPortxREG_FILE_15xx28x, fromRegsPortxREG_FILE_15xx27x, 
      fromRegsPortxREG_FILE_15xx26x, fromRegsPortxREG_FILE_15xx25x, 
      fromRegsPortxREG_FILE_15xx24x, fromRegsPortxREG_FILE_15xx23x, 
      fromRegsPortxREG_FILE_15xx22x, fromRegsPortxREG_FILE_15xx21x, 
      fromRegsPortxREG_FILE_15xx20x, fromRegsPortxREG_FILE_15xx19x, 
      fromRegsPortxREG_FILE_15xx18x, fromRegsPortxREG_FILE_15xx17x, 
      fromRegsPortxREG_FILE_15xx16x, fromRegsPortxREG_FILE_15xx15x, 
      fromRegsPortxREG_FILE_15xx14x, fromRegsPortxREG_FILE_15xx13x, 
      fromRegsPortxREG_FILE_15xx12x, fromRegsPortxREG_FILE_15xx11x, 
      fromRegsPortxREG_FILE_15xx10x, fromRegsPortxREG_FILE_15xx9x, 
      fromRegsPortxREG_FILE_15xx8x, fromRegsPortxREG_FILE_15xx7x, 
      fromRegsPortxREG_FILE_15xx6x, fromRegsPortxREG_FILE_15xx5x, 
      fromRegsPortxREG_FILE_15xx4x, fromRegsPortxREG_FILE_15xx3x, 
      fromRegsPortxREG_FILE_15xx2x, fromRegsPortxREG_FILE_15xx1x, 
      fromRegsPortxREG_FILE_15xx0x, fromRegsPortxREG_FILE_16xx31x, 
      fromRegsPortxREG_FILE_16xx30x, fromRegsPortxREG_FILE_16xx29x, 
      fromRegsPortxREG_FILE_16xx28x, fromRegsPortxREG_FILE_16xx27x, 
      fromRegsPortxREG_FILE_16xx26x, fromRegsPortxREG_FILE_16xx25x, 
      fromRegsPortxREG_FILE_16xx24x, fromRegsPortxREG_FILE_16xx23x, 
      fromRegsPortxREG_FILE_16xx22x, fromRegsPortxREG_FILE_16xx21x, 
      fromRegsPortxREG_FILE_16xx20x, fromRegsPortxREG_FILE_16xx19x, 
      fromRegsPortxREG_FILE_16xx18x, fromRegsPortxREG_FILE_16xx17x, 
      fromRegsPortxREG_FILE_16xx16x, fromRegsPortxREG_FILE_16xx15x, 
      fromRegsPortxREG_FILE_16xx14x, fromRegsPortxREG_FILE_16xx13x, 
      fromRegsPortxREG_FILE_16xx12x, fromRegsPortxREG_FILE_16xx11x, 
      fromRegsPortxREG_FILE_16xx10x, fromRegsPortxREG_FILE_16xx9x, 
      fromRegsPortxREG_FILE_16xx8x, fromRegsPortxREG_FILE_16xx7x, 
      fromRegsPortxREG_FILE_16xx6x, fromRegsPortxREG_FILE_16xx5x, 
      fromRegsPortxREG_FILE_16xx4x, fromRegsPortxREG_FILE_16xx3x, 
      fromRegsPortxREG_FILE_16xx2x, fromRegsPortxREG_FILE_16xx1x, 
      fromRegsPortxREG_FILE_16xx0x, fromRegsPortxREG_FILE_17xx31x, 
      fromRegsPortxREG_FILE_17xx30x, fromRegsPortxREG_FILE_17xx29x, 
      fromRegsPortxREG_FILE_17xx28x, fromRegsPortxREG_FILE_17xx27x, 
      fromRegsPortxREG_FILE_17xx26x, fromRegsPortxREG_FILE_17xx25x, 
      fromRegsPortxREG_FILE_17xx24x, fromRegsPortxREG_FILE_17xx23x, 
      fromRegsPortxREG_FILE_17xx22x, fromRegsPortxREG_FILE_17xx21x, 
      fromRegsPortxREG_FILE_17xx20x, fromRegsPortxREG_FILE_17xx19x, 
      fromRegsPortxREG_FILE_17xx18x, fromRegsPortxREG_FILE_17xx17x, 
      fromRegsPortxREG_FILE_17xx16x, fromRegsPortxREG_FILE_17xx15x, 
      fromRegsPortxREG_FILE_17xx14x, fromRegsPortxREG_FILE_17xx13x, 
      fromRegsPortxREG_FILE_17xx12x, fromRegsPortxREG_FILE_17xx11x, 
      fromRegsPortxREG_FILE_17xx10x, fromRegsPortxREG_FILE_17xx9x, 
      fromRegsPortxREG_FILE_17xx8x, fromRegsPortxREG_FILE_17xx7x, 
      fromRegsPortxREG_FILE_17xx6x, fromRegsPortxREG_FILE_17xx5x, 
      fromRegsPortxREG_FILE_17xx4x, fromRegsPortxREG_FILE_17xx3x, 
      fromRegsPortxREG_FILE_17xx2x, fromRegsPortxREG_FILE_17xx1x, 
      fromRegsPortxREG_FILE_17xx0x, fromRegsPortxREG_FILE_18xx31x, 
      fromRegsPortxREG_FILE_18xx30x, fromRegsPortxREG_FILE_18xx29x, 
      fromRegsPortxREG_FILE_18xx28x, fromRegsPortxREG_FILE_18xx27x, 
      fromRegsPortxREG_FILE_18xx26x, fromRegsPortxREG_FILE_18xx25x, 
      fromRegsPortxREG_FILE_18xx24x, fromRegsPortxREG_FILE_18xx23x, 
      fromRegsPortxREG_FILE_18xx22x, fromRegsPortxREG_FILE_18xx21x, 
      fromRegsPortxREG_FILE_18xx20x, fromRegsPortxREG_FILE_18xx19x, 
      fromRegsPortxREG_FILE_18xx18x, fromRegsPortxREG_FILE_18xx17x, 
      fromRegsPortxREG_FILE_18xx16x, fromRegsPortxREG_FILE_18xx15x, 
      fromRegsPortxREG_FILE_18xx14x, fromRegsPortxREG_FILE_18xx13x, 
      fromRegsPortxREG_FILE_18xx12x, fromRegsPortxREG_FILE_18xx11x, 
      fromRegsPortxREG_FILE_18xx10x, fromRegsPortxREG_FILE_18xx9x, 
      fromRegsPortxREG_FILE_18xx8x, fromRegsPortxREG_FILE_18xx7x, 
      fromRegsPortxREG_FILE_18xx6x, fromRegsPortxREG_FILE_18xx5x, 
      fromRegsPortxREG_FILE_18xx4x, fromRegsPortxREG_FILE_18xx3x, 
      fromRegsPortxREG_FILE_18xx2x, fromRegsPortxREG_FILE_18xx1x, 
      fromRegsPortxREG_FILE_18xx0x, fromRegsPortxREG_FILE_19xx31x, 
      fromRegsPortxREG_FILE_19xx30x, fromRegsPortxREG_FILE_19xx29x, 
      fromRegsPortxREG_FILE_19xx28x, fromRegsPortxREG_FILE_19xx27x, 
      fromRegsPortxREG_FILE_19xx26x, fromRegsPortxREG_FILE_19xx25x, 
      fromRegsPortxREG_FILE_19xx24x, fromRegsPortxREG_FILE_19xx23x, 
      fromRegsPortxREG_FILE_19xx22x, fromRegsPortxREG_FILE_19xx21x, 
      fromRegsPortxREG_FILE_19xx20x, fromRegsPortxREG_FILE_19xx19x, 
      fromRegsPortxREG_FILE_19xx18x, fromRegsPortxREG_FILE_19xx17x, 
      fromRegsPortxREG_FILE_19xx16x, fromRegsPortxREG_FILE_19xx15x, 
      fromRegsPortxREG_FILE_19xx14x, fromRegsPortxREG_FILE_19xx13x, 
      fromRegsPortxREG_FILE_19xx12x, fromRegsPortxREG_FILE_19xx11x, 
      fromRegsPortxREG_FILE_19xx10x, fromRegsPortxREG_FILE_19xx9x, 
      fromRegsPortxREG_FILE_19xx8x, fromRegsPortxREG_FILE_19xx7x, 
      fromRegsPortxREG_FILE_19xx6x, fromRegsPortxREG_FILE_19xx5x, 
      fromRegsPortxREG_FILE_19xx4x, fromRegsPortxREG_FILE_19xx3x, 
      fromRegsPortxREG_FILE_19xx2x, fromRegsPortxREG_FILE_19xx1x, 
      fromRegsPortxREG_FILE_19xx0x, fromRegsPortxREG_FILE_20xx31x, 
      fromRegsPortxREG_FILE_20xx30x, fromRegsPortxREG_FILE_20xx29x, 
      fromRegsPortxREG_FILE_20xx28x, fromRegsPortxREG_FILE_20xx27x, 
      fromRegsPortxREG_FILE_20xx26x, fromRegsPortxREG_FILE_20xx25x, 
      fromRegsPortxREG_FILE_20xx24x, fromRegsPortxREG_FILE_20xx23x, 
      fromRegsPortxREG_FILE_20xx22x, fromRegsPortxREG_FILE_20xx21x, 
      fromRegsPortxREG_FILE_20xx20x, fromRegsPortxREG_FILE_20xx19x, 
      fromRegsPortxREG_FILE_20xx18x, fromRegsPortxREG_FILE_20xx17x, 
      fromRegsPortxREG_FILE_20xx16x, fromRegsPortxREG_FILE_20xx15x, 
      fromRegsPortxREG_FILE_20xx14x, fromRegsPortxREG_FILE_20xx13x, 
      fromRegsPortxREG_FILE_20xx12x, fromRegsPortxREG_FILE_20xx11x, 
      fromRegsPortxREG_FILE_20xx10x, fromRegsPortxREG_FILE_20xx9x, 
      fromRegsPortxREG_FILE_20xx8x, fromRegsPortxREG_FILE_20xx7x, 
      fromRegsPortxREG_FILE_20xx6x, fromRegsPortxREG_FILE_20xx5x, 
      fromRegsPortxREG_FILE_20xx4x, fromRegsPortxREG_FILE_20xx3x, 
      fromRegsPortxREG_FILE_20xx2x, fromRegsPortxREG_FILE_20xx1x, 
      fromRegsPortxREG_FILE_20xx0x, fromRegsPortxREG_FILE_21xx31x, 
      fromRegsPortxREG_FILE_21xx30x, fromRegsPortxREG_FILE_21xx29x, 
      fromRegsPortxREG_FILE_21xx28x, fromRegsPortxREG_FILE_21xx27x, 
      fromRegsPortxREG_FILE_21xx26x, fromRegsPortxREG_FILE_21xx25x, 
      fromRegsPortxREG_FILE_21xx24x, fromRegsPortxREG_FILE_21xx23x, 
      fromRegsPortxREG_FILE_21xx22x, fromRegsPortxREG_FILE_21xx21x, 
      fromRegsPortxREG_FILE_21xx20x, fromRegsPortxREG_FILE_21xx19x, 
      fromRegsPortxREG_FILE_21xx18x, fromRegsPortxREG_FILE_21xx17x, 
      fromRegsPortxREG_FILE_21xx16x, fromRegsPortxREG_FILE_21xx15x, 
      fromRegsPortxREG_FILE_21xx14x, fromRegsPortxREG_FILE_21xx13x, 
      fromRegsPortxREG_FILE_21xx12x, fromRegsPortxREG_FILE_21xx11x, 
      fromRegsPortxREG_FILE_21xx10x, fromRegsPortxREG_FILE_21xx9x, 
      fromRegsPortxREG_FILE_21xx8x, fromRegsPortxREG_FILE_21xx7x, 
      fromRegsPortxREG_FILE_21xx6x, fromRegsPortxREG_FILE_21xx5x, 
      fromRegsPortxREG_FILE_21xx4x, fromRegsPortxREG_FILE_21xx3x, 
      fromRegsPortxREG_FILE_21xx2x, fromRegsPortxREG_FILE_21xx1x, 
      fromRegsPortxREG_FILE_21xx0x, fromRegsPortxREG_FILE_22xx31x, 
      fromRegsPortxREG_FILE_22xx30x, fromRegsPortxREG_FILE_22xx29x, 
      fromRegsPortxREG_FILE_22xx28x, fromRegsPortxREG_FILE_22xx27x, 
      fromRegsPortxREG_FILE_22xx26x, fromRegsPortxREG_FILE_22xx25x, 
      fromRegsPortxREG_FILE_22xx24x, fromRegsPortxREG_FILE_22xx23x, 
      fromRegsPortxREG_FILE_22xx22x, fromRegsPortxREG_FILE_22xx21x, 
      fromRegsPortxREG_FILE_22xx20x, fromRegsPortxREG_FILE_22xx19x, 
      fromRegsPortxREG_FILE_22xx18x, fromRegsPortxREG_FILE_22xx17x, 
      fromRegsPortxREG_FILE_22xx16x, fromRegsPortxREG_FILE_22xx15x, 
      fromRegsPortxREG_FILE_22xx14x, fromRegsPortxREG_FILE_22xx13x, 
      fromRegsPortxREG_FILE_22xx12x, fromRegsPortxREG_FILE_22xx11x, 
      fromRegsPortxREG_FILE_22xx10x, fromRegsPortxREG_FILE_22xx9x, 
      fromRegsPortxREG_FILE_22xx8x, fromRegsPortxREG_FILE_22xx7x, 
      fromRegsPortxREG_FILE_22xx6x, fromRegsPortxREG_FILE_22xx5x, 
      fromRegsPortxREG_FILE_22xx4x, fromRegsPortxREG_FILE_22xx3x, 
      fromRegsPortxREG_FILE_22xx2x, fromRegsPortxREG_FILE_22xx1x, 
      fromRegsPortxREG_FILE_22xx0x, fromRegsPortxREG_FILE_23xx31x, 
      fromRegsPortxREG_FILE_23xx30x, fromRegsPortxREG_FILE_23xx29x, 
      fromRegsPortxREG_FILE_23xx28x, fromRegsPortxREG_FILE_23xx27x, 
      fromRegsPortxREG_FILE_23xx26x, fromRegsPortxREG_FILE_23xx25x, 
      fromRegsPortxREG_FILE_23xx24x, fromRegsPortxREG_FILE_23xx23x, 
      fromRegsPortxREG_FILE_23xx22x, fromRegsPortxREG_FILE_23xx21x, 
      fromRegsPortxREG_FILE_23xx20x, fromRegsPortxREG_FILE_23xx19x, 
      fromRegsPortxREG_FILE_23xx18x, fromRegsPortxREG_FILE_23xx17x, 
      fromRegsPortxREG_FILE_23xx16x, fromRegsPortxREG_FILE_23xx15x, 
      fromRegsPortxREG_FILE_23xx14x, fromRegsPortxREG_FILE_23xx13x, 
      fromRegsPortxREG_FILE_23xx12x, fromRegsPortxREG_FILE_23xx11x, 
      fromRegsPortxREG_FILE_23xx10x, fromRegsPortxREG_FILE_23xx9x, 
      fromRegsPortxREG_FILE_23xx8x, fromRegsPortxREG_FILE_23xx7x, 
      fromRegsPortxREG_FILE_23xx6x, fromRegsPortxREG_FILE_23xx5x, 
      fromRegsPortxREG_FILE_23xx4x, fromRegsPortxREG_FILE_23xx3x, 
      fromRegsPortxREG_FILE_23xx2x, fromRegsPortxREG_FILE_23xx1x, 
      fromRegsPortxREG_FILE_23xx0x, fromRegsPortxREG_FILE_24xx31x, 
      fromRegsPortxREG_FILE_24xx30x, fromRegsPortxREG_FILE_24xx29x, 
      fromRegsPortxREG_FILE_24xx28x, fromRegsPortxREG_FILE_24xx27x, 
      fromRegsPortxREG_FILE_24xx26x, fromRegsPortxREG_FILE_24xx25x, 
      fromRegsPortxREG_FILE_24xx24x, fromRegsPortxREG_FILE_24xx23x, 
      fromRegsPortxREG_FILE_24xx22x, fromRegsPortxREG_FILE_24xx21x, 
      fromRegsPortxREG_FILE_24xx20x, fromRegsPortxREG_FILE_24xx19x, 
      fromRegsPortxREG_FILE_24xx18x, fromRegsPortxREG_FILE_24xx17x, 
      fromRegsPortxREG_FILE_24xx16x, fromRegsPortxREG_FILE_24xx15x, 
      fromRegsPortxREG_FILE_24xx14x, fromRegsPortxREG_FILE_24xx13x, 
      fromRegsPortxREG_FILE_24xx12x, fromRegsPortxREG_FILE_24xx11x, 
      fromRegsPortxREG_FILE_24xx10x, fromRegsPortxREG_FILE_24xx9x, 
      fromRegsPortxREG_FILE_24xx8x, fromRegsPortxREG_FILE_24xx7x, 
      fromRegsPortxREG_FILE_24xx6x, fromRegsPortxREG_FILE_24xx5x, 
      fromRegsPortxREG_FILE_24xx4x, fromRegsPortxREG_FILE_24xx3x, 
      fromRegsPortxREG_FILE_24xx2x, fromRegsPortxREG_FILE_24xx1x, 
      fromRegsPortxREG_FILE_24xx0x, fromRegsPortxREG_FILE_25xx31x, 
      fromRegsPortxREG_FILE_25xx30x, fromRegsPortxREG_FILE_25xx29x, 
      fromRegsPortxREG_FILE_25xx28x, fromRegsPortxREG_FILE_25xx27x, 
      fromRegsPortxREG_FILE_25xx26x, fromRegsPortxREG_FILE_25xx25x, 
      fromRegsPortxREG_FILE_25xx24x, fromRegsPortxREG_FILE_25xx23x, 
      fromRegsPortxREG_FILE_25xx22x, fromRegsPortxREG_FILE_25xx21x, 
      fromRegsPortxREG_FILE_25xx20x, fromRegsPortxREG_FILE_25xx19x, 
      fromRegsPortxREG_FILE_25xx18x, fromRegsPortxREG_FILE_25xx17x, 
      fromRegsPortxREG_FILE_25xx16x, fromRegsPortxREG_FILE_25xx15x, 
      fromRegsPortxREG_FILE_25xx14x, fromRegsPortxREG_FILE_25xx13x, 
      fromRegsPortxREG_FILE_25xx12x, fromRegsPortxREG_FILE_25xx11x, 
      fromRegsPortxREG_FILE_25xx10x, fromRegsPortxREG_FILE_25xx9x, 
      fromRegsPortxREG_FILE_25xx8x, fromRegsPortxREG_FILE_25xx7x, 
      fromRegsPortxREG_FILE_25xx6x, fromRegsPortxREG_FILE_25xx5x, 
      fromRegsPortxREG_FILE_25xx4x, fromRegsPortxREG_FILE_25xx3x, 
      fromRegsPortxREG_FILE_25xx2x, fromRegsPortxREG_FILE_25xx1x, 
      fromRegsPortxREG_FILE_25xx0x, fromRegsPortxREG_FILE_26xx31x, 
      fromRegsPortxREG_FILE_26xx30x, fromRegsPortxREG_FILE_26xx29x, 
      fromRegsPortxREG_FILE_26xx28x, fromRegsPortxREG_FILE_26xx27x, 
      fromRegsPortxREG_FILE_26xx26x, fromRegsPortxREG_FILE_26xx25x, 
      fromRegsPortxREG_FILE_26xx24x, fromRegsPortxREG_FILE_26xx23x, 
      fromRegsPortxREG_FILE_26xx22x, fromRegsPortxREG_FILE_26xx21x, 
      fromRegsPortxREG_FILE_26xx20x, fromRegsPortxREG_FILE_26xx19x, 
      fromRegsPortxREG_FILE_26xx18x, fromRegsPortxREG_FILE_26xx17x, 
      fromRegsPortxREG_FILE_26xx16x, fromRegsPortxREG_FILE_26xx15x, 
      fromRegsPortxREG_FILE_26xx14x, fromRegsPortxREG_FILE_26xx13x, 
      fromRegsPortxREG_FILE_26xx12x, fromRegsPortxREG_FILE_26xx11x, 
      fromRegsPortxREG_FILE_26xx10x, fromRegsPortxREG_FILE_26xx9x, 
      fromRegsPortxREG_FILE_26xx8x, fromRegsPortxREG_FILE_26xx7x, 
      fromRegsPortxREG_FILE_26xx6x, fromRegsPortxREG_FILE_26xx5x, 
      fromRegsPortxREG_FILE_26xx4x, fromRegsPortxREG_FILE_26xx3x, 
      fromRegsPortxREG_FILE_26xx2x, fromRegsPortxREG_FILE_26xx1x, 
      fromRegsPortxREG_FILE_26xx0x, fromRegsPortxREG_FILE_27xx31x, 
      fromRegsPortxREG_FILE_27xx30x, fromRegsPortxREG_FILE_27xx29x, 
      fromRegsPortxREG_FILE_27xx28x, fromRegsPortxREG_FILE_27xx27x, 
      fromRegsPortxREG_FILE_27xx26x, fromRegsPortxREG_FILE_27xx25x, 
      fromRegsPortxREG_FILE_27xx24x, fromRegsPortxREG_FILE_27xx23x, 
      fromRegsPortxREG_FILE_27xx22x, fromRegsPortxREG_FILE_27xx21x, 
      fromRegsPortxREG_FILE_27xx20x, fromRegsPortxREG_FILE_27xx19x, 
      fromRegsPortxREG_FILE_27xx18x, fromRegsPortxREG_FILE_27xx17x, 
      fromRegsPortxREG_FILE_27xx16x, fromRegsPortxREG_FILE_27xx15x, 
      fromRegsPortxREG_FILE_27xx14x, fromRegsPortxREG_FILE_27xx13x, 
      fromRegsPortxREG_FILE_27xx12x, fromRegsPortxREG_FILE_27xx11x, 
      fromRegsPortxREG_FILE_27xx10x, fromRegsPortxREG_FILE_27xx9x, 
      fromRegsPortxREG_FILE_27xx8x, fromRegsPortxREG_FILE_27xx7x, 
      fromRegsPortxREG_FILE_27xx6x, fromRegsPortxREG_FILE_27xx5x, 
      fromRegsPortxREG_FILE_27xx4x, fromRegsPortxREG_FILE_27xx3x, 
      fromRegsPortxREG_FILE_27xx2x, fromRegsPortxREG_FILE_27xx1x, 
      fromRegsPortxREG_FILE_27xx0x, fromRegsPortxREG_FILE_28xx31x, 
      fromRegsPortxREG_FILE_28xx30x, fromRegsPortxREG_FILE_28xx29x, 
      fromRegsPortxREG_FILE_28xx28x, fromRegsPortxREG_FILE_28xx27x, 
      fromRegsPortxREG_FILE_28xx26x, fromRegsPortxREG_FILE_28xx25x, 
      fromRegsPortxREG_FILE_28xx24x, fromRegsPortxREG_FILE_28xx23x, 
      fromRegsPortxREG_FILE_28xx22x, fromRegsPortxREG_FILE_28xx21x, 
      fromRegsPortxREG_FILE_28xx20x, fromRegsPortxREG_FILE_28xx19x, 
      fromRegsPortxREG_FILE_28xx18x, fromRegsPortxREG_FILE_28xx17x, 
      fromRegsPortxREG_FILE_28xx16x, fromRegsPortxREG_FILE_28xx15x, 
      fromRegsPortxREG_FILE_28xx14x, fromRegsPortxREG_FILE_28xx13x, 
      fromRegsPortxREG_FILE_28xx12x, fromRegsPortxREG_FILE_28xx11x, 
      fromRegsPortxREG_FILE_28xx10x, fromRegsPortxREG_FILE_28xx9x, 
      fromRegsPortxREG_FILE_28xx8x, fromRegsPortxREG_FILE_28xx7x, 
      fromRegsPortxREG_FILE_28xx6x, fromRegsPortxREG_FILE_28xx5x, 
      fromRegsPortxREG_FILE_28xx4x, fromRegsPortxREG_FILE_28xx3x, 
      fromRegsPortxREG_FILE_28xx2x, fromRegsPortxREG_FILE_28xx1x, 
      fromRegsPortxREG_FILE_28xx0x, fromRegsPortxREG_FILE_29xx31x, 
      fromRegsPortxREG_FILE_29xx30x, fromRegsPortxREG_FILE_29xx29x, 
      fromRegsPortxREG_FILE_29xx28x, fromRegsPortxREG_FILE_29xx27x, 
      fromRegsPortxREG_FILE_29xx26x, fromRegsPortxREG_FILE_29xx25x, 
      fromRegsPortxREG_FILE_29xx24x, fromRegsPortxREG_FILE_29xx23x, 
      fromRegsPortxREG_FILE_29xx22x, fromRegsPortxREG_FILE_29xx21x, 
      fromRegsPortxREG_FILE_29xx20x, fromRegsPortxREG_FILE_29xx19x, 
      fromRegsPortxREG_FILE_29xx18x, fromRegsPortxREG_FILE_29xx17x, 
      fromRegsPortxREG_FILE_29xx16x, fromRegsPortxREG_FILE_29xx15x, 
      fromRegsPortxREG_FILE_29xx14x, fromRegsPortxREG_FILE_29xx13x, 
      fromRegsPortxREG_FILE_29xx12x, fromRegsPortxREG_FILE_29xx11x, 
      fromRegsPortxREG_FILE_29xx10x, fromRegsPortxREG_FILE_29xx9x, 
      fromRegsPortxREG_FILE_29xx8x, fromRegsPortxREG_FILE_29xx7x, 
      fromRegsPortxREG_FILE_29xx6x, fromRegsPortxREG_FILE_29xx5x, 
      fromRegsPortxREG_FILE_29xx4x, fromRegsPortxREG_FILE_29xx3x, 
      fromRegsPortxREG_FILE_29xx2x, fromRegsPortxREG_FILE_29xx1x, 
      fromRegsPortxREG_FILE_29xx0x, fromRegsPortxREG_FILE_30xx31x, 
      fromRegsPortxREG_FILE_30xx30x, fromRegsPortxREG_FILE_30xx29x, 
      fromRegsPortxREG_FILE_30xx28x, fromRegsPortxREG_FILE_30xx27x, 
      fromRegsPortxREG_FILE_30xx26x, fromRegsPortxREG_FILE_30xx25x, 
      fromRegsPortxREG_FILE_30xx24x, fromRegsPortxREG_FILE_30xx23x, 
      fromRegsPortxREG_FILE_30xx22x, fromRegsPortxREG_FILE_30xx21x, 
      fromRegsPortxREG_FILE_30xx20x, fromRegsPortxREG_FILE_30xx19x, 
      fromRegsPortxREG_FILE_30xx18x, fromRegsPortxREG_FILE_30xx17x, 
      fromRegsPortxREG_FILE_30xx16x, fromRegsPortxREG_FILE_30xx15x, 
      fromRegsPortxREG_FILE_30xx14x, fromRegsPortxREG_FILE_30xx13x, 
      fromRegsPortxREG_FILE_30xx12x, fromRegsPortxREG_FILE_30xx11x, 
      fromRegsPortxREG_FILE_30xx10x, fromRegsPortxREG_FILE_30xx9x, 
      fromRegsPortxREG_FILE_30xx8x, fromRegsPortxREG_FILE_30xx7x, 
      fromRegsPortxREG_FILE_30xx6x, fromRegsPortxREG_FILE_30xx5x, 
      fromRegsPortxREG_FILE_30xx4x, fromRegsPortxREG_FILE_30xx3x, 
      fromRegsPortxREG_FILE_30xx2x, fromRegsPortxREG_FILE_30xx1x, 
      fromRegsPortxREG_FILE_30xx0x, fromRegsPortxREG_FILE_31xx31x, 
      fromRegsPortxREG_FILE_31xx30x, fromRegsPortxREG_FILE_31xx29x, 
      fromRegsPortxREG_FILE_31xx28x, fromRegsPortxREG_FILE_31xx27x, 
      fromRegsPortxREG_FILE_31xx26x, fromRegsPortxREG_FILE_31xx25x, 
      fromRegsPortxREG_FILE_31xx24x, fromRegsPortxREG_FILE_31xx23x, 
      fromRegsPortxREG_FILE_31xx22x, fromRegsPortxREG_FILE_31xx21x, 
      fromRegsPortxREG_FILE_31xx20x, fromRegsPortxREG_FILE_31xx19x, 
      fromRegsPortxREG_FILE_31xx18x, fromRegsPortxREG_FILE_31xx17x, 
      fromRegsPortxREG_FILE_31xx16x, fromRegsPortxREG_FILE_31xx15x, 
      fromRegsPortxREG_FILE_31xx14x, fromRegsPortxREG_FILE_31xx13x, 
      fromRegsPortxREG_FILE_31xx12x, fromRegsPortxREG_FILE_31xx11x, 
      fromRegsPortxREG_FILE_31xx10x, fromRegsPortxREG_FILE_31xx9x, 
      fromRegsPortxREG_FILE_31xx8x, fromRegsPortxREG_FILE_31xx7x, 
      fromRegsPortxREG_FILE_31xx6x, fromRegsPortxREG_FILE_31xx5x, 
      fromRegsPortxREG_FILE_31xx4x, fromRegsPortxREG_FILE_31xx3x, 
      fromRegsPortxREG_FILE_31xx2x, fromRegsPortxREG_FILE_31xx1x, 
      fromRegsPortxREG_FILE_31xx0x, IF_ISAxN10974, IF_ISAxN10973, IF_ISAxN10972
      , IF_ISAxN10971, IF_ISAxN10970, IF_ISAxN10969, IF_ISAxN10968, 
      IF_ISAxN10967, IF_ISAxN10966, IF_ISAxN10965, IF_ISAxN10964, IF_ISAxN10963
      , IF_ISAxN10962, IF_ISAxN10961, IF_ISAxN10960, IF_ISAxN10959, 
      IF_ISAxN10958, IF_ISAxN10957, IF_ISAxN10956, IF_ISAxN10955, IF_ISAxN10954
      , IF_ISAxN10953, IF_ISAxN10952, IF_ISAxN10951, IF_ISAxN10950, 
      IF_ISAxN10949, IF_ISAxN10948, IF_ISAxN10947, IF_ISAxN10946, IF_ISAxN10945
      , IF_ISAxN10944, IF_ISAxN10943, IF_ISAxN10942, IF_ISAxN10941, 
      IF_ISAxN10940, IF_ISAxN10939, IF_ISAxN10938, IF_ISAxN10936, IF_ISAxN10935
      , IF_ISAxN10904, IF_ISAxN10902, IF_ISAxN10869, IF_ISAxN10868, 
      IF_ISAxN10867, IF_ISAxN10866, IF_ISAxN10865, IF_ISAxN10864, IF_ISAxN10863
      , IF_ISAxN10862, IF_ISAxN10861, IF_ISAxN10860, IF_ISAxN10859, 
      IF_ISAxN10858, IF_ISAxN10857, IF_ISAxN10856, IF_ISAxN10855, IF_ISAxN10854
      , IF_ISAxN10853, IF_ISAxN10852, IF_ISAxN10851, IF_ISAxN10850, 
      IF_ISAxN10849, IF_ISAxN10848, IF_ISAxN10847, IF_ISAxN10846, IF_ISAxN10845
      , IF_ISAxN10844, IF_ISAxN10843, IF_ISAxN10842, IF_ISAxN10832, 
      IF_ISAxN10829, IF_ISAxN2460, IF_ISAxN2459, IF_ISAxpcReg_signal_2_port, 
      IF_ISAxpcReg_signal_3_port, IF_ISAxpcReg_signal_4_port, 
      IF_ISAxpcReg_signal_5_port, IF_ISAxpcReg_signal_6_port, 
      IF_ISAxpcReg_signal_7_port, IF_ISAxpcReg_signal_8_port, 
      IF_ISAxpcReg_signal_9_port, IF_ISAxpcReg_signal_10_port, 
      IF_ISAxpcReg_signal_11_port, IF_ISAxpcReg_signal_12_port, 
      IF_ISAxpcReg_signal_13_port, IF_ISAxpcReg_signal_14_port, 
      IF_ISAxpcReg_signal_15_port, IF_ISAxpcReg_signal_16_port, 
      IF_ISAxpcReg_signal_17_port, IF_ISAxpcReg_signal_18_port, 
      IF_ISAxpcReg_signal_19_port, IF_ISAxpcReg_signal_20_port, 
      IF_ISAxpcReg_signal_21_port, IF_ISAxpcReg_signal_22_port, 
      IF_ISAxpcReg_signal_23_port, IF_ISAxpcReg_signal_24_port, 
      IF_ISAxpcReg_signal_25_port, IF_ISAxpcReg_signal_26_port, 
      IF_ISAxpcReg_signal_27_port, IF_ISAxpcReg_signal_28_port, 
      IF_ISAxpcReg_signal_29_port, IF_ISAxpcReg_signal_30_port, 
      IF_ISAxpcReg_signal_31_port, IF_ISAxsection_0_port, IF_ISAxsection_2_port
      , IF_RegsxN721, IF_RegsxN720, IF_RegsxN719, IF_RegsxN718, IF_RegsxN717, 
      IF_RegsxN716, IF_RegsxN715, IF_RegsxN714, IF_RegsxN713, IF_RegsxN712, 
      IF_RegsxN711, IF_RegsxN710, IF_RegsxN709, IF_RegsxN708, IF_RegsxN707, 
      IF_RegsxN706, IF_RegsxN705, IF_RegsxN704, IF_RegsxN703, IF_RegsxN702, 
      IF_RegsxN701, IF_RegsxN700, IF_RegsxN699, IF_RegsxN698, IF_RegsxN697, 
      IF_RegsxN696, IF_RegsxN695, IF_RegsxN694, IF_RegsxN693, IF_RegsxN692, 
      IF_RegsxN691, IF_RegsxN690, IF_RegsxN689, IF_RegsxN688, IF_RegsxN687, 
      IF_RegsxN686, IF_RegsxN685, IF_RegsxN684, IF_RegsxN683, IF_RegsxN682, 
      IF_RegsxN681, IF_RegsxN680, IF_RegsxN679, IF_RegsxN678, IF_RegsxN677, 
      IF_RegsxN676, IF_RegsxN675, IF_RegsxN674, IF_RegsxN673, IF_RegsxN672, 
      IF_RegsxN671, IF_RegsxN670, IF_RegsxN669, IF_RegsxN668, IF_RegsxN667, 
      IF_RegsxN666, IF_RegsxN665, IF_RegsxN664, IF_RegsxN663, IF_RegsxN662, 
      IF_RegsxN661, IF_RegsxN660, IF_RegsxN659, net6523, net6528, net6533, 
      net6538, net6543, net6548, net6553, net6558, net6563, net6568, net6573, 
      net6578, net6583, net6588, net6593, net6598, net6603, net6608, net6613, 
      net6618, net6623, net6628, net6633, net6638, net6643, net6648, net6653, 
      net6658, net6663, net6668, net6673, net6678, net6683, net6688, net6693, 
      net6698, net6703, ashr_25xAx30x, ashr_25xAx29x, ashr_25xAx28x, 
      ashr_25xAx27x, ashr_25xAx26x, ashr_25xAx25x, ashr_25xAx24x, ashr_25xAx23x
      , ashr_25xAx22x, ashr_25xAx21x, ashr_25xAx20x, ashr_25xAx19x, 
      ashr_25xAx18x, ashr_25xAx17x, ashr_25xAx16x, ashr_25xAx15x, ashr_25xAx14x
      , ashr_25xAx13x, ashr_25xAx12x, ashr_25xAx11x, ashr_25xAx10x, 
      ashr_25xAx9x, ashr_25xAx8x, ashr_25xAx7x, ashr_25xAx6x, ashr_25xAx5x, 
      ashr_25xAx4x, ashr_25xAx3x, ashr_25xAx2x, ashr_25xAx1x, ashr_25xAx0x, 
      ashr_25xSHx4x, ashr_25xSHx3x, n3458, add_x_26xBx30x, add_x_26xBx29x, 
      add_x_26xBx28x, add_x_26xBx27x, add_x_26xBx26x, add_x_26xBx25x, 
      add_x_26xBx24x, add_x_26xBx23x, add_x_26xBx22x, add_x_26xBx21x, 
      add_x_26xBx20x, add_x_26xBx19x, add_x_26xBx18x, add_x_26xBx17x, 
      add_x_26xBx16x, add_x_26xBx15x, add_x_26xBx14x, add_x_26xBx13x, 
      add_x_26xBx12x, add_x_26xBx11x, add_x_26xBx10x, add_x_26xBx9x, 
      add_x_26xBx8x, add_x_26xBx7x, add_x_26xBx6x, add_x_26xBx5x, 
      DP_OP_679J1_122_3096xn99, DP_OP_679J1_122_3096xn98, 
      DP_OP_679J1_122_3096xn97, DP_OP_679J1_122_3096xn96, 
      DP_OP_679J1_122_3096xn95, DP_OP_679J1_122_3096xn94, 
      DP_OP_679J1_122_3096xn93, DP_OP_679J1_122_3096xn92, 
      DP_OP_679J1_122_3096xn91, DP_OP_679J1_122_3096xn90, 
      DP_OP_679J1_122_3096xn89, DP_OP_679J1_122_3096xn88, 
      DP_OP_679J1_122_3096xn87, DP_OP_679J1_122_3096xn86, 
      DP_OP_679J1_122_3096xn85, DP_OP_679J1_122_3096xn84, 
      DP_OP_679J1_122_3096xn83, DP_OP_679J1_122_3096xn82, 
      DP_OP_679J1_122_3096xn81, DP_OP_679J1_122_3096xn80, 
      DP_OP_679J1_122_3096xn79, DP_OP_679J1_122_3096xn78, 
      DP_OP_679J1_122_3096xn77, DP_OP_679J1_122_3096xn76, 
      DP_OP_679J1_122_3096xn75, DP_OP_679J1_122_3096xn74, 
      DP_OP_679J1_122_3096xn73, DP_OP_679J1_122_3096xn72, 
      DP_OP_679J1_122_3096xn71, DP_OP_679J1_122_3096xn70, 
      DP_OP_679J1_122_3096xn69, DP_OP_679J1_122_3096xn68, 
      DP_OP_679J1_122_3096xn67, DP_OP_679J1_122_3096xn66, 
      DP_OP_679J1_122_3096xn65, DP_OP_679J1_122_3096xn64, 
      DP_OP_679J1_122_3096xn63, DP_OP_679J1_122_3096xn62, 
      DP_OP_679J1_122_3096xn61, DP_OP_679J1_122_3096xn60, 
      DP_OP_679J1_122_3096xn59, DP_OP_679J1_122_3096xn58, 
      DP_OP_679J1_122_3096xn57, DP_OP_679J1_122_3096xn56, 
      DP_OP_679J1_122_3096xn55, DP_OP_679J1_122_3096xn54, 
      DP_OP_679J1_122_3096xn53, DP_OP_679J1_122_3096xn52, 
      DP_OP_679J1_122_3096xn51, DP_OP_679J1_122_3096xn50, 
      DP_OP_679J1_122_3096xn49, DP_OP_679J1_122_3096xn48, 
      DP_OP_679J1_122_3096xn47, DP_OP_679J1_122_3096xn46, 
      DP_OP_679J1_122_3096xn45, DP_OP_679J1_122_3096xn44, 
      DP_OP_679J1_122_3096xn43, DP_OP_679J1_122_3096xn42, 
      DP_OP_679J1_122_3096xn41, DP_OP_679J1_122_3096xn40, 
      DP_OP_679J1_122_3096xn39, DP_OP_679J1_122_3096xn38, 
      DP_OP_679J1_122_3096xn32, DP_OP_679J1_122_3096xn31, 
      DP_OP_679J1_122_3096xn30, DP_OP_679J1_122_3096xn29, 
      DP_OP_679J1_122_3096xn28, DP_OP_679J1_122_3096xn27, 
      DP_OP_679J1_122_3096xn26, DP_OP_679J1_122_3096xn25, 
      DP_OP_679J1_122_3096xn24, DP_OP_679J1_122_3096xn23, 
      DP_OP_679J1_122_3096xn22, DP_OP_679J1_122_3096xn21, 
      DP_OP_679J1_122_3096xn20, DP_OP_679J1_122_3096xn19, 
      DP_OP_679J1_122_3096xn18, DP_OP_679J1_122_3096xn17, 
      DP_OP_679J1_122_3096xn16, DP_OP_679J1_122_3096xn15, 
      DP_OP_679J1_122_3096xn14, DP_OP_679J1_122_3096xn13, 
      DP_OP_679J1_122_3096xn12, DP_OP_679J1_122_3096xn11, 
      DP_OP_679J1_122_3096xn10, DP_OP_679J1_122_3096xn9, 
      DP_OP_679J1_122_3096xn8, DP_OP_679J1_122_3096xn7, DP_OP_679J1_122_3096xn6
      , DP_OP_679J1_122_3096xn5, DP_OP_679J1_122_3096xn4, 
      DP_OP_679J1_122_3096xn3, DP_OP_679J1_122_3096xn2, 
      DP_OP_719J1_125_1055xn164, DP_OP_719J1_125_1055xn163, 
      DP_OP_719J1_125_1055xn162, DP_OP_719J1_125_1055xn161, 
      DP_OP_719J1_125_1055xn160, DP_OP_719J1_125_1055xn159, 
      DP_OP_719J1_125_1055xn158, DP_OP_719J1_125_1055xn157, 
      DP_OP_719J1_125_1055xn156, DP_OP_719J1_125_1055xn155, 
      DP_OP_719J1_125_1055xn154, DP_OP_719J1_125_1055xn153, 
      DP_OP_719J1_125_1055xn152, DP_OP_719J1_125_1055xn151, 
      DP_OP_719J1_125_1055xn150, DP_OP_719J1_125_1055xn149, 
      DP_OP_719J1_125_1055xn148, DP_OP_719J1_125_1055xn147, 
      DP_OP_719J1_125_1055xn146, DP_OP_719J1_125_1055xn145, 
      DP_OP_719J1_125_1055xn144, DP_OP_719J1_125_1055xn143, 
      DP_OP_719J1_125_1055xn142, DP_OP_719J1_125_1055xn141, 
      DP_OP_719J1_125_1055xn140, DP_OP_719J1_125_1055xn139, 
      DP_OP_719J1_125_1055xn138, DP_OP_719J1_125_1055xn137, 
      DP_OP_719J1_125_1055xn136, DP_OP_719J1_125_1055xn135, 
      DP_OP_719J1_125_1055xn134, DP_OP_719J1_125_1055xn99, 
      DP_OP_719J1_125_1055xn98, DP_OP_719J1_125_1055xn97, 
      DP_OP_719J1_125_1055xn96, DP_OP_719J1_125_1055xn95, 
      DP_OP_719J1_125_1055xn94, DP_OP_719J1_125_1055xn93, 
      DP_OP_719J1_125_1055xn92, DP_OP_719J1_125_1055xn91, 
      DP_OP_719J1_125_1055xn90, DP_OP_719J1_125_1055xn89, 
      DP_OP_719J1_125_1055xn88, DP_OP_719J1_125_1055xn87, 
      DP_OP_719J1_125_1055xn86, DP_OP_719J1_125_1055xn85, 
      DP_OP_719J1_125_1055xn84, DP_OP_719J1_125_1055xn83, 
      DP_OP_719J1_125_1055xn82, DP_OP_719J1_125_1055xn81, 
      DP_OP_719J1_125_1055xn80, DP_OP_719J1_125_1055xn79, 
      DP_OP_719J1_125_1055xn78, DP_OP_719J1_125_1055xn77, 
      DP_OP_719J1_125_1055xn76, DP_OP_719J1_125_1055xn75, 
      DP_OP_719J1_125_1055xn74, DP_OP_719J1_125_1055xn73, 
      DP_OP_719J1_125_1055xn72, DP_OP_719J1_125_1055xn71, 
      DP_OP_719J1_125_1055xn70, DP_OP_719J1_125_1055xn69, 
      DP_OP_719J1_125_1055xn68, DP_OP_719J1_125_1055xn67, 
      DP_OP_719J1_125_1055xn66, DP_OP_719J1_125_1055xn65, 
      DP_OP_719J1_125_1055xn64, DP_OP_719J1_125_1055xn63, 
      DP_OP_719J1_125_1055xn62, DP_OP_719J1_125_1055xn61, 
      DP_OP_719J1_125_1055xn60, DP_OP_719J1_125_1055xn59, 
      DP_OP_719J1_125_1055xn58, DP_OP_719J1_125_1055xn57, 
      DP_OP_719J1_125_1055xn56, DP_OP_719J1_125_1055xn55, 
      DP_OP_719J1_125_1055xn54, DP_OP_719J1_125_1055xn53, 
      DP_OP_719J1_125_1055xn52, DP_OP_719J1_125_1055xn51, 
      DP_OP_719J1_125_1055xn50, DP_OP_719J1_125_1055xn49, 
      DP_OP_719J1_125_1055xn48, DP_OP_719J1_125_1055xn47, 
      DP_OP_719J1_125_1055xn46, DP_OP_719J1_125_1055xn45, 
      DP_OP_719J1_125_1055xn44, DP_OP_719J1_125_1055xn43, 
      DP_OP_719J1_125_1055xn42, DP_OP_719J1_125_1055xn41, 
      DP_OP_719J1_125_1055xn40, DP_OP_719J1_125_1055xn39, 
      DP_OP_719J1_125_1055xn38, DP_OP_719J1_125_1055xn32, 
      DP_OP_719J1_125_1055xn31, DP_OP_719J1_125_1055xn30, 
      DP_OP_719J1_125_1055xn29, DP_OP_719J1_125_1055xn28, 
      DP_OP_719J1_125_1055xn27, DP_OP_719J1_125_1055xn26, 
      DP_OP_719J1_125_1055xn25, DP_OP_719J1_125_1055xn24, 
      DP_OP_719J1_125_1055xn23, DP_OP_719J1_125_1055xn22, 
      DP_OP_719J1_125_1055xn21, DP_OP_719J1_125_1055xn20, 
      DP_OP_719J1_125_1055xn19, DP_OP_719J1_125_1055xn18, 
      DP_OP_719J1_125_1055xn17, DP_OP_719J1_125_1055xn16, 
      DP_OP_719J1_125_1055xn15, DP_OP_719J1_125_1055xn14, 
      DP_OP_719J1_125_1055xn13, DP_OP_719J1_125_1055xn12, 
      DP_OP_719J1_125_1055xn11, DP_OP_719J1_125_1055xn10, 
      DP_OP_719J1_125_1055xn9, DP_OP_719J1_125_1055xn8, DP_OP_719J1_125_1055xn7
      , DP_OP_719J1_125_1055xn6, DP_OP_719J1_125_1055xn5, 
      DP_OP_719J1_125_1055xn4, DP_OP_719J1_125_1055xn3, DP_OP_719J1_125_1055xn2
      , intadd_0xBx0x, intadd_0xCI, intadd_0xSUMx28x, intadd_0xSUMx27x, 
      intadd_0xSUMx26x, intadd_0xSUMx25x, intadd_0xSUMx24x, intadd_0xSUMx23x, 
      intadd_0xSUMx22x, intadd_0xSUMx21x, intadd_0xSUMx20x, intadd_0xSUMx19x, 
      intadd_0xSUMx18x, intadd_0xSUMx17x, intadd_0xSUMx16x, intadd_0xSUMx15x, 
      intadd_0xSUMx14x, intadd_0xSUMx13x, intadd_0xSUMx12x, intadd_0xSUMx11x, 
      intadd_0xSUMx10x, intadd_0xSUMx9x, intadd_0xSUMx8x, intadd_0xSUMx7x, 
      intadd_0xSUMx6x, intadd_0xSUMx5x, intadd_0xSUMx4x, intadd_0xSUMx3x, 
      intadd_0xSUMx2x, intadd_0xSUMx1x, intadd_0xSUMx0x, intadd_0xn29, 
      intadd_0xn28, intadd_0xn27, intadd_0xn26, intadd_0xn25, intadd_0xn24, 
      intadd_0xn23, intadd_0xn22, intadd_0xn21, intadd_0xn20, intadd_0xn19, 
      intadd_0xn18, intadd_0xn17, intadd_0xn16, intadd_0xn15, intadd_0xn14, 
      intadd_0xn13, intadd_0xn12, intadd_0xn11, intadd_0xn10, intadd_0xn9, 
      intadd_0xn8, intadd_0xn7, intadd_0xn6, intadd_0xn5, intadd_0xn4, 
      intadd_0xn3, intadd_0xn2, intadd_0xn1, intadd_1xAx7x, intadd_1xAx6x, 
      intadd_1xAx5x, intadd_1xAx4x, intadd_1xAx3x, intadd_1xAx2x, intadd_1xAx1x
      , intadd_1xAx0x, intadd_1xBx7x, intadd_1xBx6x, intadd_1xBx5x, 
      intadd_1xBx4x, intadd_1xBx3x, intadd_1xBx2x, intadd_1xBx1x, intadd_1xBx0x
      , intadd_1xCI, intadd_1xSUMx7x, intadd_1xSUMx6x, intadd_1xSUMx5x, 
      intadd_1xSUMx4x, intadd_1xSUMx3x, intadd_1xSUMx2x, intadd_1xSUMx1x, 
      intadd_1xSUMx0x, intadd_1xn8, intadd_1xn7, intadd_1xn6, intadd_1xn5, 
      intadd_1xn4, intadd_1xn3, intadd_1xn2, intadd_1xn1, intadd_2xAx3x, 
      intadd_2xAx2x, intadd_2xAx1x, intadd_2xAx0x, intadd_2xBx3x, intadd_2xBx2x
      , intadd_2xBx1x, intadd_2xBx0x, intadd_2xCI, intadd_2xSUMx3x, 
      intadd_2xSUMx2x, intadd_2xSUMx1x, intadd_2xSUMx0x, intadd_2xn4, 
      intadd_2xn3, intadd_2xn2, intadd_2xn1, intadd_3xAx2x, intadd_3xAx1x, 
      intadd_3xAx0x, intadd_3xBx2x, intadd_3xBx1x, intadd_3xBx0x, intadd_3xCI, 
      intadd_3xSUMx2x, intadd_3xSUMx1x, intadd_3xSUMx0x, intadd_3xn3, 
      intadd_3xn2, intadd_3xn1, intadd_4xAx2x, intadd_4xAx1x, intadd_4xAx0x, 
      intadd_4xBx2x, intadd_4xBx1x, intadd_4xBx0x, intadd_4xCI, intadd_4xSUMx2x
      , intadd_4xSUMx1x, intadd_4xSUMx0x, intadd_4xn3, intadd_4xn2, intadd_4xn1
      , n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, 
      n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, 
      n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, 
      n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, 
      n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, 
      n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, 
      n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, 
      n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, 
      n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, 
      n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, 
      n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, 
      n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, 
      n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, 
      n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, 
      n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, 
      n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, 
      n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, 
      n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, 
      n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, 
      n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, 
      n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, 
      n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, 
      n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, 
      n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, 
      n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, 
      n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, 
      n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, 
      n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, 
      n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, 
      n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, 
      n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, 
      n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, 
      n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, 
      n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, 
      n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, 
      n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, 
      n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, 
      n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, 
      n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, 
      n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, 
      n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, 
      n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, 
      n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, 
      n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, 
      n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, 
      n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, 
      n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, 
      n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, 
      n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, 
      n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, 
      n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, 
      n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, 
      n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, 
      n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, 
      n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, 
      n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, 
      n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, 
      n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, 
      n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, 
      n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, 
      n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, 
      n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, 
      n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, 
      n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
      n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, 
      n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, 
      n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, 
      n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, 
      n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, 
      n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, 
      n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, 
      n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, 
      n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, 
      n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, 
      n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, 
      n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, 
      n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, 
      n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, 
      n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, 
      n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, 
      n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, 
      n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, 
      n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, 
      n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, 
      n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, 
      n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, 
      n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, 
      n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, 
      n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, 
      n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, 
      n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, 
      n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, 
      n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, 
      n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, 
      n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, 
      n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, 
      n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, 
      n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, 
      n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, 
      n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, 
      n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, 
      n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, 
      n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, 
      n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, 
      n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, 
      n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, 
      n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, 
      n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, 
      n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, 
      n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, 
      n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, 
      n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, 
      n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, 
      n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, 
      n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, 
      n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, 
      n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, 
      n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, 
      n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, 
      n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, 
      n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, 
      n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, 
      n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, 
      n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, 
      n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, 
      n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, 
      n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, 
      n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, 
      n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, 
      n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, 
      n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, 
      n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, 
      n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, 
      n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, 
      n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, 
      n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, 
      n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, 
      n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, 
      n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, 
      n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, 
      n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, 
      n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, 
      n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, 
      n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, 
      n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, 
      n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, 
      n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, 
      n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, 
      n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, 
      n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, 
      n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, 
      n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, 
      n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, 
      n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, 
      n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, 
      n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, 
      n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, 
      n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, 
      n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, 
      n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, 
      n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, 
      n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, 
      n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, 
      n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, 
      n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, 
      n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, 
      n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, 
      n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, 
      n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, 
      n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, 
      n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, 
      n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, 
      n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, 
      n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, 
      n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, 
      n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, 
      n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, 
      n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, 
      n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, 
      n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, 
      n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, 
      n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, 
      n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, 
      n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, 
      n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, 
      n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, 
      n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, 
      n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, 
      n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, 
      n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, 
      n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, 
      n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, 
      n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, 
      n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, 
      n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, 
      n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, 
      n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, 
      n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, 
      n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, 
      n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, 
      n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, 
      n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, 
      n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, 
      n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, 
      n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, 
      n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, 
      n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, 
      n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, 
      n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, 
      n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, 
      n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, 
      n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, 
      n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, 
      n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, 
      n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, 
      n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, 
      n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, 
      n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, 
      n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, 
      n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, 
      n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, 
      n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, 
      n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, 
      n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, 
      n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, 
      n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, 
      n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, 
      n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, 
      n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, 
      n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, 
      n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, 
      n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, 
      n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, 
      n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, 
      n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, 
      n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, 
      n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, 
      n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, 
      n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, 
      n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, 
      n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, 
      n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, 
      n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, 
      n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, 
      n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, 
      n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, 
      n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, 
      n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, 
      n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, 
      n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, 
      n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, 
      n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, 
      n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, 
      n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, 
      n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, 
      n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, 
      n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, 
      n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, 
      n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, 
      n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, 
      n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, 
      n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, 
      n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, 
      n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, 
      n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, 
      n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, 
      n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, 
      n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, 
      n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, 
      n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, 
      n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, 
      n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, 
      n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, 
      n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, 
      n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, 
      n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, 
      n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, 
      n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, 
      n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, 
      n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, 
      n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, 
      n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, 
      n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, 
      n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, 
      n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, 
      n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, 
      n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, 
      n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, 
      n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, 
      n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, 
      n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, 
      n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, 
      n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, 
      n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, 
      n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, 
      n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, 
      n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, 
      n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, 
      n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, 
      n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, 
      n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, 
      n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, 
      n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, 
      n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, 
      n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, 
      n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, 
      n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, 
      n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, 
      n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, 
      n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, 
      n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, 
      n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, 
      n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, 
      n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, 
      n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, 
      n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, 
      n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, 
      n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, 
      n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, 
      n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, 
      n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, 
      n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, 
      n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, 
      n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, 
      n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, 
      n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, 
      n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, 
      n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, 
      n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, 
      n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, 
      n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, 
      n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, 
      n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, 
      n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, 
      n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, 
      n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, 
      n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, 
      n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, 
      n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, 
      n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, 
      n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, 
      n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, 
      n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, 
      n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, 
      n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, 
      n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, 
      n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, 
      n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, 
      n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, 
      n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, 
      n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, 
      n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, 
      n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, 
      n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, 
      n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, 
      n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, 
      n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, 
      n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, 
      n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, 
      n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, 
      n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, 
      n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, 
      n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, 
      n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, 
      n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, 
      n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, 
      n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, 
      n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, 
      n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, 
      n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, 
      n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, 
      n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, 
      n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, 
      n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, 
      n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, 
      n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, 
      n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, 
      n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, 
      n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, 
      n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, 
      n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, 
      n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, 
      n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, 
      n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, 
      n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, 
      n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, 
      n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, 
      n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, 
      n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, 
      n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, 
      n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, 
      n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, 
      n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, 
      n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, 
      n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, 
      n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, 
      n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, 
      n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, 
      n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, 
      n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, 
      n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, 
      n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, 
      n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, 
      n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, 
      n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, 
      n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, 
      n7618, n7619, n7620, n7621, n7622, n7624, n_1000, n_1001, n_1002, n_1003,
      n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, 
      n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, 
      n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, 
      n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, 
      n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, 
      n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, 
      n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, 
      n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, 
      n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, 
      n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, 
      n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, 
      n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, 
      n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, 
      n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, 
      n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, 
      n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, 
      n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, 
      n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, 
      n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, 
      n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, 
      n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, 
      n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, 
      n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, 
      n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, 
      n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, 
      n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, 
      n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, 
      n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, 
      n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, 
      n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, 
      n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, 
      n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, 
      n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, 
      n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, 
      n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, 
      n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, 
      n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, 
      n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, 
      n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, 
      n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, 
      n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, 
      n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, 
      n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, 
      n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, 
      n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, 
      n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, 
      n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, 
      n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, 
      n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, 
      n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, 
      n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, 
      n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, 
      n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, 
      n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, 
      n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, 
      n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, 
      n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, 
      n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, 
      n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, 
      n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, 
      n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, 
      n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, 
      n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, 
      n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, 
      n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, 
      n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, 
      n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, 
      n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, 
      n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, 
      n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, 
      n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, 
      n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, 
      n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, 
      n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, 
      n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, 
      n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, 
      n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, 
      n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, 
      n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, 
      n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, 
      n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, 
      n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, 
      n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, 
      n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, 
      n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, 
      n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, 
      n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, 
      n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, 
      n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, 
      n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, 
      n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, 
      n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, 
      n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, 
      n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, 
      n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, 
      n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, 
      n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, 
      n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, 
      n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, 
      n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, 
      n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, 
      n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, 
      n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, 
      n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, 
      n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, 
      n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, 
      n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, 
      n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, 
      n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, 
      n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, 
      n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, 
      n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, 
      n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, 
      n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, 
      n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, 
      n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, 
      n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, 
      n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, 
      n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, 
      n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, 
      n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, 
      n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, 
      n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, 
      n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118 : 
      std_logic;

begin
   fromMemoryPort_sync_port <= bool_to_std_logic(fromMemoryPort_sync);
   fromMemoryPort_notify <= std_logic_to_bool(IF_ISAxsection_0_port);
   toMemoryPort_sync_port <= bool_to_std_logic(toMemoryPort_sync);
   toMemoryPort_notify <= std_logic_to_bool(toMemoryPort_notify_port);
   
   IF_ISAxsection_regx2x : DFF_X1 port map( D => n7551, CK => net6523, Q => 
                           IF_ISAxsection_2_port, QN => n7531);
   IF_ISAxsection_regx1x : DFF_X1 port map( D => n7550, CK => net6523, Q => 
                           n_1000, QN => n7534);
   IF_ISAxtoRegsPort_regxDSTxx0x : DFF_X1 port map( D => IF_ISAxN10970, CK => 
                           net6533, Q => toRegsPortxDSTxx0x, QN => n7532);
   IF_ISAxtoRegsPort_regxDSTxx1x : DFF_X1 port map( D => IF_ISAxN10971, CK => 
                           net6533, Q => toRegsPortxDSTxx1x, QN => n7530);
   IF_ISAxtoRegsPort_regxDSTxx2x : DFF_X1 port map( D => IF_ISAxN10972, CK => 
                           net6533, Q => toRegsPortxDSTxx2x, QN => n7533);
   IF_ISAxtoRegsPort_regxDSTxx3x : DFF_X1 port map( D => IF_ISAxN10973, CK => 
                           net6533, Q => toRegsPortxDSTxx3x, QN => n7537);
   IF_ISAxtoRegsPort_regxDSTxx4x : DFF_X1 port map( D => IF_ISAxN10974, CK => 
                           net6533, Q => toRegsPortxDSTxx4x, QN => n7535);
   IF_ISAxsection_regx0x : DFF_X1 port map( D => n7552, CK => net6523, Q => 
                           IF_ISAxsection_0_port, QN => n_1001);
   IF_ISAxpcReg_signal_regx0x : DFF_X1 port map( D => n7548, CK => net6538, Q 
                           => IF_ISAxN2459, QN => n7545);
   IF_ISAxpcReg_signal_regx1x : DFF_X1 port map( D => IF_ISAxN10904, CK => 
                           net6538, Q => IF_ISAxN2460, QN => n7538);
   IF_ISAxpcReg_signal_regx2x : DFF_X1 port map( D => n7582, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_2_port, QN => n7542);
   IF_ISAxpcReg_signal_regx3x : DFF_X1 port map( D => n7581, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_3_port, QN => n_1002);
   IF_ISAxpcReg_signal_regx4x : DFF_X1 port map( D => n7580, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_4_port, QN => n_1003);
   IF_ISAxpcReg_signal_regx5x : DFF_X1 port map( D => n7579, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_5_port, QN => n_1004);
   IF_ISAxpcReg_signal_regx6x : DFF_X1 port map( D => n7578, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_6_port, QN => n7539);
   IF_ISAxpcReg_signal_regx7x : DFF_X1 port map( D => n7577, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_7_port, QN => n_1005);
   IF_ISAxpcReg_signal_regx8x : DFF_X1 port map( D => n7576, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_8_port, QN => n7540);
   IF_ISAxpcReg_signal_regx9x : DFF_X1 port map( D => n7575, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_9_port, QN => n_1006);
   IF_ISAxpcReg_signal_regx10x : DFF_X1 port map( D => n7574, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_10_port, QN => n7541);
   IF_ISAxpcReg_signal_regx11x : DFF_X1 port map( D => n7573, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_11_port, QN => n_1007);
   IF_ISAxpcReg_signal_regx12x : DFF_X1 port map( D => n7572, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_12_port, QN => n7543);
   IF_ISAxpcReg_signal_regx13x : DFF_X1 port map( D => n7571, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_13_port, QN => n_1008);
   IF_ISAxpcReg_signal_regx14x : DFF_X1 port map( D => n7570, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_14_port, QN => n_1009);
   IF_ISAxpcReg_signal_regx15x : DFF_X1 port map( D => n7569, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_15_port, QN => n_1010);
   IF_ISAxpcReg_signal_regx16x : DFF_X1 port map( D => n7568, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_16_port, QN => n_1011);
   IF_ISAxpcReg_signal_regx17x : DFF_X1 port map( D => n7567, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_17_port, QN => n_1012);
   IF_ISAxpcReg_signal_regx18x : DFF_X1 port map( D => n7566, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_18_port, QN => n_1013);
   IF_ISAxpcReg_signal_regx19x : DFF_X1 port map( D => n7565, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_19_port, QN => n_1014);
   IF_ISAxpcReg_signal_regx20x : DFF_X1 port map( D => n7564, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_20_port, QN => n_1015);
   IF_ISAxpcReg_signal_regx21x : DFF_X1 port map( D => n7563, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_21_port, QN => n_1016);
   IF_ISAxpcReg_signal_regx22x : DFF_X1 port map( D => n7562, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_22_port, QN => n_1017);
   IF_ISAxpcReg_signal_regx23x : DFF_X1 port map( D => n7561, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_23_port, QN => n_1018);
   IF_ISAxpcReg_signal_regx24x : DFF_X1 port map( D => n7560, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_24_port, QN => n_1019);
   IF_ISAxpcReg_signal_regx25x : DFF_X1 port map( D => n7559, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_25_port, QN => n_1020);
   IF_ISAxpcReg_signal_regx26x : DFF_X1 port map( D => n7558, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_26_port, QN => n_1021);
   IF_ISAxpcReg_signal_regx27x : DFF_X1 port map( D => n7557, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_27_port, QN => n_1022);
   IF_ISAxpcReg_signal_regx28x : DFF_X1 port map( D => n7556, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_28_port, QN => n_1023);
   IF_ISAxpcReg_signal_regx29x : DFF_X1 port map( D => n7555, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_29_port, QN => n_1024);
   IF_ISAxpcReg_signal_regx30x : DFF_X1 port map( D => n7554, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_30_port, QN => n_1025);
   IF_ISAxpcReg_signal_regx31x : DFF_X1 port map( D => n7553, CK => net6538, Q 
                           => IF_ISAxpcReg_signal_31_port, QN => n7544);
   IF_ISAxtoMemoryPort_regxREQxx0x : DFF_X1 port map( D => n7591, CK => net6543
                           , Q => toMemoryPortxREQxx0x(0), QN => n_1026);
   IF_ISAxtoMemoryPort_regxMASKxx0x : DFF_X1 port map( D => n7590, CK => 
                           net6543, Q => toMemoryPortxMASKxx0x(0), QN => n_1027
                           );
   IF_ISAxtoMemoryPort_regxMASKxx1x : DFF_X1 port map( D => n7589, CK => 
                           net6543, Q => toMemoryPortxMASKxx1x(0), QN => n_1028
                           );
   IF_ISAxtoMemoryPort_regxMASKxx2x : DFF_X1 port map( D => n7588, CK => 
                           net6543, Q => toMemoryPortxMASKxx2x(0), QN => n_1029
                           );
   IF_ISAxtoMemoryPort_regxADDRINxx0x : DFF_X1 port map( D => n7548, CK => 
                           net6548, Q => toMemoryPortxADDRINxx0x(0), QN => 
                           n_1030);
   IF_ISAxtoMemoryPort_regxADDRINxx1x : DFF_X1 port map( D => n7622, CK => 
                           net6548, Q => toMemoryPortxADDRINxx1x(0), QN => 
                           n_1031);
   IF_ISAxtoMemoryPort_regxADDRINxx2x : DFF_X1 port map( D => n7621, CK => 
                           net6548, Q => toMemoryPortxADDRINxx2x(0), QN => 
                           n_1032);
   IF_ISAxtoMemoryPort_regxADDRINxx3x : DFF_X1 port map( D => n7620, CK => 
                           net6548, Q => toMemoryPortxADDRINxx3x(0), QN => 
                           n_1033);
   IF_ISAxtoMemoryPort_regxADDRINxx4x : DFF_X1 port map( D => n7619, CK => 
                           net6548, Q => toMemoryPortxADDRINxx4x(0), QN => 
                           n_1034);
   IF_ISAxtoMemoryPort_regxADDRINxx5x : DFF_X1 port map( D => n7618, CK => 
                           net6548, Q => toMemoryPortxADDRINxx5x(0), QN => 
                           n_1035);
   IF_ISAxtoMemoryPort_regxADDRINxx6x : DFF_X1 port map( D => n7617, CK => 
                           net6548, Q => toMemoryPortxADDRINxx6x(0), QN => 
                           n_1036);
   IF_ISAxtoMemoryPort_regxADDRINxx7x : DFF_X1 port map( D => n7616, CK => 
                           net6548, Q => toMemoryPortxADDRINxx7x(0), QN => 
                           n_1037);
   IF_ISAxtoMemoryPort_regxADDRINxx8x : DFF_X1 port map( D => n7615, CK => 
                           net6548, Q => toMemoryPortxADDRINxx8x(0), QN => 
                           n_1038);
   IF_ISAxtoMemoryPort_regxADDRINxx9x : DFF_X1 port map( D => n7614, CK => 
                           net6548, Q => toMemoryPortxADDRINxx9x(0), QN => 
                           n_1039);
   IF_ISAxtoMemoryPort_regxADDRINxx10x : DFF_X1 port map( D => n7613, CK => 
                           net6548, Q => toMemoryPortxADDRINxx10x(0), QN => 
                           n_1040);
   IF_ISAxtoMemoryPort_regxADDRINxx11x : DFF_X1 port map( D => n7612, CK => 
                           net6548, Q => toMemoryPortxADDRINxx11x(0), QN => 
                           n_1041);
   IF_ISAxtoMemoryPort_regxADDRINxx12x : DFF_X1 port map( D => n7611, CK => 
                           net6548, Q => toMemoryPortxADDRINxx12x(0), QN => 
                           n_1042);
   IF_ISAxtoMemoryPort_regxADDRINxx13x : DFF_X1 port map( D => n7610, CK => 
                           net6548, Q => toMemoryPortxADDRINxx13x(0), QN => 
                           n_1043);
   IF_ISAxtoMemoryPort_regxADDRINxx14x : DFF_X1 port map( D => n7609, CK => 
                           net6548, Q => toMemoryPortxADDRINxx14x(0), QN => 
                           n_1044);
   IF_ISAxtoMemoryPort_regxADDRINxx15x : DFF_X1 port map( D => n7608, CK => 
                           net6548, Q => toMemoryPortxADDRINxx15x(0), QN => 
                           n_1045);
   IF_ISAxtoMemoryPort_regxADDRINxx16x : DFF_X1 port map( D => n7607, CK => 
                           net6548, Q => toMemoryPortxADDRINxx16x(0), QN => 
                           n_1046);
   IF_ISAxtoMemoryPort_regxADDRINxx17x : DFF_X1 port map( D => n7606, CK => 
                           net6548, Q => toMemoryPortxADDRINxx17x(0), QN => 
                           n_1047);
   IF_ISAxtoMemoryPort_regxADDRINxx18x : DFF_X1 port map( D => n7605, CK => 
                           net6548, Q => toMemoryPortxADDRINxx18x(0), QN => 
                           n_1048);
   IF_ISAxtoMemoryPort_regxADDRINxx19x : DFF_X1 port map( D => n7604, CK => 
                           net6548, Q => toMemoryPortxADDRINxx19x(0), QN => 
                           n_1049);
   IF_ISAxtoMemoryPort_regxADDRINxx20x : DFF_X1 port map( D => n7603, CK => 
                           net6548, Q => toMemoryPortxADDRINxx20x(0), QN => 
                           n_1050);
   IF_ISAxtoMemoryPort_regxADDRINxx21x : DFF_X1 port map( D => n7602, CK => 
                           net6548, Q => toMemoryPortxADDRINxx21x(0), QN => 
                           n_1051);
   IF_ISAxtoMemoryPort_regxADDRINxx22x : DFF_X1 port map( D => n7601, CK => 
                           net6548, Q => toMemoryPortxADDRINxx22x(0), QN => 
                           n_1052);
   IF_ISAxtoMemoryPort_regxADDRINxx23x : DFF_X1 port map( D => n7600, CK => 
                           net6548, Q => toMemoryPortxADDRINxx23x(0), QN => 
                           n_1053);
   IF_ISAxtoMemoryPort_regxADDRINxx24x : DFF_X1 port map( D => n7599, CK => 
                           net6548, Q => toMemoryPortxADDRINxx24x(0), QN => 
                           n_1054);
   IF_ISAxtoMemoryPort_regxADDRINxx25x : DFF_X1 port map( D => n7598, CK => 
                           net6548, Q => toMemoryPortxADDRINxx25x(0), QN => 
                           n_1055);
   IF_ISAxtoMemoryPort_regxADDRINxx26x : DFF_X1 port map( D => n7597, CK => 
                           net6548, Q => toMemoryPortxADDRINxx26x(0), QN => 
                           n_1056);
   IF_ISAxtoMemoryPort_regxADDRINxx27x : DFF_X1 port map( D => n7596, CK => 
                           net6548, Q => toMemoryPortxADDRINxx27x(0), QN => 
                           n_1057);
   IF_ISAxtoMemoryPort_regxADDRINxx28x : DFF_X1 port map( D => n7595, CK => 
                           net6548, Q => toMemoryPortxADDRINxx28x(0), QN => 
                           n_1058);
   IF_ISAxtoMemoryPort_regxADDRINxx29x : DFF_X1 port map( D => n7594, CK => 
                           net6548, Q => toMemoryPortxADDRINxx29x(0), QN => 
                           n_1059);
   IF_ISAxtoMemoryPort_regxADDRINxx30x : DFF_X1 port map( D => n7593, CK => 
                           net6548, Q => toMemoryPortxADDRINxx30x(0), QN => 
                           n_1060);
   IF_ISAxtoMemoryPort_regxADDRINxx31x : DFF_X1 port map( D => n7592, CK => 
                           net6548, Q => toMemoryPortxADDRINxx31x(0), QN => 
                           n_1061);
   IF_ISAxtoMemoryPort_notify_reg : DFF_X1 port map( D => n7549, CK => net6523,
                           Q => toMemoryPort_notify_port, QN => n_1062);
   IF_ISAxtoRegsPort_notify_reg : DFF_X1 port map( D => n3458, CK => clk, Q => 
                           toRegsPort_notify, QN => n7536);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx31x, QN => n_1063);
   IF_ISAxtoRegsPort_regxDSTDATAxx31x : DFF_X1 port map( D => IF_ISAxN10968, CK
                           => net6528, Q => toRegsPortxDSTDATAxx31x, QN => 
                           n_1064);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx31x, QN => n_1065);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx31x, QN => n_1066);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx31x, QN => n_1067);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx31x, QN => n_1068);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx31x, QN => n_1069);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx31x, QN => n_1070);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx31x, QN => n_1071);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx31x, QN => n_1072);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx31x, QN => n_1073);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx31x, QN => n_1074);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx31x, QN => n_1075);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx31x, QN => n_1076);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx31x, QN => n_1077);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx31x, QN => n_1078);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx31x, QN => n_1079);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx31x, QN => n_1080);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx31x, QN => n_1081);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx31x, QN => n_1082);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx31x, QN => n_1083);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx31x, QN => n_1084);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx31x, QN => n_1085);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx31x, QN => n_1086);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx31x, QN => n_1087);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx31x, QN => n_1088);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx31x, QN => n_1089);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx31x, QN => n_1090);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx31x, QN => n_1091);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx31x, QN => n_1092);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx31x, QN => n_1093);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx31x, QN => n_1094);
   IF_ISAxtoRegsPort_regxDSTDATAxx15x : DFF_X1 port map( D => IF_ISAxN10952, CK
                           => net6528, Q => toRegsPortxDSTDATAxx15x, QN => 
                           n_1095);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx15x, QN => n_1096);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx15x, QN => n_1097);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx15x, QN => n_1098);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx15x, QN => n_1099);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx15x, QN => n_1100);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx15x, QN => n_1101);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx15x, QN => n_1102);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx15x, QN => n_1103);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx15x, QN => n_1104);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx15x, QN => n_1105);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx15x, QN => n_1106);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx15x, QN => n_1107);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx15x, QN => n_1108);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx15x, QN => n_1109);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx15x, QN => n_1110);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx15x, QN => n_1111);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx15x, QN => n_1112);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx15x, QN => n_1113);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx15x, QN => n_1114);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx15x, QN => n_1115);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx15x, QN => n_1116);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx15x, QN => n_1117);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx15x, QN => n_1118);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx15x, QN => n_1119);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx15x, QN => n_1120);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx15x, QN => n_1121);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx15x, QN => n_1122);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx15x, QN => n_1123);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx15x, QN => n_1124);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx15x, QN => n_1125);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx15x, QN => n_1126);
   IF_ISAxtoRegsPort_regxDSTDATAxx23x : DFF_X1 port map( D => IF_ISAxN10960, CK
                           => net6528, Q => toRegsPortxDSTDATAxx23x, QN => 
                           n_1127);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx23x, QN => n_1128);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx23x, QN => n_1129);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx23x, QN => n_1130);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx23x, QN => n_1131);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx23x, QN => n_1132);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx23x, QN => n_1133);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx23x, QN => n_1134);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx23x, QN => n_1135);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx23x, QN => n_1136);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx23x, QN => n_1137);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx23x, QN => n_1138);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx23x, QN => n_1139);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx23x, QN => n_1140);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx23x, QN => n_1141);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx23x, QN => n_1142);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx23x, QN => n_1143);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx23x, QN => n_1144);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx23x, QN => n_1145);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx23x, QN => n_1146);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx23x, QN => n_1147);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx23x, QN => n_1148);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx23x, QN => n_1149);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx23x, QN => n_1150);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx23x, QN => n_1151);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx23x, QN => n_1152);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx23x, QN => n_1153);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx23x, QN => n_1154);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx23x, QN => n_1155);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx23x, QN => n_1156);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx23x, QN => n_1157);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx23x, QN => n_1158);
   IF_ISAxtoRegsPort_regxDSTDATAxx27x : DFF_X1 port map( D => IF_ISAxN10964, CK
                           => net6528, Q => toRegsPortxDSTDATAxx27x, QN => 
                           n_1159);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx27x, QN => n_1160);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx27x, QN => n_1161);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx27x, QN => n_1162);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx27x, QN => n_1163);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx27x, QN => n_1164);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx27x, QN => n_1165);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx27x, QN => n_1166);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx27x, QN => n_1167);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx27x, QN => n_1168);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx27x, QN => n_1169);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx27x, QN => n_1170);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx27x, QN => n_1171);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx27x, QN => n_1172);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx27x, QN => n_1173);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx27x, QN => n_1174);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx27x, QN => n_1175);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx27x, QN => n_1176);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx27x, QN => n_1177);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx27x, QN => n_1178);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx27x, QN => n_1179);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx27x, QN => n_1180);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx27x, QN => n_1181);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx27x, QN => n_1182);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx27x, QN => n_1183);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx27x, QN => n_1184);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx27x, QN => n_1185);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx27x, QN => n_1186);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx27x, QN => n_1187);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx27x, QN => n_1188);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx27x, QN => n_1189);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx27x, QN => n_1190);
   IF_ISAxtoRegsPort_regxDSTDATAxx29x : DFF_X1 port map( D => IF_ISAxN10966, CK
                           => net6528, Q => toRegsPortxDSTDATAxx29x, QN => 
                           n_1191);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx29x, QN => n_1192);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx29x, QN => n_1193);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx29x, QN => n_1194);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx29x, QN => n_1195);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx29x, QN => n_1196);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx29x, QN => n_1197);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx29x, QN => n_1198);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx29x, QN => n_1199);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx29x, QN => n_1200);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx29x, QN => n_1201);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx29x, QN => n_1202);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx29x, QN => n_1203);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx29x, QN => n_1204);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx29x, QN => n_1205);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx29x, QN => n_1206);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx29x, QN => n_1207);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx29x, QN => n_1208);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx29x, QN => n_1209);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx29x, QN => n_1210);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx29x, QN => n_1211);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx29x, QN => n_1212);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx29x, QN => n_1213);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx29x, QN => n_1214);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx29x, QN => n_1215);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx29x, QN => n_1216);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx29x, QN => n_1217);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx29x, QN => n_1218);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx29x, QN => n_1219);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx29x, QN => n_1220);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx29x, QN => n_1221);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx29x, QN => n_1222);
   IF_ISAxtoRegsPort_regxDSTDATAxx30x : DFF_X1 port map( D => IF_ISAxN10967, CK
                           => net6528, Q => toRegsPortxDSTDATAxx30x, QN => 
                           n_1223);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx30x, QN => n_1224);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx30x, QN => n_1225);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx30x, QN => n_1226);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx30x, QN => n_1227);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx30x, QN => n_1228);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx30x, QN => n_1229);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx30x, QN => n_1230);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx30x, QN => n_1231);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx30x, QN => n_1232);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx30x, QN => n_1233);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx30x, QN => n_1234);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx30x, QN => n_1235);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx30x, QN => n_1236);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx30x, QN => n_1237);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx30x, QN => n_1238);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx30x, QN => n_1239);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx30x, QN => n_1240);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx30x, QN => n_1241);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx30x, QN => n_1242);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx30x, QN => n_1243);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx30x, QN => n_1244);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx30x, QN => n_1245);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx30x, QN => n_1246);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx30x, QN => n_1247);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx30x, QN => n_1248);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx30x, QN => n_1249);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx30x, QN => n_1250);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx30x, QN => n_1251);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx30x, QN => n_1252);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx30x, QN => n_1253);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx30x, QN => n_1254);
   IF_ISAxtoRegsPort_regxDSTDATAxx0x : DFF_X1 port map( D => IF_ISAxN10936, CK 
                           => net6528, Q => toRegsPortxDSTDATAxx0x, QN => 
                           n_1255);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx0x, QN => n_1256);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx0x, QN => n_1257);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx0x, QN => n_1258);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx0x, QN => n_1259);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx0x, QN => n_1260);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx0x, QN => n_1261);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx0x, QN => n_1262);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx0x, QN => n_1263);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx0x, QN => n_1264);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx0x, QN => n_1265);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx0x, QN => n_1266);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx0x, QN => n_1267);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx0x, QN => n_1268);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx0x, QN => n_1269);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx0x, QN => n_1270);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx0x, QN => n_1271);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx0x, QN => n_1272);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx0x, QN => n_1273);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx0x, QN => n_1274);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx0x, QN => n_1275);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx0x, QN => n_1276);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx0x, QN => n_1277);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx0x, QN => n_1278);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx0x, QN => n_1279);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx0x, QN => n_1280);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx0x, QN => n_1281);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx0x, QN => n_1282);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx0x, QN => n_1283);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx0x, QN => n_1284);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx0x, QN => n_1285);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx0x, QN => n_1286);
   IF_ISAxtoMemoryPort_regxDATAINxx0x : DFF_X1 port map( D => n7587, CK => 
                           net6543, Q => toMemoryPortxDATAINxx0x(0), QN => 
                           n_1287);
   IF_ISAxtoRegsPort_regxDSTDATAxx16x : DFF_X1 port map( D => IF_ISAxN10953, CK
                           => net6528, Q => toRegsPortxDSTDATAxx16x, QN => 
                           n_1288);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx16x, QN => n_1289);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx16x, QN => n_1290);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx16x, QN => n_1291);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx16x, QN => n_1292);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx16x, QN => n_1293);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx16x, QN => n_1294);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx16x, QN => n_1295);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx16x, QN => n_1296);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx16x, QN => n_1297);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx16x, QN => n_1298);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx16x, QN => n_1299);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx16x, QN => n_1300);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx16x, QN => n_1301);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx16x, QN => n_1302);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx16x, QN => n_1303);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx16x, QN => n_1304);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx16x, QN => n_1305);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx16x, QN => n_1306);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx16x, QN => n_1307);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx16x, QN => n_1308);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx16x, QN => n_1309);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx16x, QN => n_1310);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx16x, QN => n_1311);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx16x, QN => n_1312);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx16x, QN => n_1313);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx16x, QN => n_1314);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx16x, QN => n_1315);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx16x, QN => n_1316);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx16x, QN => n_1317);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx16x, QN => n_1318);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx16x, QN => n_1319);
   IF_ISAxtoRegsPort_regxDSTDATAxx24x : DFF_X1 port map( D => IF_ISAxN10961, CK
                           => net6528, Q => toRegsPortxDSTDATAxx24x, QN => 
                           n_1320);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx24x, QN => n_1321);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx24x, QN => n_1322);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx24x, QN => n_1323);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx24x, QN => n_1324);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx24x, QN => n_1325);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx24x, QN => n_1326);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx24x, QN => n_1327);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx24x, QN => n_1328);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx24x, QN => n_1329);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx24x, QN => n_1330);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx24x, QN => n_1331);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx24x, QN => n_1332);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx24x, QN => n_1333);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx24x, QN => n_1334);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx24x, QN => n_1335);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx24x, QN => n_1336);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx24x, QN => n_1337);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx24x, QN => n_1338);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx24x, QN => n_1339);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx24x, QN => n_1340);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx24x, QN => n_1341);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx24x, QN => n_1342);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx24x, QN => n_1343);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx24x, QN => n_1344);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx24x, QN => n_1345);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx24x, QN => n_1346);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx24x, QN => n_1347);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx24x, QN => n_1348);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx24x, QN => n_1349);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx24x, QN => n_1350);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx24x, QN => n_1351);
   IF_ISAxtoRegsPort_regxDSTDATAxx28x : DFF_X1 port map( D => IF_ISAxN10965, CK
                           => net6528, Q => toRegsPortxDSTDATAxx28x, QN => 
                           n_1352);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx28x, QN => n_1353);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx28x, QN => n_1354);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx28x, QN => n_1355);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx28x, QN => n_1356);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx28x, QN => n_1357);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx28x, QN => n_1358);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx28x, QN => n_1359);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx28x, QN => n_1360);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx28x, QN => n_1361);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx28x, QN => n_1362);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx28x, QN => n_1363);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx28x, QN => n_1364);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx28x, QN => n_1365);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx28x, QN => n_1366);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx28x, QN => n_1367);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx28x, QN => n_1368);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx28x, QN => n_1369);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx28x, QN => n_1370);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx28x, QN => n_1371);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx28x, QN => n_1372);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx28x, QN => n_1373);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx28x, QN => n_1374);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx28x, QN => n_1375);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx28x, QN => n_1376);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx28x, QN => n_1377);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx28x, QN => n_1378);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx28x, QN => n_1379);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx28x, QN => n_1380);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx28x, QN => n_1381);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx28x, QN => n_1382);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx28x, QN => n_1383);
   IF_ISAxtoRegsPort_regxDSTDATAxx10x : DFF_X1 port map( D => IF_ISAxN10947, CK
                           => net6528, Q => toRegsPortxDSTDATAxx10x, QN => 
                           n_1384);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx10x, QN => n_1385);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx10x, QN => n_1386);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx10x, QN => n_1387);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx10x, QN => n_1388);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx10x, QN => n_1389);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx10x, QN => n_1390);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx10x, QN => n_1391);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx10x, QN => n_1392);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx10x, QN => n_1393);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx10x, QN => n_1394);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx10x, QN => n_1395);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx10x, QN => n_1396);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx10x, QN => n_1397);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx10x, QN => n_1398);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx10x, QN => n_1399);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx10x, QN => n_1400);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx10x, QN => n_1401);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx10x, QN => n_1402);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx10x, QN => n_1403);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx10x, QN => n_1404);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx10x, QN => n_1405);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx10x, QN => n_1406);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx10x, QN => n_1407);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx10x, QN => n_1408);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx10x, QN => n_1409);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx10x, QN => n_1410);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx10x, QN => n_1411);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx10x, QN => n_1412);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx10x, QN => n_1413);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx10x, QN => n_1414);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx10x, QN => n_1415);
   IF_ISAxtoRegsPort_regxDSTDATAxx26x : DFF_X1 port map( D => IF_ISAxN10963, CK
                           => net6528, Q => toRegsPortxDSTDATAxx26x, QN => 
                           n_1416);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx26x, QN => n_1417);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx26x, QN => n_1418);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx26x, QN => n_1419);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx26x, QN => n_1420);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx26x, QN => n_1421);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx26x, QN => n_1422);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx26x, QN => n_1423);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx26x, QN => n_1424);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx26x, QN => n_1425);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx26x, QN => n_1426);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx26x, QN => n_1427);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx26x, QN => n_1428);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx26x, QN => n_1429);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx26x, QN => n_1430);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx26x, QN => n_1431);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx26x, QN => n_1432);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx26x, QN => n_1433);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx26x, QN => n_1434);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx26x, QN => n_1435);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx26x, QN => n_1436);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx26x, QN => n_1437);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx26x, QN => n_1438);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx26x, QN => n_1439);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx26x, QN => n_1440);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx26x, QN => n_1441);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx26x, QN => n_1442);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx26x, QN => n_1443);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx26x, QN => n_1444);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx26x, QN => n_1445);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx26x, QN => n_1446);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx26x, QN => n_1447);
   IF_ISAxtoRegsPort_regxDSTDATAxx12x : DFF_X1 port map( D => IF_ISAxN10949, CK
                           => net6528, Q => toRegsPortxDSTDATAxx12x, QN => 
                           n_1448);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx12x, QN => n_1449);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx12x, QN => n_1450);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx12x, QN => n_1451);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx12x, QN => n_1452);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx12x, QN => n_1453);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx12x, QN => n_1454);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx12x, QN => n_1455);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx12x, QN => n_1456);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx12x, QN => n_1457);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx12x, QN => n_1458);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx12x, QN => n_1459);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx12x, QN => n_1460);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx12x, QN => n_1461);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx12x, QN => n_1462);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx12x, QN => n_1463);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx12x, QN => n_1464);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx12x, QN => n_1465);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx12x, QN => n_1466);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx12x, QN => n_1467);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx12x, QN => n_1468);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx12x, QN => n_1469);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx12x, QN => n_1470);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx12x, QN => n_1471);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx12x, QN => n_1472);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx12x, QN => n_1473);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx12x, QN => n_1474);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx12x, QN => n_1475);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx12x, QN => n_1476);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx12x, QN => n_1477);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx12x, QN => n_1478);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx12x, QN => n_1479);
   IF_ISAxtoRegsPort_regxDSTDATAxx20x : DFF_X1 port map( D => IF_ISAxN10957, CK
                           => net6528, Q => toRegsPortxDSTDATAxx20x, QN => 
                           n_1480);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx20x, QN => n_1481);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx20x, QN => n_1482);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx20x, QN => n_1483);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx20x, QN => n_1484);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx20x, QN => n_1485);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx20x, QN => n_1486);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx20x, QN => n_1487);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx20x, QN => n_1488);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx20x, QN => n_1489);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx20x, QN => n_1490);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx20x, QN => n_1491);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx20x, QN => n_1492);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx20x, QN => n_1493);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx20x, QN => n_1494);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx20x, QN => n_1495);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx20x, QN => n_1496);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx20x, QN => n_1497);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx20x, QN => n_1498);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx20x, QN => n_1499);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx20x, QN => n_1500);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx20x, QN => n_1501);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx20x, QN => n_1502);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx20x, QN => n_1503);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx20x, QN => n_1504);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx20x, QN => n_1505);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx20x, QN => n_1506);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx20x, QN => n_1507);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx20x, QN => n_1508);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx20x, QN => n_1509);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx20x, QN => n_1510);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx20x, QN => n_1511);
   IF_ISAxtoRegsPort_regxDSTDATAxx22x : DFF_X1 port map( D => IF_ISAxN10959, CK
                           => net6528, Q => toRegsPortxDSTDATAxx22x, QN => 
                           n_1512);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx22x, QN => n_1513);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx22x, QN => n_1514);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx22x, QN => n_1515);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx22x, QN => n_1516);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx22x, QN => n_1517);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx22x, QN => n_1518);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx22x, QN => n_1519);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx22x, QN => n_1520);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx22x, QN => n_1521);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx22x, QN => n_1522);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx22x, QN => n_1523);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx22x, QN => n_1524);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx22x, QN => n_1525);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx22x, QN => n_1526);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx22x, QN => n_1527);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx22x, QN => n_1528);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx22x, QN => n_1529);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx22x, QN => n_1530);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx22x, QN => n_1531);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx22x, QN => n_1532);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx22x, QN => n_1533);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx22x, QN => n_1534);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx22x, QN => n_1535);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx22x, QN => n_1536);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx22x, QN => n_1537);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx22x, QN => n_1538);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx22x, QN => n_1539);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx22x, QN => n_1540);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx22x, QN => n_1541);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx22x, QN => n_1542);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx22x, QN => n_1543);
   IF_ISAxtoRegsPort_regxDSTDATAxx8x : DFF_X1 port map( D => IF_ISAxN10945, CK 
                           => net6528, Q => toRegsPortxDSTDATAxx8x, QN => 
                           n_1544);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx8x, QN => n_1545);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx8x, QN => n_1546);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx8x, QN => n_1547);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx8x, QN => n_1548);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx8x, QN => n_1549);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx8x, QN => n_1550);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx8x, QN => n_1551);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx8x, QN => n_1552);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx8x, QN => n_1553);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx8x, QN => n_1554);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx8x, QN => n_1555);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx8x, QN => n_1556);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx8x, QN => n_1557);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx8x, QN => n_1558);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx8x, QN => n_1559);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx8x, QN => n_1560);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx8x, QN => n_1561);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx8x, QN => n_1562);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx8x, QN => n_1563);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx8x, QN => n_1564);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx8x, QN => n_1565);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx8x, QN => n_1566);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx8x, QN => n_1567);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx8x, QN => n_1568);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx8x, QN => n_1569);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx8x, QN => n_1570);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx8x, QN => n_1571);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx8x, QN => n_1572);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx8x, QN => n_1573);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx8x, QN => n_1574);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx8x, QN => n_1575);
   IF_ISAxtoRegsPort_regxDSTDATAxx11x : DFF_X1 port map( D => IF_ISAxN10948, CK
                           => net6528, Q => toRegsPortxDSTDATAxx11x, QN => 
                           n_1576);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx11x, QN => n_1577);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx11x, QN => n_1578);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx11x, QN => n_1579);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx11x, QN => n_1580);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx11x, QN => n_1581);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx11x, QN => n_1582);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx11x, QN => n_1583);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx11x, QN => n_1584);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx11x, QN => n_1585);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx11x, QN => n_1586);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx11x, QN => n_1587);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx11x, QN => n_1588);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx11x, QN => n_1589);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx11x, QN => n_1590);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx11x, QN => n_1591);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx11x, QN => n_1592);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx11x, QN => n_1593);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx11x, QN => n_1594);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx11x, QN => n_1595);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx11x, QN => n_1596);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx11x, QN => n_1597);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx11x, QN => n_1598);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx11x, QN => n_1599);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx11x, QN => n_1600);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx11x, QN => n_1601);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx11x, QN => n_1602);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx11x, QN => n_1603);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx11x, QN => n_1604);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx11x, QN => n_1605);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx11x, QN => n_1606);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx11x, QN => n_1607);
   IF_ISAxtoRegsPort_regxDSTDATAxx13x : DFF_X1 port map( D => IF_ISAxN10950, CK
                           => net6528, Q => toRegsPortxDSTDATAxx13x, QN => 
                           n_1608);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx13x, QN => n_1609);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx13x, QN => n_1610);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx13x, QN => n_1611);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx13x, QN => n_1612);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx13x, QN => n_1613);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx13x, QN => n_1614);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx13x, QN => n_1615);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx13x, QN => n_1616);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx13x, QN => n_1617);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx13x, QN => n_1618);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx13x, QN => n_1619);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx13x, QN => n_1620);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx13x, QN => n_1621);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx13x, QN => n_1622);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx13x, QN => n_1623);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx13x, QN => n_1624);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx13x, QN => n_1625);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx13x, QN => n_1626);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx13x, QN => n_1627);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx13x, QN => n_1628);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx13x, QN => n_1629);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx13x, QN => n_1630);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx13x, QN => n_1631);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx13x, QN => n_1632);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx13x, QN => n_1633);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx13x, QN => n_1634);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx13x, QN => n_1635);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx13x, QN => n_1636);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx13x, QN => n_1637);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx13x, QN => n_1638);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx13x, QN => n_1639);
   IF_ISAxtoRegsPort_regxDSTDATAxx14x : DFF_X1 port map( D => IF_ISAxN10951, CK
                           => net6528, Q => toRegsPortxDSTDATAxx14x, QN => 
                           n_1640);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx14x, QN => n_1641);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx14x, QN => n_1642);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx14x, QN => n_1643);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx14x, QN => n_1644);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx14x, QN => n_1645);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx14x, QN => n_1646);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx14x, QN => n_1647);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx14x, QN => n_1648);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx14x, QN => n_1649);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx14x, QN => n_1650);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx14x, QN => n_1651);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx14x, QN => n_1652);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx14x, QN => n_1653);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx14x, QN => n_1654);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx14x, QN => n_1655);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx14x, QN => n_1656);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx14x, QN => n_1657);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx14x, QN => n_1658);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx14x, QN => n_1659);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx14x, QN => n_1660);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx14x, QN => n_1661);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx14x, QN => n_1662);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx14x, QN => n_1663);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx14x, QN => n_1664);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx14x, QN => n_1665);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx14x, QN => n_1666);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx14x, QN => n_1667);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx14x, QN => n_1668);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx14x, QN => n_1669);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx14x, QN => n_1670);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx14x, QN => n_1671);
   IF_ISAxtoRegsPort_regxDSTDATAxx4x : DFF_X1 port map( D => IF_ISAxN10941, CK 
                           => net6528, Q => toRegsPortxDSTDATAxx4x, QN => 
                           n_1672);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx4x, QN => n_1673);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx4x, QN => n_1674);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx4x, QN => n_1675);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx4x, QN => n_1676);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx4x, QN => n_1677);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx4x, QN => n_1678);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx4x, QN => n_1679);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx4x, QN => n_1680);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx4x, QN => n_1681);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx4x, QN => n_1682);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx4x, QN => n_1683);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx4x, QN => n_1684);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx4x, QN => n_1685);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx4x, QN => n_1686);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx4x, QN => n_1687);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx4x, QN => n_1688);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx4x, QN => n_1689);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx4x, QN => n_1690);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx4x, QN => n_1691);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx4x, QN => n_1692);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx4x, QN => n_1693);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx4x, QN => n_1694);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx4x, QN => n_1695);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx4x, QN => n_1696);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx4x, QN => n_1697);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx4x, QN => n_1698);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx4x, QN => n_1699);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx4x, QN => n_1700);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx4x, QN => n_1701);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx4x, QN => n_1702);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx4x, QN => n_1703);
   IF_ISAxtoMemoryPort_regxDATAINxx4x : DFF_X1 port map( D => n7586, CK => 
                           net6543, Q => toMemoryPortxDATAINxx4x(0), QN => 
                           n_1704);
   IF_ISAxtoRegsPort_regxDSTDATAxx17x : DFF_X1 port map( D => IF_ISAxN10954, CK
                           => net6528, Q => toRegsPortxDSTDATAxx17x, QN => 
                           n_1705);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx17x, QN => n_1706);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx17x, QN => n_1707);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx17x, QN => n_1708);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx17x, QN => n_1709);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx17x, QN => n_1710);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx17x, QN => n_1711);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx17x, QN => n_1712);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx17x, QN => n_1713);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx17x, QN => n_1714);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx17x, QN => n_1715);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx17x, QN => n_1716);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx17x, QN => n_1717);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx17x, QN => n_1718);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx17x, QN => n_1719);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx17x, QN => n_1720);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx17x, QN => n_1721);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx17x, QN => n_1722);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx17x, QN => n_1723);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx17x, QN => n_1724);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx17x, QN => n_1725);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx17x, QN => n_1726);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx17x, QN => n_1727);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx17x, QN => n_1728);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx17x, QN => n_1729);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx17x, QN => n_1730);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx17x, QN => n_1731);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx17x, QN => n_1732);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx17x, QN => n_1733);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx17x, QN => n_1734);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx17x, QN => n_1735);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx17x, QN => n_1736);
   IF_ISAxtoRegsPort_regxDSTDATAxx25x : DFF_X1 port map( D => IF_ISAxN10962, CK
                           => net6528, Q => toRegsPortxDSTDATAxx25x, QN => 
                           n_1737);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx25x, QN => n_1738);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx25x, QN => n_1739);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx25x, QN => n_1740);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx25x, QN => n_1741);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx25x, QN => n_1742);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx25x, QN => n_1743);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx25x, QN => n_1744);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx25x, QN => n_1745);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx25x, QN => n_1746);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx25x, QN => n_1747);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx25x, QN => n_1748);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx25x, QN => n_1749);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx25x, QN => n_1750);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx25x, QN => n_1751);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx25x, QN => n_1752);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx25x, QN => n_1753);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx25x, QN => n_1754);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx25x, QN => n_1755);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx25x, QN => n_1756);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx25x, QN => n_1757);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx25x, QN => n_1758);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx25x, QN => n_1759);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx25x, QN => n_1760);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx25x, QN => n_1761);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx25x, QN => n_1762);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx25x, QN => n_1763);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx25x, QN => n_1764);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx25x, QN => n_1765);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx25x, QN => n_1766);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx25x, QN => n_1767);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx25x, QN => n_1768);
   IF_ISAxtoRegsPort_regxDSTDATAxx18x : DFF_X1 port map( D => IF_ISAxN10955, CK
                           => net6528, Q => toRegsPortxDSTDATAxx18x, QN => 
                           n_1769);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx18x, QN => n_1770);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx18x, QN => n_1771);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx18x, QN => n_1772);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx18x, QN => n_1773);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx18x, QN => n_1774);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx18x, QN => n_1775);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx18x, QN => n_1776);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx18x, QN => n_1777);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx18x, QN => n_1778);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx18x, QN => n_1779);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx18x, QN => n_1780);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx18x, QN => n_1781);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx18x, QN => n_1782);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx18x, QN => n_1783);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx18x, QN => n_1784);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx18x, QN => n_1785);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx18x, QN => n_1786);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx18x, QN => n_1787);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx18x, QN => n_1788);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx18x, QN => n_1789);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx18x, QN => n_1790);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx18x, QN => n_1791);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx18x, QN => n_1792);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx18x, QN => n_1793);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx18x, QN => n_1794);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx18x, QN => n_1795);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx18x, QN => n_1796);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx18x, QN => n_1797);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx18x, QN => n_1798);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx18x, QN => n_1799);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx18x, QN => n_1800);
   IF_ISAxtoRegsPort_regxDSTDATAxx19x : DFF_X1 port map( D => IF_ISAxN10956, CK
                           => net6528, Q => toRegsPortxDSTDATAxx19x, QN => 
                           n_1801);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx19x, QN => n_1802);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx19x, QN => n_1803);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx19x, QN => n_1804);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx19x, QN => n_1805);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx19x, QN => n_1806);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx19x, QN => n_1807);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx19x, QN => n_1808);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx19x, QN => n_1809);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx19x, QN => n_1810);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx19x, QN => n_1811);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx19x, QN => n_1812);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx19x, QN => n_1813);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx19x, QN => n_1814);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx19x, QN => n_1815);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx19x, QN => n_1816);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx19x, QN => n_1817);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx19x, QN => n_1818);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx19x, QN => n_1819);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx19x, QN => n_1820);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx19x, QN => n_1821);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx19x, QN => n_1822);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx19x, QN => n_1823);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx19x, QN => n_1824);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx19x, QN => n_1825);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx19x, QN => n_1826);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx19x, QN => n_1827);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx19x, QN => n_1828);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx19x, QN => n_1829);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx19x, QN => n_1830);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx19x, QN => n_1831);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx19x, QN => n_1832);
   IF_ISAxtoRegsPort_regxDSTDATAxx6x : DFF_X1 port map( D => IF_ISAxN10943, CK 
                           => net6528, Q => toRegsPortxDSTDATAxx6x, QN => 
                           n_1833);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx6x, QN => n_1834);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx6x, QN => n_1835);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx6x, QN => n_1836);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx6x, QN => n_1837);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx6x, QN => n_1838);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx6x, QN => n_1839);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx6x, QN => n_1840);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx6x, QN => n_1841);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx6x, QN => n_1842);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx6x, QN => n_1843);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx6x, QN => n_1844);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx6x, QN => n_1845);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx6x, QN => n_1846);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx6x, QN => n_1847);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx6x, QN => n_1848);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx6x, QN => n_1849);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx6x, QN => n_1850);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx6x, QN => n_1851);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx6x, QN => n_1852);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx6x, QN => n_1853);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx6x, QN => n_1854);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx6x, QN => n_1855);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx6x, QN => n_1856);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx6x, QN => n_1857);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx6x, QN => n_1858);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx6x, QN => n_1859);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx6x, QN => n_1860);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx6x, QN => n_1861);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx6x, QN => n_1862);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx6x, QN => n_1863);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx6x, QN => n_1864);
   IF_ISAxtoRegsPort_regxDSTDATAxx7x : DFF_X1 port map( D => IF_ISAxN10944, CK 
                           => net6528, Q => toRegsPortxDSTDATAxx7x, QN => 
                           n_1865);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx7x, QN => n_1866);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx7x, QN => n_1867);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx7x, QN => n_1868);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx7x, QN => n_1869);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx7x, QN => n_1870);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx7x, QN => n_1871);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx7x, QN => n_1872);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx7x, QN => n_1873);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx7x, QN => n_1874);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx7x, QN => n_1875);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx7x, QN => n_1876);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx7x, QN => n_1877);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx7x, QN => n_1878);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx7x, QN => n_1879);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx7x, QN => n_1880);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx7x, QN => n_1881);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx7x, QN => n_1882);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx7x, QN => n_1883);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx7x, QN => n_1884);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx7x, QN => n_1885);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx7x, QN => n_1886);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx7x, QN => n_1887);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx7x, QN => n_1888);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx7x, QN => n_1889);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx7x, QN => n_1890);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx7x, QN => n_1891);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx7x, QN => n_1892);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx7x, QN => n_1893);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx7x, QN => n_1894);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx7x, QN => n_1895);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx7x, QN => n_1896);
   IF_ISAxtoRegsPort_regxDSTDATAxx2x : DFF_X1 port map( D => IF_ISAxN10939, CK 
                           => net6528, Q => toRegsPortxDSTDATAxx2x, QN => 
                           n_1897);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx2x, QN => n_1898);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx2x, QN => n_1899);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx2x, QN => n_1900);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx2x, QN => n_1901);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx2x, QN => n_1902);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx2x, QN => n_1903);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx2x, QN => n_1904);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx2x, QN => n_1905);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx2x, QN => n_1906);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx2x, QN => n_1907);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx2x, QN => n_1908);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx2x, QN => n_1909);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx2x, QN => n_1910);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx2x, QN => n_1911);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx2x, QN => n_1912);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx2x, QN => n_1913);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx2x, QN => n_1914);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx2x, QN => n_1915);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx2x, QN => n_1916);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx2x, QN => n_1917);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx2x, QN => n_1918);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx2x, QN => n_1919);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx2x, QN => n_1920);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx2x, QN => n_1921);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx2x, QN => n_1922);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx2x, QN => n_1923);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx2x, QN => n_1924);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx2x, QN => n_1925);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx2x, QN => n_1926);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx2x, QN => n_1927);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx2x, QN => n_1928);
   IF_ISAxtoMemoryPort_regxDATAINxx2x : DFF_X1 port map( D => n7585, CK => 
                           net6543, Q => toMemoryPortxDATAINxx2x(0), QN => 
                           n_1929);
   IF_ISAxtoRegsPort_regxDSTDATAxx3x : DFF_X1 port map( D => IF_ISAxN10940, CK 
                           => net6528, Q => toRegsPortxDSTDATAxx3x, QN => 
                           n_1930);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx3x, QN => n_1931);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx3x, QN => n_1932);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx3x, QN => n_1933);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx3x, QN => n_1934);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx3x, QN => n_1935);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx3x, QN => n_1936);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx3x, QN => n_1937);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx3x, QN => n_1938);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx3x, QN => n_1939);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx3x, QN => n_1940);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx3x, QN => n_1941);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx3x, QN => n_1942);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx3x, QN => n_1943);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx3x, QN => n_1944);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx3x, QN => n_1945);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx3x, QN => n_1946);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx3x, QN => n_1947);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx3x, QN => n_1948);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx3x, QN => n_1949);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx3x, QN => n_1950);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx3x, QN => n_1951);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx3x, QN => n_1952);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx3x, QN => n_1953);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx3x, QN => n_1954);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx3x, QN => n_1955);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx3x, QN => n_1956);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx3x, QN => n_1957);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx3x, QN => n_1958);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx3x, QN => n_1959);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx3x, QN => n_1960);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx3x, QN => n_1961);
   IF_ISAxtoMemoryPort_regxDATAINxx3x : DFF_X1 port map( D => n7584, CK => 
                           net6543, Q => toMemoryPortxDATAINxx3x(0), QN => 
                           n_1962);
   IF_ISAxtoRegsPort_regxDSTDATAxx21x : DFF_X1 port map( D => IF_ISAxN10958, CK
                           => net6528, Q => toRegsPortxDSTDATAxx21x, QN => 
                           n_1963);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx21x, QN => n_1964);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx21x, QN => n_1965);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx21x, QN => n_1966);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx21x, QN => n_1967);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx21x, QN => n_1968);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx21x, QN => n_1969);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx21x, QN => n_1970);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx21x, QN => n_1971);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx21x, QN => n_1972);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx21x, QN => n_1973);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx21x, QN => n_1974);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx21x, QN => n_1975);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx21x, QN => n_1976);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx21x, QN => n_1977);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx21x, QN => n_1978);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx21x, QN => n_1979);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx21x, QN => n_1980);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx21x, QN => n_1981);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx21x, QN => n_1982);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx21x, QN => n_1983);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx21x, QN => n_1984);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx21x, QN => n_1985);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx21x, QN => n_1986);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx21x, QN => n_1987);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx21x, QN => n_1988);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx21x, QN => n_1989);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx21x, QN => n_1990);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx21x, QN => n_1991);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx21x, QN => n_1992);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx21x, QN => n_1993);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx21x, QN => n_1994);
   IF_ISAxtoRegsPort_regxDSTDATAxx5x : DFF_X1 port map( D => IF_ISAxN10942, CK 
                           => net6528, Q => toRegsPortxDSTDATAxx5x, QN => 
                           n_1995);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx5x, QN => n_1996);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx5x, QN => n_1997);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx5x, QN => n_1998);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx5x, QN => n_1999);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx5x, QN => n_2000);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx5x, QN => n_2001);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx5x, QN => n_2002);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx5x, QN => n_2003);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx5x, QN => n_2004);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx5x, QN => n_2005);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx5x, QN => n_2006);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx5x, QN => n_2007);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx5x, QN => n_2008);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx5x, QN => n_2009);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx5x, QN => n_2010);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx5x, QN => n_2011);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx5x, QN => n_2012);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx5x, QN => n_2013);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx5x, QN => n_2014);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx5x, QN => n_2015);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx5x, QN => n_2016);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx5x, QN => n_2017);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx5x, QN => n_2018);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx5x, QN => n_2019);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx5x, QN => n_2020);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx5x, QN => n_2021);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx5x, QN => n_2022);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx5x, QN => n_2023);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx5x, QN => n_2024);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx5x, QN => n_2025);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx5x, QN => n_2026);
   IF_ISAxtoRegsPort_regxDSTDATAxx9x : DFF_X1 port map( D => IF_ISAxN10946, CK 
                           => net6528, Q => toRegsPortxDSTDATAxx9x, QN => 
                           n_2027);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx9x, QN => n_2028);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx9x, QN => n_2029);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx9x, QN => n_2030);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx9x, QN => n_2031);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx9x, QN => n_2032);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx9x, QN => n_2033);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx9x, QN => n_2034);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx9x, QN => n_2035);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx9x, QN => n_2036);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx9x, QN => n_2037);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx9x, QN => n_2038);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx9x, QN => n_2039);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx9x, QN => n_2040);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx9x, QN => n_2041);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx9x, QN => n_2042);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx9x, QN => n_2043);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx9x, QN => n_2044);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx9x, QN => n_2045);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx9x, QN => n_2046);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx9x, QN => n_2047);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx9x, QN => n_2048);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx9x, QN => n_2049);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx9x, QN => n_2050);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx9x, QN => n_2051);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx9x, QN => n_2052);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx9x, QN => n_2053);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx9x, QN => n_2054);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx9x, QN => n_2055);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx9x, QN => n_2056);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx9x, QN => n_2057);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx9x, QN => n_2058);
   IF_ISAxtoRegsPort_regxDSTDATAxx1x : DFF_X1 port map( D => IF_ISAxN10938, CK 
                           => net6528, Q => toRegsPortxDSTDATAxx1x, QN => 
                           n_2059);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6553, Q => 
                           fromRegsPortxREG_FILE_31xx1x, QN => n_2060);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6703, Q => 
                           fromRegsPortxREG_FILE_01xx1x, QN => n_2061);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6698, Q => 
                           fromRegsPortxREG_FILE_02xx1x, QN => n_2062);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6693, Q => 
                           fromRegsPortxREG_FILE_03xx1x, QN => n_2063);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6688, Q => 
                           fromRegsPortxREG_FILE_04xx1x, QN => n_2064);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6683, Q => 
                           fromRegsPortxREG_FILE_05xx1x, QN => n_2065);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6678, Q => 
                           fromRegsPortxREG_FILE_06xx1x, QN => n_2066);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6673, Q => 
                           fromRegsPortxREG_FILE_07xx1x, QN => n_2067);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6668, Q => 
                           fromRegsPortxREG_FILE_08xx1x, QN => n_2068);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6663, Q => 
                           fromRegsPortxREG_FILE_09xx1x, QN => n_2069);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6658, Q => 
                           fromRegsPortxREG_FILE_10xx1x, QN => n_2070);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6653, Q => 
                           fromRegsPortxREG_FILE_11xx1x, QN => n_2071);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6648, Q => 
                           fromRegsPortxREG_FILE_12xx1x, QN => n_2072);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6643, Q => 
                           fromRegsPortxREG_FILE_13xx1x, QN => n_2073);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6638, Q => 
                           fromRegsPortxREG_FILE_14xx1x, QN => n_2074);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6633, Q => 
                           fromRegsPortxREG_FILE_15xx1x, QN => n_2075);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6628, Q => 
                           fromRegsPortxREG_FILE_16xx1x, QN => n_2076);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6623, Q => 
                           fromRegsPortxREG_FILE_17xx1x, QN => n_2077);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6618, Q => 
                           fromRegsPortxREG_FILE_18xx1x, QN => n_2078);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6613, Q => 
                           fromRegsPortxREG_FILE_19xx1x, QN => n_2079);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6608, Q => 
                           fromRegsPortxREG_FILE_20xx1x, QN => n_2080);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6603, Q => 
                           fromRegsPortxREG_FILE_21xx1x, QN => n_2081);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6598, Q => 
                           fromRegsPortxREG_FILE_22xx1x, QN => n_2082);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6593, Q => 
                           fromRegsPortxREG_FILE_23xx1x, QN => n_2083);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6588, Q => 
                           fromRegsPortxREG_FILE_24xx1x, QN => n_2084);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6583, Q => 
                           fromRegsPortxREG_FILE_25xx1x, QN => n_2085);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6578, Q => 
                           fromRegsPortxREG_FILE_26xx1x, QN => n_2086);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6573, Q => 
                           fromRegsPortxREG_FILE_27xx1x, QN => n_2087);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6568, Q => 
                           fromRegsPortxREG_FILE_28xx1x, QN => n_2088);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6563, Q => 
                           fromRegsPortxREG_FILE_29xx1x, QN => n_2089);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net6558, Q => 
                           fromRegsPortxREG_FILE_30xx1x, QN => n_2090);
   IF_ISAxtoMemoryPort_regxDATAINxx1x : DFF_X1 port map( D => n7583, CK => 
                           net6543, Q => toMemoryPortxDATAINxx1x(0), QN => 
                           n_2091);
   IF_ISAxtoMemoryPort_regxDATAINxx9x : DFF_X1 port map( D => IF_ISAxN10846, CK
                           => net6543, Q => toMemoryPortxDATAINxx9x(0), QN => 
                           n_2092);
   IF_ISAxtoMemoryPort_regxDATAINxx5x : DFF_X1 port map( D => IF_ISAxN10842, CK
                           => net6543, Q => toMemoryPortxDATAINxx5x(0), QN => 
                           n_2093);
   IF_ISAxtoMemoryPort_regxDATAINxx21x : DFF_X1 port map( D => IF_ISAxN10858, 
                           CK => net6543, Q => toMemoryPortxDATAINxx21x(0), QN 
                           => n_2094);
   IF_ISAxtoMemoryPort_regxDATAINxx7x : DFF_X1 port map( D => IF_ISAxN10844, CK
                           => net6543, Q => toMemoryPortxDATAINxx7x(0), QN => 
                           n_2095);
   IF_ISAxtoMemoryPort_regxDATAINxx6x : DFF_X1 port map( D => IF_ISAxN10843, CK
                           => net6543, Q => toMemoryPortxDATAINxx6x(0), QN => 
                           n_2096);
   IF_ISAxtoMemoryPort_regxDATAINxx19x : DFF_X1 port map( D => IF_ISAxN10856, 
                           CK => net6543, Q => toMemoryPortxDATAINxx19x(0), QN 
                           => n_2097);
   IF_ISAxtoMemoryPort_regxDATAINxx18x : DFF_X1 port map( D => IF_ISAxN10855, 
                           CK => net6543, Q => toMemoryPortxDATAINxx18x(0), QN 
                           => n_2098);
   IF_ISAxtoMemoryPort_regxDATAINxx25x : DFF_X1 port map( D => IF_ISAxN10862, 
                           CK => net6543, Q => toMemoryPortxDATAINxx25x(0), QN 
                           => n_2099);
   IF_ISAxtoMemoryPort_regxDATAINxx17x : DFF_X1 port map( D => IF_ISAxN10854, 
                           CK => net6543, Q => toMemoryPortxDATAINxx17x(0), QN 
                           => n_2100);
   IF_ISAxtoMemoryPort_regxDATAINxx14x : DFF_X1 port map( D => IF_ISAxN10851, 
                           CK => net6543, Q => toMemoryPortxDATAINxx14x(0), QN 
                           => n_2101);
   IF_ISAxtoMemoryPort_regxDATAINxx13x : DFF_X1 port map( D => IF_ISAxN10850, 
                           CK => net6543, Q => toMemoryPortxDATAINxx13x(0), QN 
                           => n_2102);
   IF_ISAxtoMemoryPort_regxDATAINxx11x : DFF_X1 port map( D => IF_ISAxN10848, 
                           CK => net6543, Q => toMemoryPortxDATAINxx11x(0), QN 
                           => n_2103);
   IF_ISAxtoMemoryPort_regxDATAINxx8x : DFF_X1 port map( D => IF_ISAxN10845, CK
                           => net6543, Q => toMemoryPortxDATAINxx8x(0), QN => 
                           n_2104);
   IF_ISAxtoMemoryPort_regxDATAINxx22x : DFF_X1 port map( D => IF_ISAxN10859, 
                           CK => net6543, Q => toMemoryPortxDATAINxx22x(0), QN 
                           => n_2105);
   IF_ISAxtoMemoryPort_regxDATAINxx20x : DFF_X1 port map( D => IF_ISAxN10857, 
                           CK => net6543, Q => toMemoryPortxDATAINxx20x(0), QN 
                           => n_2106);
   IF_ISAxtoMemoryPort_regxDATAINxx12x : DFF_X1 port map( D => IF_ISAxN10849, 
                           CK => net6543, Q => toMemoryPortxDATAINxx12x(0), QN 
                           => n_2107);
   IF_ISAxtoMemoryPort_regxDATAINxx26x : DFF_X1 port map( D => IF_ISAxN10863, 
                           CK => net6543, Q => toMemoryPortxDATAINxx26x(0), QN 
                           => n_2108);
   IF_ISAxtoMemoryPort_regxDATAINxx10x : DFF_X1 port map( D => IF_ISAxN10847, 
                           CK => net6543, Q => toMemoryPortxDATAINxx10x(0), QN 
                           => n_2109);
   IF_ISAxtoMemoryPort_regxDATAINxx28x : DFF_X1 port map( D => IF_ISAxN10865, 
                           CK => net6543, Q => toMemoryPortxDATAINxx28x(0), QN 
                           => n_2110);
   IF_ISAxtoMemoryPort_regxDATAINxx24x : DFF_X1 port map( D => IF_ISAxN10861, 
                           CK => net6543, Q => toMemoryPortxDATAINxx24x(0), QN 
                           => n_2111);
   IF_ISAxtoMemoryPort_regxDATAINxx16x : DFF_X1 port map( D => IF_ISAxN10853, 
                           CK => net6543, Q => toMemoryPortxDATAINxx16x(0), QN 
                           => n_2112);
   IF_ISAxtoMemoryPort_regxDATAINxx30x : DFF_X1 port map( D => IF_ISAxN10867, 
                           CK => net6543, Q => toMemoryPortxDATAINxx30x(0), QN 
                           => n_2113);
   IF_ISAxtoMemoryPort_regxDATAINxx29x : DFF_X1 port map( D => IF_ISAxN10866, 
                           CK => net6543, Q => toMemoryPortxDATAINxx29x(0), QN 
                           => n_2114);
   IF_ISAxtoMemoryPort_regxDATAINxx27x : DFF_X1 port map( D => IF_ISAxN10864, 
                           CK => net6543, Q => toMemoryPortxDATAINxx27x(0), QN 
                           => n_2115);
   IF_ISAxtoMemoryPort_regxDATAINxx23x : DFF_X1 port map( D => IF_ISAxN10860, 
                           CK => net6543, Q => toMemoryPortxDATAINxx23x(0), QN 
                           => n_2116);
   IF_ISAxtoMemoryPort_regxDATAINxx15x : DFF_X1 port map( D => IF_ISAxN10852, 
                           CK => net6543, Q => toMemoryPortxDATAINxx15x(0), QN 
                           => n_2117);
   IF_ISAxtoMemoryPort_regxDATAINxx31x : DFF_X1 port map( D => IF_ISAxN10868, 
                           CK => net6543, Q => toMemoryPortxDATAINxx31x(0), QN 
                           => n_2118);
   DP_OP_679J1_122_3096xU33 : FA_X1 port map( A => ashr_25xAx0x, B => n7547, CI
                           => DP_OP_679J1_122_3096xn68, CO => 
                           DP_OP_679J1_122_3096xn32, S => 
                           DP_OP_679J1_122_3096xn69);
   DP_OP_679J1_122_3096xU32 : FA_X1 port map( A => DP_OP_679J1_122_3096xn67, B 
                           => ashr_25xAx1x, CI => DP_OP_679J1_122_3096xn32, CO 
                           => DP_OP_679J1_122_3096xn31, S => 
                           DP_OP_679J1_122_3096xn70);
   DP_OP_679J1_122_3096xU31 : FA_X1 port map( A => DP_OP_679J1_122_3096xn66, B 
                           => ashr_25xAx2x, CI => DP_OP_679J1_122_3096xn31, CO 
                           => DP_OP_679J1_122_3096xn30, S => 
                           DP_OP_679J1_122_3096xn71);
   DP_OP_679J1_122_3096xU30 : FA_X1 port map( A => DP_OP_679J1_122_3096xn65, B 
                           => ashr_25xAx3x, CI => DP_OP_679J1_122_3096xn30, CO 
                           => DP_OP_679J1_122_3096xn29, S => 
                           DP_OP_679J1_122_3096xn72);
   DP_OP_679J1_122_3096xU29 : FA_X1 port map( A => DP_OP_679J1_122_3096xn64, B 
                           => ashr_25xAx4x, CI => DP_OP_679J1_122_3096xn29, CO 
                           => DP_OP_679J1_122_3096xn28, S => 
                           DP_OP_679J1_122_3096xn73);
   DP_OP_679J1_122_3096xU28 : FA_X1 port map( A => DP_OP_679J1_122_3096xn63, B 
                           => ashr_25xAx5x, CI => DP_OP_679J1_122_3096xn28, CO 
                           => DP_OP_679J1_122_3096xn27, S => 
                           DP_OP_679J1_122_3096xn74);
   DP_OP_679J1_122_3096xU27 : FA_X1 port map( A => DP_OP_679J1_122_3096xn62, B 
                           => ashr_25xAx6x, CI => DP_OP_679J1_122_3096xn27, CO 
                           => DP_OP_679J1_122_3096xn26, S => 
                           DP_OP_679J1_122_3096xn75);
   DP_OP_679J1_122_3096xU26 : FA_X1 port map( A => DP_OP_679J1_122_3096xn61, B 
                           => ashr_25xAx7x, CI => DP_OP_679J1_122_3096xn26, CO 
                           => DP_OP_679J1_122_3096xn25, S => 
                           DP_OP_679J1_122_3096xn76);
   DP_OP_679J1_122_3096xU25 : FA_X1 port map( A => DP_OP_679J1_122_3096xn60, B 
                           => ashr_25xAx8x, CI => DP_OP_679J1_122_3096xn25, CO 
                           => DP_OP_679J1_122_3096xn24, S => 
                           DP_OP_679J1_122_3096xn77);
   DP_OP_679J1_122_3096xU24 : FA_X1 port map( A => DP_OP_679J1_122_3096xn59, B 
                           => ashr_25xAx9x, CI => DP_OP_679J1_122_3096xn24, CO 
                           => DP_OP_679J1_122_3096xn23, S => 
                           DP_OP_679J1_122_3096xn78);
   DP_OP_679J1_122_3096xU23 : FA_X1 port map( A => DP_OP_679J1_122_3096xn58, B 
                           => ashr_25xAx10x, CI => DP_OP_679J1_122_3096xn23, CO
                           => DP_OP_679J1_122_3096xn22, S => 
                           DP_OP_679J1_122_3096xn79);
   DP_OP_679J1_122_3096xU22 : FA_X1 port map( A => DP_OP_679J1_122_3096xn57, B 
                           => ashr_25xAx11x, CI => DP_OP_679J1_122_3096xn22, CO
                           => DP_OP_679J1_122_3096xn21, S => 
                           DP_OP_679J1_122_3096xn80);
   DP_OP_679J1_122_3096xU21 : FA_X1 port map( A => DP_OP_679J1_122_3096xn56, B 
                           => ashr_25xAx12x, CI => DP_OP_679J1_122_3096xn21, CO
                           => DP_OP_679J1_122_3096xn20, S => 
                           DP_OP_679J1_122_3096xn81);
   DP_OP_679J1_122_3096xU20 : FA_X1 port map( A => DP_OP_679J1_122_3096xn55, B 
                           => ashr_25xAx13x, CI => DP_OP_679J1_122_3096xn20, CO
                           => DP_OP_679J1_122_3096xn19, S => 
                           DP_OP_679J1_122_3096xn82);
   DP_OP_679J1_122_3096xU19 : FA_X1 port map( A => DP_OP_679J1_122_3096xn54, B 
                           => ashr_25xAx14x, CI => DP_OP_679J1_122_3096xn19, CO
                           => DP_OP_679J1_122_3096xn18, S => 
                           DP_OP_679J1_122_3096xn83);
   DP_OP_679J1_122_3096xU18 : FA_X1 port map( A => DP_OP_679J1_122_3096xn53, B 
                           => ashr_25xAx15x, CI => DP_OP_679J1_122_3096xn18, CO
                           => DP_OP_679J1_122_3096xn17, S => 
                           DP_OP_679J1_122_3096xn84);
   DP_OP_679J1_122_3096xU17 : FA_X1 port map( A => DP_OP_679J1_122_3096xn52, B 
                           => ashr_25xAx16x, CI => DP_OP_679J1_122_3096xn17, CO
                           => DP_OP_679J1_122_3096xn16, S => 
                           DP_OP_679J1_122_3096xn85);
   DP_OP_679J1_122_3096xU16 : FA_X1 port map( A => DP_OP_679J1_122_3096xn51, B 
                           => ashr_25xAx17x, CI => DP_OP_679J1_122_3096xn16, CO
                           => DP_OP_679J1_122_3096xn15, S => 
                           DP_OP_679J1_122_3096xn86);
   DP_OP_679J1_122_3096xU15 : FA_X1 port map( A => DP_OP_679J1_122_3096xn50, B 
                           => ashr_25xAx18x, CI => DP_OP_679J1_122_3096xn15, CO
                           => DP_OP_679J1_122_3096xn14, S => 
                           DP_OP_679J1_122_3096xn87);
   DP_OP_679J1_122_3096xU14 : FA_X1 port map( A => DP_OP_679J1_122_3096xn49, B 
                           => ashr_25xAx19x, CI => DP_OP_679J1_122_3096xn14, CO
                           => DP_OP_679J1_122_3096xn13, S => 
                           DP_OP_679J1_122_3096xn88);
   DP_OP_679J1_122_3096xU13 : FA_X1 port map( A => DP_OP_679J1_122_3096xn48, B 
                           => ashr_25xAx20x, CI => DP_OP_679J1_122_3096xn13, CO
                           => DP_OP_679J1_122_3096xn12, S => 
                           DP_OP_679J1_122_3096xn89);
   DP_OP_679J1_122_3096xU12 : FA_X1 port map( A => DP_OP_679J1_122_3096xn47, B 
                           => ashr_25xAx21x, CI => DP_OP_679J1_122_3096xn12, CO
                           => DP_OP_679J1_122_3096xn11, S => 
                           DP_OP_679J1_122_3096xn90);
   DP_OP_679J1_122_3096xU11 : FA_X1 port map( A => DP_OP_679J1_122_3096xn46, B 
                           => ashr_25xAx22x, CI => DP_OP_679J1_122_3096xn11, CO
                           => DP_OP_679J1_122_3096xn10, S => 
                           DP_OP_679J1_122_3096xn91);
   DP_OP_679J1_122_3096xU10 : FA_X1 port map( A => DP_OP_679J1_122_3096xn45, B 
                           => ashr_25xAx23x, CI => DP_OP_679J1_122_3096xn10, CO
                           => DP_OP_679J1_122_3096xn9, S => 
                           DP_OP_679J1_122_3096xn92);
   DP_OP_679J1_122_3096xU9 : FA_X1 port map( A => DP_OP_679J1_122_3096xn44, B 
                           => ashr_25xAx24x, CI => DP_OP_679J1_122_3096xn9, CO 
                           => DP_OP_679J1_122_3096xn8, S => 
                           DP_OP_679J1_122_3096xn93);
   DP_OP_679J1_122_3096xU8 : FA_X1 port map( A => DP_OP_679J1_122_3096xn43, B 
                           => ashr_25xAx25x, CI => DP_OP_679J1_122_3096xn8, CO 
                           => DP_OP_679J1_122_3096xn7, S => 
                           DP_OP_679J1_122_3096xn94);
   DP_OP_679J1_122_3096xU7 : FA_X1 port map( A => DP_OP_679J1_122_3096xn42, B 
                           => ashr_25xAx26x, CI => DP_OP_679J1_122_3096xn7, CO 
                           => DP_OP_679J1_122_3096xn6, S => 
                           DP_OP_679J1_122_3096xn95);
   DP_OP_679J1_122_3096xU6 : FA_X1 port map( A => DP_OP_679J1_122_3096xn41, B 
                           => ashr_25xAx27x, CI => DP_OP_679J1_122_3096xn6, CO 
                           => DP_OP_679J1_122_3096xn5, S => 
                           DP_OP_679J1_122_3096xn96);
   DP_OP_679J1_122_3096xU5 : FA_X1 port map( A => DP_OP_679J1_122_3096xn40, B 
                           => ashr_25xAx28x, CI => DP_OP_679J1_122_3096xn5, CO 
                           => DP_OP_679J1_122_3096xn4, S => 
                           DP_OP_679J1_122_3096xn97);
   DP_OP_679J1_122_3096xU4 : FA_X1 port map( A => DP_OP_679J1_122_3096xn39, B 
                           => ashr_25xAx29x, CI => DP_OP_679J1_122_3096xn4, CO 
                           => DP_OP_679J1_122_3096xn3, S => 
                           DP_OP_679J1_122_3096xn98);
   DP_OP_679J1_122_3096xU3 : FA_X1 port map( A => DP_OP_679J1_122_3096xn38, B 
                           => ashr_25xAx30x, CI => DP_OP_679J1_122_3096xn3, CO 
                           => DP_OP_679J1_122_3096xn2, S => 
                           DP_OP_679J1_122_3096xn99);
   DP_OP_719J1_125_1055xU33 : FA_X1 port map( A => DP_OP_719J1_125_1055xn134, B
                           => n7546, CI => DP_OP_719J1_125_1055xn68, CO => 
                           DP_OP_719J1_125_1055xn32, S => 
                           DP_OP_719J1_125_1055xn69);
   DP_OP_719J1_125_1055xU32 : FA_X1 port map( A => DP_OP_719J1_125_1055xn67, B 
                           => DP_OP_719J1_125_1055xn135, CI => 
                           DP_OP_719J1_125_1055xn32, CO => 
                           DP_OP_719J1_125_1055xn31, S => 
                           DP_OP_719J1_125_1055xn70);
   DP_OP_719J1_125_1055xU31 : FA_X1 port map( A => DP_OP_719J1_125_1055xn66, B 
                           => DP_OP_719J1_125_1055xn136, CI => 
                           DP_OP_719J1_125_1055xn31, CO => 
                           DP_OP_719J1_125_1055xn30, S => 
                           DP_OP_719J1_125_1055xn71);
   DP_OP_719J1_125_1055xU30 : FA_X1 port map( A => DP_OP_719J1_125_1055xn65, B 
                           => DP_OP_719J1_125_1055xn137, CI => 
                           DP_OP_719J1_125_1055xn30, CO => 
                           DP_OP_719J1_125_1055xn29, S => 
                           DP_OP_719J1_125_1055xn72);
   DP_OP_719J1_125_1055xU29 : FA_X1 port map( A => DP_OP_719J1_125_1055xn64, B 
                           => DP_OP_719J1_125_1055xn138, CI => 
                           DP_OP_719J1_125_1055xn29, CO => 
                           DP_OP_719J1_125_1055xn28, S => 
                           DP_OP_719J1_125_1055xn73);
   DP_OP_719J1_125_1055xU28 : FA_X1 port map( A => DP_OP_719J1_125_1055xn63, B 
                           => DP_OP_719J1_125_1055xn139, CI => 
                           DP_OP_719J1_125_1055xn28, CO => 
                           DP_OP_719J1_125_1055xn27, S => 
                           DP_OP_719J1_125_1055xn74);
   DP_OP_719J1_125_1055xU27 : FA_X1 port map( A => DP_OP_719J1_125_1055xn62, B 
                           => DP_OP_719J1_125_1055xn140, CI => 
                           DP_OP_719J1_125_1055xn27, CO => 
                           DP_OP_719J1_125_1055xn26, S => 
                           DP_OP_719J1_125_1055xn75);
   DP_OP_719J1_125_1055xU26 : FA_X1 port map( A => DP_OP_719J1_125_1055xn61, B 
                           => DP_OP_719J1_125_1055xn141, CI => 
                           DP_OP_719J1_125_1055xn26, CO => 
                           DP_OP_719J1_125_1055xn25, S => 
                           DP_OP_719J1_125_1055xn76);
   DP_OP_719J1_125_1055xU25 : FA_X1 port map( A => DP_OP_719J1_125_1055xn60, B 
                           => DP_OP_719J1_125_1055xn142, CI => 
                           DP_OP_719J1_125_1055xn25, CO => 
                           DP_OP_719J1_125_1055xn24, S => 
                           DP_OP_719J1_125_1055xn77);
   DP_OP_719J1_125_1055xU24 : FA_X1 port map( A => DP_OP_719J1_125_1055xn59, B 
                           => DP_OP_719J1_125_1055xn143, CI => 
                           DP_OP_719J1_125_1055xn24, CO => 
                           DP_OP_719J1_125_1055xn23, S => 
                           DP_OP_719J1_125_1055xn78);
   DP_OP_719J1_125_1055xU23 : FA_X1 port map( A => DP_OP_719J1_125_1055xn58, B 
                           => DP_OP_719J1_125_1055xn144, CI => 
                           DP_OP_719J1_125_1055xn23, CO => 
                           DP_OP_719J1_125_1055xn22, S => 
                           DP_OP_719J1_125_1055xn79);
   DP_OP_719J1_125_1055xU22 : FA_X1 port map( A => DP_OP_719J1_125_1055xn57, B 
                           => DP_OP_719J1_125_1055xn145, CI => 
                           DP_OP_719J1_125_1055xn22, CO => 
                           DP_OP_719J1_125_1055xn21, S => 
                           DP_OP_719J1_125_1055xn80);
   DP_OP_719J1_125_1055xU21 : FA_X1 port map( A => DP_OP_719J1_125_1055xn56, B 
                           => DP_OP_719J1_125_1055xn146, CI => 
                           DP_OP_719J1_125_1055xn21, CO => 
                           DP_OP_719J1_125_1055xn20, S => 
                           DP_OP_719J1_125_1055xn81);
   DP_OP_719J1_125_1055xU20 : FA_X1 port map( A => DP_OP_719J1_125_1055xn55, B 
                           => DP_OP_719J1_125_1055xn147, CI => 
                           DP_OP_719J1_125_1055xn20, CO => 
                           DP_OP_719J1_125_1055xn19, S => 
                           DP_OP_719J1_125_1055xn82);
   DP_OP_719J1_125_1055xU19 : FA_X1 port map( A => DP_OP_719J1_125_1055xn54, B 
                           => DP_OP_719J1_125_1055xn148, CI => 
                           DP_OP_719J1_125_1055xn19, CO => 
                           DP_OP_719J1_125_1055xn18, S => 
                           DP_OP_719J1_125_1055xn83);
   DP_OP_719J1_125_1055xU18 : FA_X1 port map( A => DP_OP_719J1_125_1055xn53, B 
                           => DP_OP_719J1_125_1055xn149, CI => 
                           DP_OP_719J1_125_1055xn18, CO => 
                           DP_OP_719J1_125_1055xn17, S => 
                           DP_OP_719J1_125_1055xn84);
   DP_OP_719J1_125_1055xU17 : FA_X1 port map( A => DP_OP_719J1_125_1055xn52, B 
                           => DP_OP_719J1_125_1055xn150, CI => 
                           DP_OP_719J1_125_1055xn17, CO => 
                           DP_OP_719J1_125_1055xn16, S => 
                           DP_OP_719J1_125_1055xn85);
   DP_OP_719J1_125_1055xU16 : FA_X1 port map( A => DP_OP_719J1_125_1055xn51, B 
                           => DP_OP_719J1_125_1055xn151, CI => 
                           DP_OP_719J1_125_1055xn16, CO => 
                           DP_OP_719J1_125_1055xn15, S => 
                           DP_OP_719J1_125_1055xn86);
   DP_OP_719J1_125_1055xU15 : FA_X1 port map( A => DP_OP_719J1_125_1055xn50, B 
                           => DP_OP_719J1_125_1055xn152, CI => 
                           DP_OP_719J1_125_1055xn15, CO => 
                           DP_OP_719J1_125_1055xn14, S => 
                           DP_OP_719J1_125_1055xn87);
   DP_OP_719J1_125_1055xU14 : FA_X1 port map( A => DP_OP_719J1_125_1055xn49, B 
                           => DP_OP_719J1_125_1055xn153, CI => 
                           DP_OP_719J1_125_1055xn14, CO => 
                           DP_OP_719J1_125_1055xn13, S => 
                           DP_OP_719J1_125_1055xn88);
   DP_OP_719J1_125_1055xU13 : FA_X1 port map( A => DP_OP_719J1_125_1055xn48, B 
                           => DP_OP_719J1_125_1055xn154, CI => 
                           DP_OP_719J1_125_1055xn13, CO => 
                           DP_OP_719J1_125_1055xn12, S => 
                           DP_OP_719J1_125_1055xn89);
   DP_OP_719J1_125_1055xU12 : FA_X1 port map( A => DP_OP_719J1_125_1055xn47, B 
                           => DP_OP_719J1_125_1055xn155, CI => 
                           DP_OP_719J1_125_1055xn12, CO => 
                           DP_OP_719J1_125_1055xn11, S => 
                           DP_OP_719J1_125_1055xn90);
   DP_OP_719J1_125_1055xU11 : FA_X1 port map( A => DP_OP_719J1_125_1055xn46, B 
                           => DP_OP_719J1_125_1055xn156, CI => 
                           DP_OP_719J1_125_1055xn11, CO => 
                           DP_OP_719J1_125_1055xn10, S => 
                           DP_OP_719J1_125_1055xn91);
   DP_OP_719J1_125_1055xU10 : FA_X1 port map( A => DP_OP_719J1_125_1055xn45, B 
                           => DP_OP_719J1_125_1055xn157, CI => 
                           DP_OP_719J1_125_1055xn10, CO => 
                           DP_OP_719J1_125_1055xn9, S => 
                           DP_OP_719J1_125_1055xn92);
   DP_OP_719J1_125_1055xU9 : FA_X1 port map( A => DP_OP_719J1_125_1055xn44, B 
                           => DP_OP_719J1_125_1055xn158, CI => 
                           DP_OP_719J1_125_1055xn9, CO => 
                           DP_OP_719J1_125_1055xn8, S => 
                           DP_OP_719J1_125_1055xn93);
   DP_OP_719J1_125_1055xU8 : FA_X1 port map( A => DP_OP_719J1_125_1055xn43, B 
                           => DP_OP_719J1_125_1055xn159, CI => 
                           DP_OP_719J1_125_1055xn8, CO => 
                           DP_OP_719J1_125_1055xn7, S => 
                           DP_OP_719J1_125_1055xn94);
   DP_OP_719J1_125_1055xU7 : FA_X1 port map( A => DP_OP_719J1_125_1055xn42, B 
                           => DP_OP_719J1_125_1055xn160, CI => 
                           DP_OP_719J1_125_1055xn7, CO => 
                           DP_OP_719J1_125_1055xn6, S => 
                           DP_OP_719J1_125_1055xn95);
   DP_OP_719J1_125_1055xU6 : FA_X1 port map( A => DP_OP_719J1_125_1055xn41, B 
                           => DP_OP_719J1_125_1055xn161, CI => 
                           DP_OP_719J1_125_1055xn6, CO => 
                           DP_OP_719J1_125_1055xn5, S => 
                           DP_OP_719J1_125_1055xn96);
   DP_OP_719J1_125_1055xU5 : FA_X1 port map( A => DP_OP_719J1_125_1055xn40, B 
                           => DP_OP_719J1_125_1055xn162, CI => 
                           DP_OP_719J1_125_1055xn5, CO => 
                           DP_OP_719J1_125_1055xn4, S => 
                           DP_OP_719J1_125_1055xn97);
   DP_OP_719J1_125_1055xU4 : FA_X1 port map( A => DP_OP_719J1_125_1055xn39, B 
                           => DP_OP_719J1_125_1055xn163, CI => 
                           DP_OP_719J1_125_1055xn4, CO => 
                           DP_OP_719J1_125_1055xn3, S => 
                           DP_OP_719J1_125_1055xn98);
   DP_OP_719J1_125_1055xU3 : FA_X1 port map( A => DP_OP_719J1_125_1055xn38, B 
                           => DP_OP_719J1_125_1055xn164, CI => 
                           DP_OP_719J1_125_1055xn3, CO => 
                           DP_OP_719J1_125_1055xn2, S => 
                           DP_OP_719J1_125_1055xn99);
   intadd_0xU30 : FA_X1 port map( A => IF_ISAxpcReg_signal_2_port, B => 
                           intadd_0xBx0x, CI => intadd_0xCI, CO => intadd_0xn29
                           , S => intadd_0xSUMx0x);
   intadd_0xU29 : FA_X1 port map( A => IF_ISAxpcReg_signal_3_port, B => 
                           ashr_25xSHx3x, CI => intadd_0xn29, CO => 
                           intadd_0xn28, S => intadd_0xSUMx1x);
   intadd_0xU28 : FA_X1 port map( A => IF_ISAxpcReg_signal_4_port, B => 
                           ashr_25xSHx4x, CI => intadd_0xn28, CO => 
                           intadd_0xn27, S => intadd_0xSUMx2x);
   intadd_0xU27 : FA_X1 port map( A => IF_ISAxpcReg_signal_5_port, B => 
                           add_x_26xBx5x, CI => intadd_0xn27, CO => 
                           intadd_0xn26, S => intadd_0xSUMx3x);
   intadd_0xU26 : FA_X1 port map( A => IF_ISAxpcReg_signal_6_port, B => 
                           add_x_26xBx6x, CI => intadd_0xn26, CO => 
                           intadd_0xn25, S => intadd_0xSUMx4x);
   intadd_0xU25 : FA_X1 port map( A => IF_ISAxpcReg_signal_7_port, B => 
                           add_x_26xBx7x, CI => intadd_0xn25, CO => 
                           intadd_0xn24, S => intadd_0xSUMx5x);
   intadd_0xU24 : FA_X1 port map( A => IF_ISAxpcReg_signal_8_port, B => 
                           add_x_26xBx8x, CI => intadd_0xn24, CO => 
                           intadd_0xn23, S => intadd_0xSUMx6x);
   intadd_0xU23 : FA_X1 port map( A => IF_ISAxpcReg_signal_9_port, B => 
                           add_x_26xBx9x, CI => intadd_0xn23, CO => 
                           intadd_0xn22, S => intadd_0xSUMx7x);
   intadd_0xU22 : FA_X1 port map( A => IF_ISAxpcReg_signal_10_port, B => 
                           add_x_26xBx10x, CI => intadd_0xn22, CO => 
                           intadd_0xn21, S => intadd_0xSUMx8x);
   intadd_0xU21 : FA_X1 port map( A => IF_ISAxpcReg_signal_11_port, B => 
                           add_x_26xBx11x, CI => intadd_0xn21, CO => 
                           intadd_0xn20, S => intadd_0xSUMx9x);
   intadd_0xU20 : FA_X1 port map( A => IF_ISAxpcReg_signal_12_port, B => 
                           add_x_26xBx12x, CI => intadd_0xn20, CO => 
                           intadd_0xn19, S => intadd_0xSUMx10x);
   intadd_0xU19 : FA_X1 port map( A => IF_ISAxpcReg_signal_13_port, B => 
                           add_x_26xBx13x, CI => intadd_0xn19, CO => 
                           intadd_0xn18, S => intadd_0xSUMx11x);
   intadd_0xU18 : FA_X1 port map( A => IF_ISAxpcReg_signal_14_port, B => 
                           add_x_26xBx14x, CI => intadd_0xn18, CO => 
                           intadd_0xn17, S => intadd_0xSUMx12x);
   intadd_0xU17 : FA_X1 port map( A => IF_ISAxpcReg_signal_15_port, B => 
                           add_x_26xBx15x, CI => intadd_0xn17, CO => 
                           intadd_0xn16, S => intadd_0xSUMx13x);
   intadd_0xU16 : FA_X1 port map( A => IF_ISAxpcReg_signal_16_port, B => 
                           add_x_26xBx16x, CI => intadd_0xn16, CO => 
                           intadd_0xn15, S => intadd_0xSUMx14x);
   intadd_0xU15 : FA_X1 port map( A => IF_ISAxpcReg_signal_17_port, B => 
                           add_x_26xBx17x, CI => intadd_0xn15, CO => 
                           intadd_0xn14, S => intadd_0xSUMx15x);
   intadd_0xU14 : FA_X1 port map( A => IF_ISAxpcReg_signal_18_port, B => 
                           add_x_26xBx18x, CI => intadd_0xn14, CO => 
                           intadd_0xn13, S => intadd_0xSUMx16x);
   intadd_0xU13 : FA_X1 port map( A => IF_ISAxpcReg_signal_19_port, B => 
                           add_x_26xBx19x, CI => intadd_0xn13, CO => 
                           intadd_0xn12, S => intadd_0xSUMx17x);
   intadd_0xU12 : FA_X1 port map( A => IF_ISAxpcReg_signal_20_port, B => 
                           add_x_26xBx20x, CI => intadd_0xn12, CO => 
                           intadd_0xn11, S => intadd_0xSUMx18x);
   intadd_0xU11 : FA_X1 port map( A => IF_ISAxpcReg_signal_21_port, B => 
                           add_x_26xBx21x, CI => intadd_0xn11, CO => 
                           intadd_0xn10, S => intadd_0xSUMx19x);
   intadd_0xU10 : FA_X1 port map( A => IF_ISAxpcReg_signal_22_port, B => 
                           add_x_26xBx22x, CI => intadd_0xn10, CO => 
                           intadd_0xn9, S => intadd_0xSUMx20x);
   intadd_0xU9 : FA_X1 port map( A => IF_ISAxpcReg_signal_23_port, B => 
                           add_x_26xBx23x, CI => intadd_0xn9, CO => intadd_0xn8
                           , S => intadd_0xSUMx21x);
   intadd_0xU8 : FA_X1 port map( A => IF_ISAxpcReg_signal_24_port, B => 
                           add_x_26xBx24x, CI => intadd_0xn8, CO => intadd_0xn7
                           , S => intadd_0xSUMx22x);
   intadd_0xU7 : FA_X1 port map( A => IF_ISAxpcReg_signal_25_port, B => 
                           add_x_26xBx25x, CI => intadd_0xn7, CO => intadd_0xn6
                           , S => intadd_0xSUMx23x);
   intadd_0xU6 : FA_X1 port map( A => IF_ISAxpcReg_signal_26_port, B => 
                           add_x_26xBx26x, CI => intadd_0xn6, CO => intadd_0xn5
                           , S => intadd_0xSUMx24x);
   intadd_0xU5 : FA_X1 port map( A => IF_ISAxpcReg_signal_27_port, B => 
                           add_x_26xBx27x, CI => intadd_0xn5, CO => intadd_0xn4
                           , S => intadd_0xSUMx25x);
   intadd_0xU4 : FA_X1 port map( A => IF_ISAxpcReg_signal_28_port, B => 
                           add_x_26xBx28x, CI => intadd_0xn4, CO => intadd_0xn3
                           , S => intadd_0xSUMx26x);
   intadd_0xU3 : FA_X1 port map( A => IF_ISAxpcReg_signal_29_port, B => 
                           add_x_26xBx29x, CI => intadd_0xn3, CO => intadd_0xn2
                           , S => intadd_0xSUMx27x);
   intadd_0xU2 : FA_X1 port map( A => IF_ISAxpcReg_signal_30_port, B => 
                           add_x_26xBx30x, CI => intadd_0xn2, CO => intadd_0xn1
                           , S => intadd_0xSUMx28x);
   intadd_1xU9 : FA_X1 port map( A => intadd_1xAx0x, B => intadd_1xBx0x, CI => 
                           intadd_1xCI, CO => intadd_1xn8, S => intadd_1xSUMx0x
                           );
   intadd_1xU8 : FA_X1 port map( A => intadd_1xAx1x, B => intadd_1xBx1x, CI => 
                           intadd_1xn8, CO => intadd_1xn7, S => intadd_1xSUMx1x
                           );
   intadd_1xU7 : FA_X1 port map( A => intadd_1xAx2x, B => intadd_1xBx2x, CI => 
                           intadd_1xn7, CO => intadd_1xn6, S => intadd_1xSUMx2x
                           );
   intadd_1xU6 : FA_X1 port map( A => intadd_1xAx3x, B => intadd_1xBx3x, CI => 
                           intadd_1xn6, CO => intadd_1xn5, S => intadd_1xSUMx3x
                           );
   intadd_1xU5 : FA_X1 port map( A => intadd_1xAx4x, B => intadd_1xBx4x, CI => 
                           intadd_1xn5, CO => intadd_1xn4, S => intadd_1xSUMx4x
                           );
   intadd_1xU4 : FA_X1 port map( A => intadd_1xAx5x, B => intadd_1xBx5x, CI => 
                           intadd_1xn4, CO => intadd_1xn3, S => intadd_1xSUMx5x
                           );
   intadd_1xU3 : FA_X1 port map( A => intadd_1xAx6x, B => intadd_1xBx6x, CI => 
                           intadd_1xn3, CO => intadd_1xn2, S => intadd_1xSUMx6x
                           );
   intadd_1xU2 : FA_X1 port map( A => intadd_1xAx7x, B => intadd_1xBx7x, CI => 
                           intadd_1xn2, CO => intadd_1xn1, S => intadd_1xSUMx7x
                           );
   intadd_2xU5 : FA_X1 port map( A => intadd_2xAx0x, B => intadd_2xBx0x, CI => 
                           intadd_2xCI, CO => intadd_2xn4, S => intadd_2xSUMx0x
                           );
   intadd_2xU4 : FA_X1 port map( A => intadd_2xAx1x, B => intadd_2xBx1x, CI => 
                           intadd_2xn4, CO => intadd_2xn3, S => intadd_2xSUMx1x
                           );
   intadd_2xU3 : FA_X1 port map( A => intadd_2xAx2x, B => intadd_2xBx2x, CI => 
                           intadd_2xn3, CO => intadd_2xn2, S => intadd_2xSUMx2x
                           );
   intadd_2xU2 : FA_X1 port map( A => intadd_2xAx3x, B => intadd_2xBx3x, CI => 
                           intadd_2xn2, CO => intadd_2xn1, S => intadd_2xSUMx3x
                           );
   intadd_3xU4 : FA_X1 port map( A => intadd_3xAx0x, B => intadd_3xBx0x, CI => 
                           intadd_3xCI, CO => intadd_3xn3, S => intadd_3xSUMx0x
                           );
   intadd_3xU3 : FA_X1 port map( A => intadd_3xAx1x, B => intadd_3xBx1x, CI => 
                           intadd_3xn3, CO => intadd_3xn2, S => intadd_3xSUMx1x
                           );
   intadd_3xU2 : FA_X1 port map( A => intadd_3xAx2x, B => intadd_3xBx2x, CI => 
                           intadd_3xn2, CO => intadd_3xn1, S => intadd_3xSUMx2x
                           );
   intadd_4xU4 : FA_X1 port map( A => intadd_4xAx0x, B => intadd_4xBx0x, CI => 
                           intadd_4xCI, CO => intadd_4xn3, S => intadd_4xSUMx0x
                           );
   intadd_4xU3 : FA_X1 port map( A => intadd_4xAx1x, B => intadd_4xBx1x, CI => 
                           intadd_4xn3, CO => intadd_4xn2, S => intadd_4xSUMx1x
                           );
   intadd_4xU2 : FA_X1 port map( A => intadd_4xAx2x, B => intadd_4xBx2x, CI => 
                           intadd_4xn2, CO => intadd_4xn1, S => intadd_4xSUMx2x
                           );
   U3775 : AOI21_X2 port map( B1 => n7431, B2 => n7345, A => n6313, ZN => n7349
                           );
   U3776 : NOR2_X2 port map( A1 => n5716, A2 => n5715, ZN => n7248);
   U3777 : CLKBUF_X2 port map( A => n7231, Z => intadd_4xBx2x);
   U3778 : NOR2_X2 port map( A1 => n5701, A2 => n7246, ZN => n7223);
   U3779 : NOR3_X4 port map( A1 => n5713, A2 => n5716, A3 => n5712, ZN => n7315
                           );
   U3780 : AOI21_X2 port map( B1 => n5117, B2 => n5313, A => n5116, ZN => n7081
                           );
   U3781 : NAND2_X2 port map( A1 => n3564, A2 => n3563, ZN => ashr_25xSHx3x);
   U3782 : OR2_X1 port map( A1 => n3622, A2 => n3621, ZN => n3558);
   U3783 : INV_X1 port map( A => n5438, ZN => n5657);
   U3784 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(0), A2 => 
                           fromMemoryPortxLOADEDDATAx(1), ZN => n3559);
   U3785 : NOR4_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(2), A2 => 
                           fromMemoryPortxLOADEDDATAx(4), A3 => 
                           fromMemoryPortxLOADEDDATAx(3), A4 => n3559, ZN => 
                           n3561);
   U3786 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(5), A2 => n3561, 
                           ZN => n7442);
   U3787 : NAND2_X1 port map( A1 => n7442, A2 => fromMemoryPortxLOADEDDATAx(10)
                           , ZN => n3564);
   U3788 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(2), A2 => 
                           fromMemoryPortxLOADEDDATAx(6), ZN => n5769);
   U3789 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(4), ZN => n6294);
   U3790 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(5), A2 => n6294,
                           ZN => n5770);
   U3791 : NOR3_X1 port map( A1 => n5769, A2 => n3559, A3 => n5770, ZN => n7441
                           );
   U3792 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(5), ZN => n3560);
   U3793 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(6), ZN => n6388);
   U3794 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(3), ZN => n5760);
   U3795 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(4), A2 => n6388,
                           A3 => n5760, ZN => n5776);
   U3796 : NOR2_X1 port map( A1 => n3559, A2 => n5776, ZN => n6113);
   U3797 : CLKBUF_X1 port map( A => n6113, Z => n7112);
   U3798 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(2), ZN => n6182);
   U3799 : NAND2_X1 port map( A1 => n7112, A2 => n6182, ZN => n5680);
   U3800 : INV_X1 port map( A => n5680, ZN => n3565);
   U3801 : NAND2_X1 port map( A1 => n3560, A2 => n3565, ZN => n5712);
   U3802 : NAND2_X1 port map( A1 => n3561, A2 => n6388, ZN => n7486);
   U3803 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(5), A2 => n7486, 
                           ZN => n7440);
   U3804 : INV_X1 port map( A => n7440, ZN => n7448);
   U3805 : NAND2_X1 port map( A1 => n5712, A2 => n7448, ZN => n3562);
   U3806 : OR2_X1 port map( A1 => n7441, A2 => n3562, ZN => n3644);
   U3807 : NAND2_X1 port map( A1 => n3644, A2 => fromMemoryPortxLOADEDDATAx(23)
                           , ZN => n3563);
   U3808 : INV_X1 port map( A => n7441, ZN => n3570);
   U3809 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(14), A2 => 
                           fromMemoryPortxLOADEDDATAx(12), ZN => n5975);
   U3810 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(13), A2 => n5975,
                           ZN => n3601);
   U3811 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(5), A2 => n3565, 
                           ZN => n6043);
   U3812 : NOR4_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(29), A2 => 
                           fromMemoryPortxLOADEDDATAx(25), A3 => 
                           fromMemoryPortxLOADEDDATAx(27), A4 => 
                           fromMemoryPortxLOADEDDATAx(26), ZN => n3566);
   U3813 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(28), ZN => n7244);
   U3814 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(31), ZN => n7436);
   U3815 : NAND3_X1 port map( A1 => n3566, A2 => n7244, A3 => n7436, ZN => 
                           n3597);
   U3816 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(30), ZN => n7358);
   U3817 : NOR2_X1 port map( A1 => n3597, A2 => n7358, ZN => n3589);
   U3818 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(13), ZN => n6703);
   U3819 : AND2_X1 port map( A1 => n3589, A2 => n6703, ZN => n3573);
   U3820 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(12), B2 => 
                           fromMemoryPortxLOADEDDATAx(14), A => n5975, ZN => 
                           n3590);
   U3821 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(14), ZN => n6751);
   U3822 : NAND2_X1 port map( A1 => n6703, A2 => n6751, ZN => n3586);
   U3823 : OAI21_X1 port map( B1 => n3573, B2 => n3590, A => n3586, ZN => n3567
                           );
   U3824 : AND2_X1 port map( A1 => n7442, A2 => fromMemoryPortxLOADEDDATAx(6), 
                           ZN => n4875);
   U3825 : INV_X1 port map( A => n4875, ZN => n7453);
   U3826 : OAI22_X1 port map( A1 => n5712, A2 => n3567, B1 => n7453, B2 => 
                           n3590, ZN => n3568);
   U3827 : AOI21_X1 port map( B1 => n3601, B2 => n6043, A => n3568, ZN => n3569
                           );
   U3828 : AND2_X1 port map( A1 => n7442, A2 => n6388, ZN => n7456);
   U3829 : INV_X1 port map( A => n7456, ZN => n5984);
   U3830 : NAND3_X1 port map( A1 => n3570, A2 => n3569, A3 => n5984, ZN => 
                           n5700);
   U3831 : INV_X1 port map( A => n5700, ZN => n3611);
   U3832 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(30), A2 => n3597,
                           ZN => n3591);
   U3833 : INV_X1 port map( A => n3586, ZN => n5976);
   U3834 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(12), ZN => n5762);
   U3835 : NAND2_X1 port map( A1 => n5976, A2 => n5762, ZN => n3598);
   U3836 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(14), A2 => n6703
                           , ZN => n3575);
   U3837 : OAI21_X1 port map( B1 => n3591, B2 => n3598, A => n3575, ZN => n3571
                           );
   U3838 : INV_X1 port map( A => n3571, ZN => n3574);
   U3839 : INV_X1 port map( A => n6043, ZN => n5708);
   U3840 : INV_X1 port map( A => n5712, ZN => n6045);
   U3841 : OAI21_X1 port map( B1 => n3586, B2 => fromMemoryPortxLOADEDDATAx(12)
                           , A => n6045, ZN => n3584);
   U3842 : NAND2_X1 port map( A1 => n6703, A2 => n5762, ZN => n3572);
   U3843 : OAI21_X1 port map( B1 => n6751, B2 => n3573, A => n3572, ZN => n3585
                           );
   U3844 : NAND2_X1 port map( A1 => n6703, A2 => n3585, ZN => n3577);
   U3845 : INV_X1 port map( A => n7442, ZN => n3595);
   U3846 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(13), A2 => n6751
                           , ZN => n5441);
   U3847 : OAI222_X1 port map( A1 => n3574, A2 => n5708, B1 => n3584, B2 => 
                           n3577, C1 => n3595, C2 => n5441, ZN => n3608);
   U3848 : AND2_X1 port map( A1 => n7112, A2 => fromMemoryPortxLOADEDDATAx(2), 
                           ZN => n5692);
   U3849 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(13), A2 => n5762
                           , B1 => fromMemoryPortxLOADEDDATAx(12), B2 => n6703,
                           ZN => n3579);
   U3850 : INV_X1 port map( A => n3575, ZN => n3592);
   U3851 : NAND2_X1 port map( A1 => n3592, A2 => n3597, ZN => n3576);
   U3852 : AOI22_X1 port map( A1 => n6045, A2 => n3577, B1 => n6043, B2 => 
                           n3576, ZN => n3578);
   U3853 : AOI21_X1 port map( B1 => n3579, B2 => n5441, A => n3578, ZN => n3580
                           );
   U3854 : AOI211_X1 port map( C1 => fromMemoryPortxLOADEDDATAx(5), C2 => n5692
                           , A => n7456, B => n3580, ZN => n3607);
   U3855 : INV_X1 port map( A => n3607, ZN => n3613);
   U3856 : OR2_X1 port map( A1 => n3608, A2 => n3613, ZN => n3603);
   U3857 : NOR2_X1 port map( A1 => n3611, A2 => n3603, ZN => n5636);
   U3858 : AOI21_X1 port map( B1 => n4875, B2 => n3590, A => n7441, ZN => n3583
                           );
   U3859 : INV_X1 port map( A => n5441, ZN => n3581);
   U3860 : OAI221_X1 port map( B1 => n3581, B2 => n3592, C1 => n3581, C2 => 
                           fromMemoryPortxLOADEDDATAx(12), A => n6043, ZN => 
                           n3582);
   U3861 : OAI211_X1 port map( C1 => n3585, C2 => n3584, A => n3583, B => n3582
                           , ZN => n3621);
   U3862 : OAI21_X1 port map( B1 => n6703, B2 => n5975, A => n3586, ZN => n3587
                           );
   U3863 : INV_X1 port map( A => n3587, ZN => n3588);
   U3864 : AOI221_X1 port map( B1 => n3589, B2 => n3588, C1 => n5762, C2 => 
                           n3588, A => n5708, ZN => n3599);
   U3865 : AOI211_X1 port map( C1 => n3592, C2 => n3591, A => n5712, B => n3590
                           , ZN => n3593);
   U3866 : INV_X1 port map( A => n3593, ZN => n3594);
   U3867 : OAI21_X1 port map( B1 => n3595, B2 => n5762, A => n3594, ZN => n3596
                           );
   U3868 : AOI222_X1 port map( A1 => n3599, A2 => n3598, B1 => n3599, B2 => 
                           n3597, C1 => n3598, C2 => n3596, ZN => n3600);
   U3869 : INV_X1 port map( A => n3600, ZN => n3633);
   U3870 : NOR2_X1 port map( A1 => n3621, A2 => n3633, ZN => n3609);
   U3871 : OAI21_X1 port map( B1 => n3601, B2 => n7453, A => n5708, ZN => n3602
                           );
   U3872 : NOR2_X1 port map( A1 => n7456, A2 => n3602, ZN => n3610);
   U3873 : NOR2_X1 port map( A1 => n5700, A2 => n3603, ZN => n3612);
   U3874 : NAND2_X1 port map( A1 => n3612, A2 => n3621, ZN => n5638);
   U3875 : INV_X1 port map( A => n5636, ZN => n3604);
   U3876 : INV_X1 port map( A => n3621, ZN => n5635);
   U3877 : NAND2_X1 port map( A1 => n3633, A2 => n5635, ZN => n3616);
   U3878 : NOR2_X1 port map( A1 => n3604, A2 => n3616, ZN => n3635);
   U3879 : INV_X1 port map( A => n3635, ZN => n3605);
   U3880 : NAND2_X1 port map( A1 => n5638, A2 => n3605, ZN => n3606);
   U3881 : AOI22_X1 port map( A1 => n5636, A2 => n3609, B1 => n3610, B2 => 
                           n3606, ZN => n3630);
   U3882 : NAND2_X1 port map( A1 => n3600, A2 => n3610, ZN => n3615);
   U3883 : NOR2_X1 port map( A1 => n3600, A2 => n3610, ZN => n3620);
   U3884 : INV_X1 port map( A => n3620, ZN => n3625);
   U3885 : NAND2_X1 port map( A1 => n3615, A2 => n3625, ZN => n3623);
   U3886 : INV_X1 port map( A => n3623, ZN => n3619);
   U3887 : NOR2_X1 port map( A1 => n5635, A2 => n3607, ZN => n3637);
   U3888 : NAND2_X1 port map( A1 => n3609, A2 => n3608, ZN => n3626);
   U3889 : AOI21_X1 port map( B1 => n3611, B2 => n3610, A => n3626, ZN => n3618
                           );
   U3890 : INV_X1 port map( A => n3612, ZN => n3622);
   U3891 : NOR2_X1 port map( A1 => n3620, A2 => n5700, ZN => n3614);
   U3892 : NAND2_X1 port map( A1 => n5635, A2 => n3613, ZN => n5699);
   U3893 : OR2_X1 port map( A1 => n3614, A2 => n5699, ZN => n3624);
   U3894 : AOI21_X2 port map( B1 => n5700, B2 => n3615, A => n3624, ZN => n7246
                           );
   U3895 : INV_X1 port map( A => n7246, ZN => n7383);
   U3896 : OAI21_X1 port map( B1 => n3616, B2 => n3622, A => n7383, ZN => n3617
                           );
   U3897 : AOI211_X1 port map( C1 => n3619, C2 => n3637, A => n3618, B => n3617
                           , ZN => n5697);
   U3898 : NAND2_X1 port map( A1 => n3630, A2 => n5697, ZN => n5629);
   U3899 : NAND2_X1 port map( A1 => n3620, A2 => n5700, ZN => n3636);
   U3900 : NOR2_X1 port map( A1 => n5699, A2 => n3636, ZN => n3631);
   U3901 : OAI21_X1 port map( B1 => n3624, B2 => n3623, A => n3558, ZN => n3638
                           );
   U3902 : INV_X1 port map( A => n3637, ZN => n3628);
   U3903 : XNOR2_X1 port map( A => n5700, B => n3625, ZN => n3627);
   U3904 : OAI22_X1 port map( A1 => n3628, A2 => n3627, B1 => n5700, B2 => 
                           n3626, ZN => n3629);
   U3905 : NOR3_X1 port map( A1 => n3631, A2 => n3638, A3 => n3629, ZN => n5631
                           );
   U3906 : NAND2_X1 port map( A1 => n3630, A2 => n5631, ZN => n5696);
   U3907 : NAND2_X1 port map( A1 => n5629, A2 => n5696, ZN => n5716);
   U3908 : INV_X1 port map( A => n3631, ZN => n3632);
   U3909 : OAI21_X1 port map( B1 => n3633, B2 => n5638, A => n3632, ZN => n3634
                           );
   U3910 : AOI211_X1 port map( C1 => n3637, C2 => n3636, A => n3635, B => n3634
                           , ZN => n5690);
   U3911 : NOR2_X1 port map( A1 => n3638, A2 => n7246, ZN => n5713);
   U3912 : AND2_X1 port map( A1 => n5690, A2 => n5713, ZN => n5688);
   U3913 : INV_X1 port map( A => n5688, ZN => n5695);
   U3914 : NOR2_X1 port map( A1 => n5716, A2 => n5695, ZN => n5679);
   U3915 : INV_X1 port map( A => n5679, ZN => n3639);
   U3916 : NOR2_X1 port map( A1 => n3639, A2 => n5708, ZN => n4349);
   U3917 : CLKBUF_X1 port map( A => n4349, Z => n7546);
   U3918 : INV_X1 port map( A => ashr_25xSHx3x, ZN => n7231);
   U3919 : NAND2_X1 port map( A1 => n7442, A2 => fromMemoryPortxLOADEDDATAx(9),
                           ZN => n3641);
   U3920 : NAND2_X1 port map( A1 => n3644, A2 => fromMemoryPortxLOADEDDATAx(22)
                           , ZN => n3640);
   U3921 : NAND2_X1 port map( A1 => n3641, A2 => n3640, ZN => n7046);
   U3922 : CLKBUF_X1 port map( A => n7046, Z => intadd_0xBx0x);
   U3923 : NAND2_X1 port map( A1 => n7442, A2 => fromMemoryPortxLOADEDDATAx(8),
                           ZN => n3643);
   U3924 : NAND2_X1 port map( A1 => n3644, A2 => fromMemoryPortxLOADEDDATAx(21)
                           , ZN => n3642);
   U3925 : NAND2_X1 port map( A1 => n3643, A2 => n3642, ZN => n7254);
   U3926 : CLKBUF_X1 port map( A => n7254, Z => n7412);
   U3927 : INV_X1 port map( A => n7412, ZN => intadd_4xBx0x);
   U3928 : NAND2_X1 port map( A1 => n7442, A2 => fromMemoryPortxLOADEDDATAx(11)
                           , ZN => n3646);
   U3929 : NAND2_X1 port map( A1 => n3644, A2 => fromMemoryPortxLOADEDDATAx(24)
                           , ZN => n3645);
   U3930 : NAND2_X1 port map( A1 => n3646, A2 => n3645, ZN => ashr_25xSHx4x);
   U3931 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(13), A2 => n5762,
                           ZN => n3648);
   U3932 : NAND2_X1 port map( A1 => n7441, A2 => n5760, ZN => n5215);
   U3933 : AND2_X1 port map( A1 => n7486, A2 => n5215, ZN => n3647);
   U3934 : OAI21_X1 port map( B1 => n5712, B2 => n3648, A => n3647, ZN => n4640
                           );
   U3935 : OR3_X1 port map( A1 => n4875, A2 => n7441, A3 => n4640, ZN => n5052)
                           ;
   U3936 : NAND2_X1 port map( A1 => n5052, A2 => fromMemoryPortxLOADEDDATAx(31)
                           , ZN => n4611);
   U3937 : INV_X1 port map( A => n5692, ZN => n4641);
   U3938 : NAND2_X1 port map( A1 => n4611, A2 => n4641, ZN => n4552);
   U3939 : NAND2_X1 port map( A1 => n4611, A2 => n7200, ZN => n3649);
   U3940 : AND2_X1 port map( A1 => n4552, A2 => n3649, ZN => add_x_26xBx27x);
   U3941 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(27), A2 => n5052,
                           ZN => add_x_26xBx7x);
   U3942 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(28), A2 => n5052,
                           ZN => add_x_26xBx8x);
   U3943 : INV_X1 port map( A => rst, ZN => n7519);
   U3944 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx26x, A2 => n7519, ZN => 
                           IF_RegsxN686);
   U3945 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx10x, A2 => n7519, ZN => 
                           IF_RegsxN670);
   U3946 : CLKBUF_X1 port map( A => n7519, Z => n7516);
   U3947 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx28x, A2 => n7516, ZN => 
                           IF_RegsxN688);
   U3948 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx12x, A2 => n7519, ZN => 
                           IF_RegsxN672);
   U3949 : CLKBUF_X1 port map( A => n7519, Z => n7505);
   U3950 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx11x, A2 => n7505, ZN => 
                           IF_RegsxN671);
   U3951 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx8x, A2 => n7505, ZN => 
                           IF_RegsxN668);
   U3952 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx22x, A2 => n7519, ZN => 
                           IF_RegsxN682);
   U3953 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx20x, A2 => n7519, ZN => 
                           IF_RegsxN680);
   U3954 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx27x, A2 => n7505, ZN => 
                           IF_RegsxN687);
   U3955 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx23x, A2 => n7505, ZN => 
                           IF_RegsxN683);
   U3956 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx15x, A2 => n7505, ZN => 
                           IF_RegsxN675);
   U3957 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx31x, A2 => n7519, ZN => 
                           IF_RegsxN691);
   U3958 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx24x, A2 => n7519, ZN => 
                           IF_RegsxN684);
   U3959 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx16x, A2 => n7519, ZN => 
                           IF_RegsxN676);
   U3960 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx30x, A2 => n7519, ZN => 
                           IF_RegsxN690);
   U3961 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx29x, A2 => n7519, ZN => 
                           IF_RegsxN689);
   U3962 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx3x, A2 => n7519, ZN => 
                           IF_RegsxN663);
   U3963 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx2x, A2 => n7505, ZN => 
                           IF_RegsxN662);
   U3964 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx7x, A2 => n7519, ZN => 
                           IF_RegsxN667);
   U3965 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx1x, A2 => n7505, ZN => 
                           IF_RegsxN661);
   U3966 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx9x, A2 => n7516, ZN => 
                           IF_RegsxN669);
   U3967 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx5x, A2 => n7519, ZN => 
                           IF_RegsxN665);
   U3968 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx21x, A2 => n7505, ZN => 
                           IF_RegsxN681);
   U3969 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx0x, A2 => n7505, ZN => 
                           IF_RegsxN660);
   U3970 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx17x, A2 => n7505, ZN => 
                           IF_RegsxN677);
   U3971 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx4x, A2 => n7505, ZN => 
                           IF_RegsxN664);
   U3972 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx14x, A2 => n7519, ZN => 
                           IF_RegsxN674);
   U3973 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx13x, A2 => n7505, ZN => 
                           IF_RegsxN673);
   U3974 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx19x, A2 => n7505, ZN => 
                           IF_RegsxN679);
   U3975 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx18x, A2 => n7519, ZN => 
                           IF_RegsxN678);
   U3976 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx6x, A2 => n7505, ZN => 
                           IF_RegsxN666);
   U3977 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx25x, A2 => n7505, ZN => 
                           IF_RegsxN685);
   U3978 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(26), A2 => n5052,
                           ZN => add_x_26xBx6x);
   U3979 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(16), A2 => 
                           fromMemoryPortxLOADEDDATAx(15), ZN => n3654);
   U3980 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(17), ZN => n6867);
   U3981 : NAND2_X1 port map( A1 => n3654, A2 => n6867, ZN => n3667);
   U3982 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(18), ZN => n6907);
   U3983 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(19), A2 => n6907
                           , ZN => n3660);
   U3984 : NOR2_X1 port map( A1 => n3667, A2 => n3660, ZN => n3938);
   U3985 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(15), ZN => n6794);
   U3986 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(16), A2 => n6867
                           , A3 => n6794, ZN => n3673);
   U3987 : NOR2_X1 port map( A1 => n3660, A2 => n3673, ZN => n3985);
   U3988 : AOI22_X1 port map( A1 => n3938, A2 => fromRegsPortxREG_FILE_16xx12x,
                           B1 => n3985, B2 => fromRegsPortxREG_FILE_18xx12x, ZN
                           => n3653);
   U3989 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(18), A2 => 
                           fromMemoryPortxLOADEDDATAx(19), ZN => n3674);
   U3990 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(17), A2 => 
                           fromMemoryPortxLOADEDDATAx(16), A3 => 
                           fromMemoryPortxLOADEDDATAx(15), ZN => n3670);
   U3991 : NOR2_X1 port map( A1 => n3674, A2 => n3670, ZN => n3986);
   U3992 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(19), ZN => n6945);
   U3993 : NAND2_X1 port map( A1 => n6907, A2 => n6945, ZN => n3671);
   U3994 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(16), A2 => 
                           fromMemoryPortxLOADEDDATAx(15), A3 => n6867, ZN => 
                           n3672);
   U3995 : NOR2_X1 port map( A1 => n3671, A2 => n3672, ZN => n4128);
   U3996 : AOI22_X1 port map( A1 => n3986, A2 => fromRegsPortxREG_FILE_31xx12x,
                           B1 => n4128, B2 => fromRegsPortxREG_FILE_03xx12x, ZN
                           => n3652);
   U3997 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(16), A2 => 
                           fromMemoryPortxLOADEDDATAx(17), A3 => n6794, ZN => 
                           n3669);
   U3998 : NOR2_X1 port map( A1 => n3671, A2 => n3669, ZN => n4058);
   U3999 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(18), A2 => n6945
                           , ZN => n3661);
   U4000 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(16), ZN => n6828);
   U4001 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(17), A2 => 
                           fromMemoryPortxLOADEDDATAx(15), A3 => n6828, ZN => 
                           n3666);
   U4002 : NOR2_X1 port map( A1 => n3661, A2 => n3666, ZN => n4204);
   U4003 : AOI22_X1 port map( A1 => n4058, A2 => fromRegsPortxREG_FILE_06xx12x,
                           B1 => n4204, B2 => fromRegsPortxREG_FILE_13xx12x, ZN
                           => n3651);
   U4004 : NOR2_X1 port map( A1 => n3660, A2 => n3670, ZN => n4091);
   U4005 : NOR2_X1 port map( A1 => n3661, A2 => n3673, ZN => n3971);
   U4006 : AOI22_X1 port map( A1 => n4091, A2 => fromRegsPortxREG_FILE_23xx12x,
                           B1 => n3971, B2 => fromRegsPortxREG_FILE_10xx12x, ZN
                           => n3650);
   U4007 : AND4_X1 port map( A1 => n3653, A2 => n3652, A3 => n3651, A4 => n3650
                           , ZN => n3682);
   U4008 : NOR2_X1 port map( A1 => n3661, A2 => n3670, ZN => n4281);
   U4009 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(17), A2 => n3654
                           , ZN => n3659);
   U4010 : NOR2_X1 port map( A1 => n3661, A2 => n3659, ZN => n4109);
   U4011 : AOI22_X1 port map( A1 => n4281, A2 => fromRegsPortxREG_FILE_15xx12x,
                           B1 => n4109, B2 => fromRegsPortxREG_FILE_12xx12x, ZN
                           => n3658);
   U4012 : NOR2_X1 port map( A1 => n3674, A2 => n3666, ZN => n3999);
   U4013 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(15), A2 => n6867
                           , A3 => n6828, ZN => n3668);
   U4014 : NOR2_X1 port map( A1 => n3668, A2 => n3660, ZN => n4063);
   U4015 : AOI22_X1 port map( A1 => n3999, A2 => fromRegsPortxREG_FILE_29xx12x,
                           B1 => n4063, B2 => fromRegsPortxREG_FILE_17xx12x, ZN
                           => n3657);
   U4016 : NOR2_X1 port map( A1 => n3661, A2 => n3667, ZN => n3980);
   U4017 : NOR2_X1 port map( A1 => n3674, A2 => n3659, ZN => n4119);
   U4018 : AOI22_X1 port map( A1 => n3980, A2 => fromRegsPortxREG_FILE_08xx12x,
                           B1 => n4119, B2 => fromRegsPortxREG_FILE_28xx12x, ZN
                           => n3656);
   U4019 : NOR2_X1 port map( A1 => n3668, A2 => n3674, ZN => n4151);
   U4020 : NOR2_X1 port map( A1 => n3671, A2 => n3659, ZN => n5354);
   U4021 : CLKBUF_X1 port map( A => n5354, Z => n5253);
   U4022 : AOI22_X1 port map( A1 => n4151, A2 => fromRegsPortxREG_FILE_25xx12x,
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx12x, ZN
                           => n3655);
   U4023 : AND4_X1 port map( A1 => n3658, A2 => n3657, A3 => n3656, A4 => n3655
                           , ZN => n3681);
   U4024 : NOR2_X1 port map( A1 => n3661, A2 => n3672, ZN => n4114);
   U4025 : CLKBUF_X1 port map( A => n4114, Z => n5338);
   U4026 : NOR2_X1 port map( A1 => n3661, A2 => n3668, ZN => n4142);
   U4027 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_11xx12x,
                           B1 => n4142, B2 => fromRegsPortxREG_FILE_09xx12x, ZN
                           => n3665);
   U4028 : NOR2_X1 port map( A1 => n3660, A2 => n3659, ZN => n3970);
   U4029 : NOR2_X1 port map( A1 => n3669, A2 => n3660, ZN => n4186);
   U4030 : AOI22_X1 port map( A1 => n3970, A2 => fromRegsPortxREG_FILE_20xx12x,
                           B1 => n4186, B2 => fromRegsPortxREG_FILE_22xx12x, ZN
                           => n3664);
   U4031 : NOR2_X1 port map( A1 => n3671, A2 => n3673, ZN => n4024);
   U4032 : NOR2_X1 port map( A1 => n3666, A2 => n3660, ZN => n5258);
   U4033 : AOI22_X1 port map( A1 => n4024, A2 => fromRegsPortxREG_FILE_02xx12x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_21xx12x, ZN
                           => n3663);
   U4034 : NOR2_X1 port map( A1 => n3660, A2 => n3672, ZN => n4089);
   U4035 : CLKBUF_X1 port map( A => n4089, Z => n5364);
   U4036 : NOR2_X1 port map( A1 => n3661, A2 => n3669, ZN => n4185);
   U4037 : AOI22_X1 port map( A1 => n5364, A2 => fromRegsPortxREG_FILE_19xx12x,
                           B1 => n4185, B2 => fromRegsPortxREG_FILE_14xx12x, ZN
                           => n3662);
   U4038 : AND4_X1 port map( A1 => n3665, A2 => n3664, A3 => n3663, A4 => n3662
                           , ZN => n3680);
   U4039 : NOR2_X1 port map( A1 => n3671, A2 => n3666, ZN => n4129);
   U4040 : NOR2_X1 port map( A1 => n3667, A2 => n3674, ZN => n4096);
   U4041 : AOI22_X1 port map( A1 => n4129, A2 => fromRegsPortxREG_FILE_05xx12x,
                           B1 => n4096, B2 => fromRegsPortxREG_FILE_24xx12x, ZN
                           => n3678);
   U4042 : NOR2_X1 port map( A1 => n3668, A2 => n3671, ZN => n4041);
   U4043 : CLKBUF_X1 port map( A => n4041, Z => n5377);
   U4044 : NOR2_X1 port map( A1 => n3674, A2 => n3669, ZN => n4072);
   U4045 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx12x,
                           B1 => n4072, B2 => fromRegsPortxREG_FILE_30xx12x, ZN
                           => n3677);
   U4046 : NOR2_X1 port map( A1 => n3671, A2 => n3670, ZN => n4090);
   U4047 : CLKBUF_X1 port map( A => n4090, Z => n5340);
   U4048 : NAND2_X1 port map( A1 => n5340, A2 => fromRegsPortxREG_FILE_07xx12x,
                           ZN => n3676);
   U4049 : NOR2_X1 port map( A1 => n3674, A2 => n3672, ZN => n4172);
   U4050 : NOR2_X1 port map( A1 => n3674, A2 => n3673, ZN => n4195);
   U4051 : AOI22_X1 port map( A1 => n4172, A2 => fromRegsPortxREG_FILE_27xx12x,
                           B1 => n4195, B2 => fromRegsPortxREG_FILE_26xx12x, ZN
                           => n3675);
   U4052 : AND4_X1 port map( A1 => n3678, A2 => n3677, A3 => n3676, A4 => n3675
                           , ZN => n3679);
   U4053 : NAND4_X1 port map( A1 => n3682, A2 => n3681, A3 => n3680, A4 => 
                           n3679, ZN => ashr_25xAx12x);
   U4054 : INV_X1 port map( A => ashr_25xAx12x, ZN => intadd_2xAx1x);
   U4055 : CLKBUF_X1 port map( A => n4129, Z => n5371);
   U4056 : CLKBUF_X1 port map( A => n3971, Z => n5366);
   U4057 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx2x, 
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx2x, ZN 
                           => n3686);
   U4058 : CLKBUF_X1 port map( A => n3970, Z => n5351);
   U4059 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx2x, 
                           B1 => n4089, B2 => fromRegsPortxREG_FILE_19xx2x, ZN 
                           => n3685);
   U4060 : CLKBUF_X1 port map( A => n4142, Z => n5337);
   U4061 : AOI22_X1 port map( A1 => n3938, A2 => fromRegsPortxREG_FILE_16xx2x, 
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx2x, ZN 
                           => n3684);
   U4062 : CLKBUF_X1 port map( A => n3980, Z => n5375);
   U4063 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx2x, 
                           B1 => n4041, B2 => fromRegsPortxREG_FILE_01xx2x, ZN 
                           => n3683);
   U4064 : AND4_X1 port map( A1 => n3686, A2 => n3685, A3 => n3684, A4 => n3683
                           , ZN => n3702);
   U4065 : CLKBUF_X1 port map( A => n4119, Z => n5374);
   U4066 : CLKBUF_X1 port map( A => n5258, Z => n5339);
   U4067 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_28xx2x, 
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx2x, ZN 
                           => n3690);
   U4068 : CLKBUF_X1 port map( A => n4058, Z => n5359);
   U4069 : CLKBUF_X1 port map( A => n4109, Z => n5353);
   U4070 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx2x, 
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_12xx2x, ZN 
                           => n3689);
   U4071 : CLKBUF_X1 port map( A => n4186, Z => n5349);
   U4072 : AOI22_X1 port map( A1 => n4024, A2 => fromRegsPortxREG_FILE_02xx2x, 
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx2x, ZN 
                           => n3688);
   U4073 : CLKBUF_X1 port map( A => n4091, Z => n5335);
   U4074 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx2x, 
                           B1 => n4114, B2 => fromRegsPortxREG_FILE_11xx2x, ZN 
                           => n3687);
   U4075 : AND4_X1 port map( A1 => n3690, A2 => n3689, A3 => n3688, A4 => n3687
                           , ZN => n3701);
   U4076 : CLKBUF_X1 port map( A => n3999, Z => n5348);
   U4077 : CLKBUF_X1 port map( A => n3985, Z => n5361);
   U4078 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx2x, 
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx2x, ZN 
                           => n3694);
   U4079 : CLKBUF_X1 port map( A => n4128, Z => n5352);
   U4080 : CLKBUF_X1 port map( A => n4185, Z => n5365);
   U4081 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx2x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx2x, ZN 
                           => n3693);
   U4082 : CLKBUF_X1 port map( A => n4072, Z => n5336);
   U4083 : CLKBUF_X1 port map( A => n4204, Z => n5363);
   U4084 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx2x, 
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx2x, ZN 
                           => n3692);
   U4085 : CLKBUF_X1 port map( A => n4281, Z => n5341);
   U4086 : CLKBUF_X1 port map( A => n4096, Z => n5373);
   U4087 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx2x, 
                           B1 => n5373, B2 => fromRegsPortxREG_FILE_24xx2x, ZN 
                           => n3691);
   U4088 : AND4_X1 port map( A1 => n3694, A2 => n3693, A3 => n3692, A4 => n3691
                           , ZN => n3700);
   U4089 : CLKBUF_X1 port map( A => n4063, Z => n5347);
   U4090 : CLKBUF_X1 port map( A => n3986, Z => n5376);
   U4091 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx2x, 
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_31xx2x, ZN 
                           => n3698);
   U4092 : CLKBUF_X1 port map( A => n4172, Z => n5350);
   U4093 : AOI22_X1 port map( A1 => n5340, A2 => fromRegsPortxREG_FILE_07xx2x, 
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx2x, ZN 
                           => n3697);
   U4094 : CLKBUF_X1 port map( A => n4151, Z => n5360);
   U4095 : CLKBUF_X1 port map( A => n4195, Z => n5362);
   U4096 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx2x, 
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx2x, ZN 
                           => n3696);
   U4097 : NAND2_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_04xx2x, 
                           ZN => n3695);
   U4098 : AND4_X1 port map( A1 => n3698, A2 => n3697, A3 => n3696, A4 => n3695
                           , ZN => n3699);
   U4099 : NAND4_X1 port map( A1 => n3702, A2 => n3701, A3 => n3700, A4 => 
                           n3699, ZN => ashr_25xAx2x);
   U4100 : INV_X1 port map( A => ashr_25xAx2x, ZN => intadd_4xAx1x);
   U4101 : AOI22_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_12xx3x, 
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx3x, ZN 
                           => n3706);
   U4102 : CLKBUF_X1 port map( A => n4024, Z => n5372);
   U4103 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx3x, 
                           B1 => n5372, B2 => fromRegsPortxREG_FILE_02xx3x, ZN 
                           => n3705);
   U4104 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx3x, 
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx3x, ZN 
                           => n3704);
   U4105 : AOI22_X1 port map( A1 => n5364, A2 => fromRegsPortxREG_FILE_19xx3x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx3x, ZN 
                           => n3703);
   U4106 : AND4_X1 port map( A1 => n3706, A2 => n3705, A3 => n3704, A4 => n3703
                           , ZN => n3724);
   U4107 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_27xx3x, 
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx3x, ZN 
                           => n3708);
   U4108 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx3x, 
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx3x, ZN 
                           => n3707);
   U4109 : NAND2_X1 port map( A1 => n3708, A2 => n3707, ZN => n3713);
   U4110 : AOI22_X1 port map( A1 => n3938, A2 => fromRegsPortxREG_FILE_16xx3x, 
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx3x, ZN 
                           => n3711);
   U4111 : NAND2_X1 port map( A1 => n5340, A2 => fromRegsPortxREG_FILE_07xx3x, 
                           ZN => n3710);
   U4112 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx3x, 
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_31xx3x, ZN 
                           => n3709);
   U4113 : NAND3_X1 port map( A1 => n3711, A2 => n3710, A3 => n3709, ZN => 
                           n3712);
   U4114 : NOR2_X1 port map( A1 => n3713, A2 => n3712, ZN => n3723);
   U4115 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx3x, 
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx3x, ZN 
                           => n3717);
   U4116 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx3x, 
                           B1 => n3971, B2 => fromRegsPortxREG_FILE_10xx3x, ZN 
                           => n3716);
   U4117 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx3x, 
                           B1 => n4041, B2 => fromRegsPortxREG_FILE_01xx3x, ZN 
                           => n3715);
   U4118 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx3x, 
                           B1 => n4114, B2 => fromRegsPortxREG_FILE_11xx3x, ZN 
                           => n3714);
   U4119 : AND4_X1 port map( A1 => n3717, A2 => n3716, A3 => n3715, A4 => n3714
                           , ZN => n3722);
   U4120 : AOI22_X1 port map( A1 => n3970, A2 => fromRegsPortxREG_FILE_20xx3x, 
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_28xx3x, ZN 
                           => n3720);
   U4121 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx3x, 
                           B1 => n5371, B2 => fromRegsPortxREG_FILE_05xx3x, ZN 
                           => n3719);
   U4122 : AOI22_X1 port map( A1 => n5373, A2 => fromRegsPortxREG_FILE_24xx3x, 
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx3x, ZN 
                           => n3718);
   U4123 : AND3_X1 port map( A1 => n3720, A2 => n3719, A3 => n3718, ZN => n3721
                           );
   U4124 : NAND4_X1 port map( A1 => n3724, A2 => n3723, A3 => n3722, A4 => 
                           n3721, ZN => ashr_25xAx3x);
   U4125 : INV_X1 port map( A => ashr_25xAx3x, ZN => intadd_4xAx2x);
   U4126 : CLKBUF_X1 port map( A => n7046, Z => n6337);
   U4127 : INV_X2 port map( A => n6337, ZN => intadd_4xBx1x);
   U4128 : CLKBUF_X2 port map( A => n5679, Z => n7547);
   U4129 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx0x, 
                           B1 => n5351, B2 => fromRegsPortxREG_FILE_20xx0x, ZN 
                           => n3727);
   U4130 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx0x, 
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx0x, ZN 
                           => n3726);
   U4131 : AOI22_X1 port map( A1 => n5364, A2 => fromRegsPortxREG_FILE_19xx0x, 
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx0x, ZN 
                           => n3725);
   U4132 : AND3_X1 port map( A1 => n3727, A2 => n3726, A3 => n3725, ZN => n3746
                           );
   U4133 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx0x, 
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_28xx0x, ZN 
                           => n3729);
   U4134 : CLKBUF_X1 port map( A => n3938, Z => n5342);
   U4135 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx0x, 
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_16xx0x, ZN 
                           => n3728);
   U4136 : NAND2_X1 port map( A1 => n3729, A2 => n3728, ZN => n3734);
   U4137 : AOI22_X1 port map( A1 => n5373, A2 => fromRegsPortxREG_FILE_24xx0x, 
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx0x, ZN 
                           => n3732);
   U4138 : NAND2_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_04xx0x, 
                           ZN => n3731);
   U4139 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx0x, 
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_31xx0x, ZN 
                           => n3730);
   U4140 : NAND3_X1 port map( A1 => n3732, A2 => n3731, A3 => n3730, ZN => 
                           n3733);
   U4141 : NOR2_X1 port map( A1 => n3734, A2 => n3733, ZN => n3745);
   U4142 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx0x, 
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx0x, ZN 
                           => n3738);
   U4143 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_11xx0x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx0x, ZN 
                           => n3737);
   U4144 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx0x, 
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx0x, ZN 
                           => n3736);
   U4145 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx0x, 
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx0x, ZN 
                           => n3735);
   U4146 : AND4_X1 port map( A1 => n3738, A2 => n3737, A3 => n3736, A4 => n3735
                           , ZN => n3744);
   U4147 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx0x, 
                           B1 => n5372, B2 => fromRegsPortxREG_FILE_02xx0x, ZN 
                           => n3742);
   U4148 : AOI22_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_12xx0x, 
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx0x, ZN 
                           => n3741);
   U4149 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx0x, 
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx0x, ZN 
                           => n3740);
   U4150 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx0x, 
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx0x, ZN 
                           => n3739);
   U4151 : AND4_X1 port map( A1 => n3742, A2 => n3741, A3 => n3740, A4 => n3739
                           , ZN => n3743);
   U4152 : NAND4_X1 port map( A1 => n3746, A2 => n3745, A3 => n3744, A4 => 
                           n3743, ZN => ashr_25xAx0x);
   U4153 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx1x, 
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_31xx1x, ZN 
                           => n3750);
   U4154 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx1x, 
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx1x, ZN 
                           => n3749);
   U4155 : AOI22_X1 port map( A1 => n5373, A2 => fromRegsPortxREG_FILE_24xx1x, 
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx1x, ZN 
                           => n3748);
   U4156 : NAND2_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_28xx1x, 
                           ZN => n3747);
   U4157 : AND4_X1 port map( A1 => n3750, A2 => n3749, A3 => n3748, A4 => n3747
                           , ZN => n3766);
   U4158 : AOI22_X1 port map( A1 => n5337, A2 => fromRegsPortxREG_FILE_09xx1x, 
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx1x, ZN 
                           => n3754);
   U4159 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx1x, 
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx1x, ZN 
                           => n3753);
   U4160 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx1x, 
                           B1 => n5335, B2 => fromRegsPortxREG_FILE_23xx1x, ZN 
                           => n3752);
   U4161 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx1x, 
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_11xx1x, ZN 
                           => n3751);
   U4162 : AND4_X1 port map( A1 => n3754, A2 => n3753, A3 => n3752, A4 => n3751
                           , ZN => n3765);
   U4163 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx1x, 
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx1x, ZN 
                           => n3758);
   U4164 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx1x, 
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx1x, ZN 
                           => n3757);
   U4165 : AOI22_X1 port map( A1 => n5372, A2 => fromRegsPortxREG_FILE_02xx1x, 
                           B1 => n5354, B2 => fromRegsPortxREG_FILE_04xx1x, ZN 
                           => n3756);
   U4166 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx1x, 
                           B1 => n5341, B2 => fromRegsPortxREG_FILE_15xx1x, ZN 
                           => n3755);
   U4167 : AND4_X1 port map( A1 => n3758, A2 => n3757, A3 => n3756, A4 => n3755
                           , ZN => n3764);
   U4168 : AOI22_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_12xx1x, 
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx1x, ZN 
                           => n3762);
   U4169 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx1x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx1x, ZN 
                           => n3761);
   U4170 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx1x, 
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_19xx1x, ZN 
                           => n3760);
   U4171 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx1x, 
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx1x, ZN 
                           => n3759);
   U4172 : AND4_X1 port map( A1 => n3762, A2 => n3761, A3 => n3760, A4 => n3759
                           , ZN => n3763);
   U4173 : NAND4_X1 port map( A1 => n3766, A2 => n3765, A3 => n3764, A4 => 
                           n3763, ZN => ashr_25xAx1x);
   U4174 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_31xx4x, 
                           B1 => n4129, B2 => fromRegsPortxREG_FILE_05xx4x, ZN 
                           => n3770);
   U4175 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx4x, 
                           B1 => n5359, B2 => fromRegsPortxREG_FILE_06xx4x, ZN 
                           => n3769);
   U4176 : AOI22_X1 port map( A1 => n5349, A2 => fromRegsPortxREG_FILE_22xx4x, 
                           B1 => n4089, B2 => fromRegsPortxREG_FILE_19xx4x, ZN 
                           => n3768);
   U4177 : AOI22_X1 port map( A1 => n4172, A2 => fromRegsPortxREG_FILE_27xx4x, 
                           B1 => n3985, B2 => fromRegsPortxREG_FILE_18xx4x, ZN 
                           => n3767);
   U4178 : AND4_X1 port map( A1 => n3770, A2 => n3769, A3 => n3768, A4 => n3767
                           , ZN => n3786);
   U4179 : AOI22_X1 port map( A1 => n4142, A2 => fromRegsPortxREG_FILE_09xx4x, 
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx4x, ZN 
                           => n3774);
   U4180 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx4x, 
                           B1 => n4109, B2 => fromRegsPortxREG_FILE_12xx4x, ZN 
                           => n3773);
   U4181 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx4x, 
                           B1 => n3970, B2 => fromRegsPortxREG_FILE_20xx4x, ZN 
                           => n3772);
   U4182 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx4x, 
                           B1 => n4119, B2 => fromRegsPortxREG_FILE_28xx4x, ZN 
                           => n3771);
   U4183 : AND4_X1 port map( A1 => n3774, A2 => n3773, A3 => n3772, A4 => n3771
                           , ZN => n3785);
   U4184 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_11xx4x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx4x, ZN 
                           => n3778);
   U4185 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx4x, 
                           B1 => n3971, B2 => fromRegsPortxREG_FILE_10xx4x, ZN 
                           => n3777);
   U4186 : AOI22_X1 port map( A1 => n4041, A2 => fromRegsPortxREG_FILE_01xx4x, 
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx4x, ZN 
                           => n3776);
   U4187 : AOI22_X1 port map( A1 => n3938, A2 => fromRegsPortxREG_FILE_16xx4x, 
                           B1 => n4281, B2 => fromRegsPortxREG_FILE_15xx4x, ZN 
                           => n3775);
   U4188 : AND4_X1 port map( A1 => n3778, A2 => n3777, A3 => n3776, A4 => n3775
                           , ZN => n3784);
   U4189 : AOI22_X1 port map( A1 => n5373, A2 => fromRegsPortxREG_FILE_24xx4x, 
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx4x, ZN 
                           => n3782);
   U4190 : NAND2_X1 port map( A1 => n4024, A2 => fromRegsPortxREG_FILE_02xx4x, 
                           ZN => n3781);
   U4191 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_13xx4x, 
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx4x, ZN 
                           => n3780);
   U4192 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx4x, 
                           B1 => n5336, B2 => fromRegsPortxREG_FILE_30xx4x, ZN 
                           => n3779);
   U4193 : AND4_X1 port map( A1 => n3782, A2 => n3781, A3 => n3780, A4 => n3779
                           , ZN => n3783);
   U4194 : NAND4_X1 port map( A1 => n3786, A2 => n3785, A3 => n3784, A4 => 
                           n3783, ZN => ashr_25xAx4x);
   U4195 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_04xx5x, 
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx5x, ZN 
                           => n3790);
   U4196 : AOI22_X1 port map( A1 => n3999, A2 => fromRegsPortxREG_FILE_29xx5x, 
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx5x, ZN 
                           => n3789);
   U4197 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx5x, 
                           B1 => n4072, B2 => fromRegsPortxREG_FILE_30xx5x, ZN 
                           => n3788);
   U4198 : NAND2_X1 port map( A1 => n4096, A2 => fromRegsPortxREG_FILE_24xx5x, 
                           ZN => n3787);
   U4199 : AND4_X1 port map( A1 => n3790, A2 => n3789, A3 => n3788, A4 => n3787
                           , ZN => n3806);
   U4200 : AOI22_X1 port map( A1 => n4058, A2 => fromRegsPortxREG_FILE_06xx5x, 
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_16xx5x, ZN 
                           => n3794);
   U4201 : AOI22_X1 port map( A1 => n3986, A2 => fromRegsPortxREG_FILE_31xx5x, 
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx5x, ZN 
                           => n3793);
   U4202 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx5x, 
                           B1 => n4119, B2 => fromRegsPortxREG_FILE_28xx5x, ZN 
                           => n3792);
   U4203 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx5x, 
                           B1 => n4109, B2 => fromRegsPortxREG_FILE_12xx5x, ZN 
                           => n3791);
   U4204 : AND4_X1 port map( A1 => n3794, A2 => n3793, A3 => n3792, A4 => n3791
                           , ZN => n3805);
   U4205 : AOI22_X1 port map( A1 => n5364, A2 => fromRegsPortxREG_FILE_19xx5x, 
                           B1 => n3971, B2 => fromRegsPortxREG_FILE_10xx5x, ZN 
                           => n3798);
   U4206 : AOI22_X1 port map( A1 => n3970, A2 => fromRegsPortxREG_FILE_20xx5x, 
                           B1 => n4185, B2 => fromRegsPortxREG_FILE_14xx5x, ZN 
                           => n3797);
   U4207 : AOI22_X1 port map( A1 => n4186, A2 => fromRegsPortxREG_FILE_22xx5x, 
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx5x, ZN 
                           => n3796);
   U4208 : AOI22_X1 port map( A1 => n4041, A2 => fromRegsPortxREG_FILE_01xx5x, 
                           B1 => n4114, B2 => fromRegsPortxREG_FILE_11xx5x, ZN 
                           => n3795);
   U4209 : AND4_X1 port map( A1 => n3798, A2 => n3797, A3 => n3796, A4 => n3795
                           , ZN => n3804);
   U4210 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx5x, 
                           B1 => n5372, B2 => fromRegsPortxREG_FILE_02xx5x, ZN 
                           => n3802);
   U4211 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx5x, 
                           B1 => n4129, B2 => fromRegsPortxREG_FILE_05xx5x, ZN 
                           => n3801);
   U4212 : AOI22_X1 port map( A1 => n4142, A2 => fromRegsPortxREG_FILE_09xx5x, 
                           B1 => n3985, B2 => fromRegsPortxREG_FILE_18xx5x, ZN 
                           => n3800);
   U4213 : AOI22_X1 port map( A1 => n3980, A2 => fromRegsPortxREG_FILE_08xx5x, 
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx5x, ZN 
                           => n3799);
   U4214 : AND4_X1 port map( A1 => n3802, A2 => n3801, A3 => n3800, A4 => n3799
                           , ZN => n3803);
   U4215 : NAND4_X1 port map( A1 => n3806, A2 => n3805, A3 => n3804, A4 => 
                           n3803, ZN => ashr_25xAx5x);
   U4216 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_28xx6x, 
                           B1 => n4089, B2 => fromRegsPortxREG_FILE_19xx6x, ZN 
                           => n3810);
   U4217 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx6x, 
                           B1 => n3985, B2 => fromRegsPortxREG_FILE_18xx6x, ZN 
                           => n3809);
   U4218 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_26xx6x, 
                           B1 => n3971, B2 => fromRegsPortxREG_FILE_10xx6x, ZN 
                           => n3808);
   U4219 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx6x, 
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx6x, ZN 
                           => n3807);
   U4220 : AND4_X1 port map( A1 => n3810, A2 => n3809, A3 => n3808, A4 => n3807
                           , ZN => n3826);
   U4221 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx6x, 
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx6x, ZN 
                           => n3814);
   U4222 : AOI22_X1 port map( A1 => n3980, A2 => fromRegsPortxREG_FILE_08xx6x, 
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx6x, ZN 
                           => n3813);
   U4223 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx6x, 
                           B1 => n5351, B2 => fromRegsPortxREG_FILE_20xx6x, ZN 
                           => n3812);
   U4224 : AOI22_X1 port map( A1 => n4090, A2 => fromRegsPortxREG_FILE_07xx6x, 
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx6x, ZN 
                           => n3811);
   U4225 : AND4_X1 port map( A1 => n3814, A2 => n3813, A3 => n3812, A4 => n3811
                           , ZN => n3825);
   U4226 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx6x, 
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx6x, ZN 
                           => n3818);
   U4227 : AOI22_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_12xx6x, 
                           B1 => n4185, B2 => fromRegsPortxREG_FILE_14xx6x, ZN 
                           => n3817);
   U4228 : AOI22_X1 port map( A1 => n3938, A2 => fromRegsPortxREG_FILE_16xx6x, 
                           B1 => n4041, B2 => fromRegsPortxREG_FILE_01xx6x, ZN 
                           => n3816);
   U4229 : AOI22_X1 port map( A1 => n5373, A2 => fromRegsPortxREG_FILE_24xx6x, 
                           B1 => n4114, B2 => fromRegsPortxREG_FILE_11xx6x, ZN 
                           => n3815);
   U4230 : AND4_X1 port map( A1 => n3818, A2 => n3817, A3 => n3816, A4 => n3815
                           , ZN => n3824);
   U4231 : AOI22_X1 port map( A1 => n3986, A2 => fromRegsPortxREG_FILE_31xx6x, 
                           B1 => n4129, B2 => fromRegsPortxREG_FILE_05xx6x, ZN 
                           => n3822);
   U4232 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx6x, 
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx6x, ZN 
                           => n3821);
   U4233 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx6x, 
                           B1 => n4072, B2 => fromRegsPortxREG_FILE_30xx6x, ZN 
                           => n3820);
   U4234 : NAND2_X1 port map( A1 => n4024, A2 => fromRegsPortxREG_FILE_02xx6x, 
                           ZN => n3819);
   U4235 : AND4_X1 port map( A1 => n3822, A2 => n3821, A3 => n3820, A4 => n3819
                           , ZN => n3823);
   U4236 : NAND4_X1 port map( A1 => n3826, A2 => n3825, A3 => n3824, A4 => 
                           n3823, ZN => ashr_25xAx6x);
   U4237 : AOI22_X1 port map( A1 => n3980, A2 => fromRegsPortxREG_FILE_08xx7x, 
                           B1 => n4128, B2 => fromRegsPortxREG_FILE_03xx7x, ZN 
                           => n3830);
   U4238 : AOI22_X1 port map( A1 => n4204, A2 => fromRegsPortxREG_FILE_13xx7x, 
                           B1 => n3985, B2 => fromRegsPortxREG_FILE_18xx7x, ZN 
                           => n3829);
   U4239 : AOI22_X1 port map( A1 => n5373, A2 => fromRegsPortxREG_FILE_24xx7x, 
                           B1 => n4185, B2 => fromRegsPortxREG_FILE_14xx7x, ZN 
                           => n3828);
   U4240 : AOI22_X1 port map( A1 => n5349, A2 => fromRegsPortxREG_FILE_22xx7x, 
                           B1 => n3971, B2 => fromRegsPortxREG_FILE_10xx7x, ZN 
                           => n3827);
   U4241 : AND4_X1 port map( A1 => n3830, A2 => n3829, A3 => n3828, A4 => n3827
                           , ZN => n3846);
   U4242 : AOI22_X1 port map( A1 => n4041, A2 => fromRegsPortxREG_FILE_01xx7x, 
                           B1 => n4109, B2 => fromRegsPortxREG_FILE_12xx7x, ZN 
                           => n3834);
   U4243 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx7x, 
                           B1 => n4119, B2 => fromRegsPortxREG_FILE_28xx7x, ZN 
                           => n3833);
   U4244 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx7x, 
                           B1 => n5351, B2 => fromRegsPortxREG_FILE_20xx7x, ZN 
                           => n3832);
   U4245 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx7x, 
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx7x, ZN 
                           => n3831);
   U4246 : AND4_X1 port map( A1 => n3834, A2 => n3833, A3 => n3832, A4 => n3831
                           , ZN => n3845);
   U4247 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx7x, 
                           B1 => n4114, B2 => fromRegsPortxREG_FILE_11xx7x, ZN 
                           => n3838);
   U4248 : AOI22_X1 port map( A1 => n3986, A2 => fromRegsPortxREG_FILE_31xx7x, 
                           B1 => n4089, B2 => fromRegsPortxREG_FILE_19xx7x, ZN 
                           => n3837);
   U4249 : AOI22_X1 port map( A1 => n3938, A2 => fromRegsPortxREG_FILE_16xx7x, 
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx7x, ZN 
                           => n3836);
   U4250 : AOI22_X1 port map( A1 => n3999, A2 => fromRegsPortxREG_FILE_29xx7x, 
                           B1 => n4281, B2 => fromRegsPortxREG_FILE_15xx7x, ZN 
                           => n3835);
   U4251 : AND4_X1 port map( A1 => n3838, A2 => n3837, A3 => n3836, A4 => n3835
                           , ZN => n3844);
   U4252 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx7x, 
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx7x, ZN 
                           => n3842);
   U4253 : AOI22_X1 port map( A1 => n4024, A2 => fromRegsPortxREG_FILE_02xx7x, 
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx7x, ZN 
                           => n3841);
   U4254 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx7x, 
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx7x, ZN 
                           => n3840);
   U4255 : NAND2_X1 port map( A1 => n4142, A2 => fromRegsPortxREG_FILE_09xx7x, 
                           ZN => n3839);
   U4256 : AND4_X1 port map( A1 => n3842, A2 => n3841, A3 => n3840, A4 => n3839
                           , ZN => n3843);
   U4257 : NAND4_X1 port map( A1 => n3846, A2 => n3845, A3 => n3844, A4 => 
                           n3843, ZN => ashr_25xAx7x);
   U4258 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx8x, 
                           B1 => n4128, B2 => fromRegsPortxREG_FILE_03xx8x, ZN 
                           => n3850);
   U4259 : AOI22_X1 port map( A1 => n4072, A2 => fromRegsPortxREG_FILE_30xx8x, 
                           B1 => n5372, B2 => fromRegsPortxREG_FILE_02xx8x, ZN 
                           => n3849);
   U4260 : AOI22_X1 port map( A1 => n4091, A2 => fromRegsPortxREG_FILE_23xx8x, 
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx8x, ZN 
                           => n3848);
   U4261 : AOI22_X1 port map( A1 => n5373, A2 => fromRegsPortxREG_FILE_24xx8x, 
                           B1 => n3985, B2 => fromRegsPortxREG_FILE_18xx8x, ZN 
                           => n3847);
   U4262 : AND4_X1 port map( A1 => n3850, A2 => n3849, A3 => n3848, A4 => n3847
                           , ZN => n3866);
   U4263 : AOI22_X1 port map( A1 => n3970, A2 => fromRegsPortxREG_FILE_20xx8x, 
                           B1 => n4109, B2 => fromRegsPortxREG_FILE_12xx8x, ZN 
                           => n3854);
   U4264 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx8x, 
                           B1 => n4186, B2 => fromRegsPortxREG_FILE_22xx8x, ZN 
                           => n3853);
   U4265 : AOI22_X1 port map( A1 => n4058, A2 => fromRegsPortxREG_FILE_06xx8x, 
                           B1 => n4119, B2 => fromRegsPortxREG_FILE_28xx8x, ZN 
                           => n3852);
   U4266 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx8x, 
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx8x, ZN 
                           => n3851);
   U4267 : AND4_X1 port map( A1 => n3854, A2 => n3853, A3 => n3852, A4 => n3851
                           , ZN => n3865);
   U4268 : AOI22_X1 port map( A1 => n4090, A2 => fromRegsPortxREG_FILE_07xx8x, 
                           B1 => n4114, B2 => fromRegsPortxREG_FILE_11xx8x, ZN 
                           => n3858);
   U4269 : AOI22_X1 port map( A1 => n5366, A2 => fromRegsPortxREG_FILE_10xx8x, 
                           B1 => n4185, B2 => fromRegsPortxREG_FILE_14xx8x, ZN 
                           => n3857);
   U4270 : AOI22_X1 port map( A1 => n3938, A2 => fromRegsPortxREG_FILE_16xx8x, 
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx8x, ZN 
                           => n3856);
   U4271 : AOI22_X1 port map( A1 => n4063, A2 => fromRegsPortxREG_FILE_17xx8x, 
                           B1 => n4281, B2 => fromRegsPortxREG_FILE_15xx8x, ZN 
                           => n3855);
   U4272 : AND4_X1 port map( A1 => n3858, A2 => n3857, A3 => n3856, A4 => n3855
                           , ZN => n3864);
   U4273 : AOI22_X1 port map( A1 => n4142, A2 => fromRegsPortxREG_FILE_09xx8x, 
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx8x, ZN 
                           => n3862);
   U4274 : AOI22_X1 port map( A1 => n3980, A2 => fromRegsPortxREG_FILE_08xx8x, 
                           B1 => n3999, B2 => fromRegsPortxREG_FILE_29xx8x, ZN 
                           => n3861);
   U4275 : NAND2_X1 port map( A1 => n5364, A2 => fromRegsPortxREG_FILE_19xx8x, 
                           ZN => n3860);
   U4276 : AOI22_X1 port map( A1 => n3986, A2 => fromRegsPortxREG_FILE_31xx8x, 
                           B1 => n4172, B2 => fromRegsPortxREG_FILE_27xx8x, ZN 
                           => n3859);
   U4277 : AND4_X1 port map( A1 => n3862, A2 => n3861, A3 => n3860, A4 => n3859
                           , ZN => n3863);
   U4278 : NAND4_X1 port map( A1 => n3866, A2 => n3865, A3 => n3864, A4 => 
                           n3863, ZN => ashr_25xAx8x);
   U4279 : AOI22_X1 port map( A1 => n3938, A2 => fromRegsPortxREG_FILE_16xx9x, 
                           B1 => n3985, B2 => fromRegsPortxREG_FILE_18xx9x, ZN 
                           => n3870);
   U4280 : AOI22_X1 port map( A1 => n4281, A2 => fromRegsPortxREG_FILE_15xx9x, 
                           B1 => n5372, B2 => fromRegsPortxREG_FILE_02xx9x, ZN 
                           => n3869);
   U4281 : AOI22_X1 port map( A1 => n4091, A2 => fromRegsPortxREG_FILE_23xx9x, 
                           B1 => n4204, B2 => fromRegsPortxREG_FILE_13xx9x, ZN 
                           => n3868);
   U4282 : AOI22_X1 port map( A1 => n3970, A2 => fromRegsPortxREG_FILE_20xx9x, 
                           B1 => n4185, B2 => fromRegsPortxREG_FILE_14xx9x, ZN 
                           => n3867);
   U4283 : AND4_X1 port map( A1 => n3870, A2 => n3869, A3 => n3868, A4 => n3867
                           , ZN => n3886);
   U4284 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx9x, 
                           B1 => n4063, B2 => fromRegsPortxREG_FILE_17xx9x, ZN 
                           => n3874);
   U4285 : AOI22_X1 port map( A1 => n4128, A2 => fromRegsPortxREG_FILE_03xx9x, 
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx9x, ZN 
                           => n3873);
   U4286 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_04xx9x, 
                           B1 => n4109, B2 => fromRegsPortxREG_FILE_12xx9x, ZN 
                           => n3872);
   U4287 : AOI22_X1 port map( A1 => n3999, A2 => fromRegsPortxREG_FILE_29xx9x, 
                           B1 => n4119, B2 => fromRegsPortxREG_FILE_28xx9x, ZN 
                           => n3871);
   U4288 : AND4_X1 port map( A1 => n3874, A2 => n3873, A3 => n3872, A4 => n3871
                           , ZN => n3885);
   U4289 : AOI22_X1 port map( A1 => n4172, A2 => fromRegsPortxREG_FILE_27xx9x, 
                           B1 => n3971, B2 => fromRegsPortxREG_FILE_10xx9x, ZN 
                           => n3878);
   U4290 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_21xx9x, 
                           B1 => n4089, B2 => fromRegsPortxREG_FILE_19xx9x, ZN 
                           => n3877);
   U4291 : AOI22_X1 port map( A1 => n3986, A2 => fromRegsPortxREG_FILE_31xx9x, 
                           B1 => n4142, B2 => fromRegsPortxREG_FILE_09xx9x, ZN 
                           => n3876);
   U4292 : AOI22_X1 port map( A1 => n4129, A2 => fromRegsPortxREG_FILE_05xx9x, 
                           B1 => n4114, B2 => fromRegsPortxREG_FILE_11xx9x, ZN 
                           => n3875);
   U4293 : AND4_X1 port map( A1 => n3878, A2 => n3877, A3 => n3876, A4 => n3875
                           , ZN => n3884);
   U4294 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx9x, 
                           B1 => n4090, B2 => fromRegsPortxREG_FILE_07xx9x, ZN 
                           => n3882);
   U4295 : AOI22_X1 port map( A1 => n4058, A2 => fromRegsPortxREG_FILE_06xx9x, 
                           B1 => n4096, B2 => fromRegsPortxREG_FILE_24xx9x, ZN 
                           => n3881);
   U4296 : AOI22_X1 port map( A1 => n3980, A2 => fromRegsPortxREG_FILE_08xx9x, 
                           B1 => n4072, B2 => fromRegsPortxREG_FILE_30xx9x, ZN 
                           => n3880);
   U4297 : NAND2_X1 port map( A1 => n4195, A2 => fromRegsPortxREG_FILE_26xx9x, 
                           ZN => n3879);
   U4298 : AND4_X1 port map( A1 => n3882, A2 => n3881, A3 => n3880, A4 => n3879
                           , ZN => n3883);
   U4299 : NAND4_X1 port map( A1 => n3886, A2 => n3885, A3 => n3884, A4 => 
                           n3883, ZN => ashr_25xAx9x);
   U4300 : AOI22_X1 port map( A1 => n3980, A2 => fromRegsPortxREG_FILE_08xx10x,
                           B1 => n4058, B2 => fromRegsPortxREG_FILE_06xx10x, ZN
                           => n3890);
   U4301 : AOI22_X1 port map( A1 => n3999, A2 => fromRegsPortxREG_FILE_29xx10x,
                           B1 => n4128, B2 => fromRegsPortxREG_FILE_03xx10x, ZN
                           => n3889);
   U4302 : AOI22_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_12xx10x,
                           B1 => n4089, B2 => fromRegsPortxREG_FILE_19xx10x, ZN
                           => n3888);
   U4303 : AOI22_X1 port map( A1 => n4195, A2 => fromRegsPortxREG_FILE_26xx10x,
                           B1 => n3985, B2 => fromRegsPortxREG_FILE_18xx10x, ZN
                           => n3887);
   U4304 : AND4_X1 port map( A1 => n3890, A2 => n3889, A3 => n3888, A4 => n3887
                           , ZN => n3906);
   U4305 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_04xx10x,
                           B1 => n3971, B2 => fromRegsPortxREG_FILE_10xx10x, ZN
                           => n3894);
   U4306 : AOI22_X1 port map( A1 => n4024, A2 => fromRegsPortxREG_FILE_02xx10x,
                           B1 => n4185, B2 => fromRegsPortxREG_FILE_14xx10x, ZN
                           => n3893);
   U4307 : AOI22_X1 port map( A1 => n4063, A2 => fromRegsPortxREG_FILE_17xx10x,
                           B1 => n4091, B2 => fromRegsPortxREG_FILE_23xx10x, ZN
                           => n3892);
   U4308 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx10x,
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx10x, ZN
                           => n3891);
   U4309 : AND4_X1 port map( A1 => n3894, A2 => n3893, A3 => n3892, A4 => n3891
                           , ZN => n3905);
   U4310 : AOI22_X1 port map( A1 => n3938, A2 => fromRegsPortxREG_FILE_16xx10x,
                           B1 => n4281, B2 => fromRegsPortxREG_FILE_15xx10x, ZN
                           => n3898);
   U4311 : AOI22_X1 port map( A1 => n3986, A2 => fromRegsPortxREG_FILE_31xx10x,
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx10x, ZN
                           => n3897);
   U4312 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_28xx10x,
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx10x, ZN
                           => n3896);
   U4313 : AOI22_X1 port map( A1 => n3970, A2 => fromRegsPortxREG_FILE_20xx10x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx10x, ZN
                           => n3895);
   U4314 : AND4_X1 port map( A1 => n3898, A2 => n3897, A3 => n3896, A4 => n3895
                           , ZN => n3904);
   U4315 : AOI22_X1 port map( A1 => n4072, A2 => fromRegsPortxREG_FILE_30xx10x,
                           B1 => n4090, B2 => fromRegsPortxREG_FILE_07xx10x, ZN
                           => n3902);
   U4316 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx10x,
                           B1 => n4096, B2 => fromRegsPortxREG_FILE_24xx10x, ZN
                           => n3901);
   U4317 : NAND2_X1 port map( A1 => n4041, A2 => fromRegsPortxREG_FILE_01xx10x,
                           ZN => n3900);
   U4318 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_11xx10x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx10x, ZN
                           => n3899);
   U4319 : AND4_X1 port map( A1 => n3902, A2 => n3901, A3 => n3900, A4 => n3899
                           , ZN => n3903);
   U4320 : NAND4_X1 port map( A1 => n3906, A2 => n3905, A3 => n3904, A4 => 
                           n3903, ZN => ashr_25xAx10x);
   U4321 : AOI22_X1 port map( A1 => n3986, A2 => fromRegsPortxREG_FILE_31xx11x,
                           B1 => n4128, B2 => fromRegsPortxREG_FILE_03xx11x, ZN
                           => n3910);
   U4322 : AOI22_X1 port map( A1 => n4072, A2 => fromRegsPortxREG_FILE_30xx11x,
                           B1 => n3985, B2 => fromRegsPortxREG_FILE_18xx11x, ZN
                           => n3909);
   U4323 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx11x,
                           B1 => n3971, B2 => fromRegsPortxREG_FILE_10xx11x, ZN
                           => n3908);
   U4324 : AOI22_X1 port map( A1 => n3999, A2 => fromRegsPortxREG_FILE_29xx11x,
                           B1 => n4089, B2 => fromRegsPortxREG_FILE_19xx11x, ZN
                           => n3907);
   U4325 : AND4_X1 port map( A1 => n3910, A2 => n3909, A3 => n3908, A4 => n3907
                           , ZN => n3926);
   U4326 : AOI22_X1 port map( A1 => n3970, A2 => fromRegsPortxREG_FILE_20xx11x,
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx11x, ZN
                           => n3914);
   U4327 : AOI22_X1 port map( A1 => n4024, A2 => fromRegsPortxREG_FILE_02xx11x,
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx11x, ZN
                           => n3913);
   U4328 : AOI22_X1 port map( A1 => n3980, A2 => fromRegsPortxREG_FILE_08xx11x,
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx11x, ZN
                           => n3912);
   U4329 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx11x,
                           B1 => n4063, B2 => fromRegsPortxREG_FILE_17xx11x, ZN
                           => n3911);
   U4330 : AND4_X1 port map( A1 => n3914, A2 => n3913, A3 => n3912, A4 => n3911
                           , ZN => n3925);
   U4331 : AOI22_X1 port map( A1 => n4041, A2 => fromRegsPortxREG_FILE_01xx11x,
                           B1 => n4091, B2 => fromRegsPortxREG_FILE_23xx11x, ZN
                           => n3918);
   U4332 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_11xx11x,
                           B1 => n4185, B2 => fromRegsPortxREG_FILE_14xx11x, ZN
                           => n3917);
   U4333 : AOI22_X1 port map( A1 => n3938, A2 => fromRegsPortxREG_FILE_16xx11x,
                           B1 => n4281, B2 => fromRegsPortxREG_FILE_15xx11x, ZN
                           => n3916);
   U4334 : AOI22_X1 port map( A1 => n4090, A2 => fromRegsPortxREG_FILE_07xx11x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx11x, ZN
                           => n3915);
   U4335 : AND4_X1 port map( A1 => n3918, A2 => n3917, A3 => n3916, A4 => n3915
                           , ZN => n3924);
   U4336 : AOI22_X1 port map( A1 => n4119, A2 => fromRegsPortxREG_FILE_28xx11x,
                           B1 => n4096, B2 => fromRegsPortxREG_FILE_24xx11x, ZN
                           => n3922);
   U4337 : AOI22_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_12xx11x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx11x, ZN
                           => n3921);
   U4338 : AOI22_X1 port map( A1 => n4058, A2 => fromRegsPortxREG_FILE_06xx11x,
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx11x, ZN
                           => n3920);
   U4339 : NAND2_X1 port map( A1 => n4204, A2 => fromRegsPortxREG_FILE_13xx11x,
                           ZN => n3919);
   U4340 : AND4_X1 port map( A1 => n3922, A2 => n3921, A3 => n3920, A4 => n3919
                           , ZN => n3923);
   U4341 : NAND4_X1 port map( A1 => n3926, A2 => n3925, A3 => n3924, A4 => 
                           n3923, ZN => ashr_25xAx11x);
   U4342 : AOI22_X1 port map( A1 => n3999, A2 => fromRegsPortxREG_FILE_29xx13x,
                           B1 => n3985, B2 => fromRegsPortxREG_FILE_18xx13x, ZN
                           => n3930);
   U4343 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx13x,
                           B1 => n5372, B2 => fromRegsPortxREG_FILE_02xx13x, ZN
                           => n3929);
   U4344 : AOI22_X1 port map( A1 => n4058, A2 => fromRegsPortxREG_FILE_06xx13x,
                           B1 => n4089, B2 => fromRegsPortxREG_FILE_19xx13x, ZN
                           => n3928);
   U4345 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx13x,
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx13x, ZN
                           => n3927);
   U4346 : AND4_X1 port map( A1 => n3930, A2 => n3929, A3 => n3928, A4 => n3927
                           , ZN => n3949);
   U4347 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_04xx13x,
                           B1 => n4186, B2 => fromRegsPortxREG_FILE_22xx13x, ZN
                           => n3932);
   U4348 : AOI22_X1 port map( A1 => n4119, A2 => fromRegsPortxREG_FILE_28xx13x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_21xx13x, ZN
                           => n3931);
   U4349 : NAND2_X1 port map( A1 => n3932, A2 => n3931, ZN => n3937);
   U4350 : AOI22_X1 port map( A1 => n3980, A2 => fromRegsPortxREG_FILE_08xx13x,
                           B1 => n4109, B2 => fromRegsPortxREG_FILE_12xx13x, ZN
                           => n3935);
   U4351 : NAND2_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_11xx13x,
                           ZN => n3934);
   U4352 : AOI22_X1 port map( A1 => n4172, A2 => fromRegsPortxREG_FILE_27xx13x,
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx13x, ZN
                           => n3933);
   U4353 : NAND3_X1 port map( A1 => n3935, A2 => n3934, A3 => n3933, ZN => 
                           n3936);
   U4354 : NOR2_X1 port map( A1 => n3937, A2 => n3936, ZN => n3948);
   U4355 : AOI22_X1 port map( A1 => n3938, A2 => fromRegsPortxREG_FILE_16xx13x,
                           B1 => n4185, B2 => fromRegsPortxREG_FILE_14xx13x, ZN
                           => n3942);
   U4356 : AOI22_X1 port map( A1 => n3986, A2 => fromRegsPortxREG_FILE_31xx13x,
                           B1 => n3971, B2 => fromRegsPortxREG_FILE_10xx13x, ZN
                           => n3941);
   U4357 : AOI22_X1 port map( A1 => n4063, A2 => fromRegsPortxREG_FILE_17xx13x,
                           B1 => n4091, B2 => fromRegsPortxREG_FILE_23xx13x, ZN
                           => n3940);
   U4358 : AOI22_X1 port map( A1 => n5373, A2 => fromRegsPortxREG_FILE_24xx13x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx13x, ZN
                           => n3939);
   U4359 : AND4_X1 port map( A1 => n3942, A2 => n3941, A3 => n3940, A4 => n3939
                           , ZN => n3947);
   U4360 : AOI22_X1 port map( A1 => n4128, A2 => fromRegsPortxREG_FILE_03xx13x,
                           B1 => n3970, B2 => fromRegsPortxREG_FILE_20xx13x, ZN
                           => n3945);
   U4361 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx13x,
                           B1 => n4090, B2 => fromRegsPortxREG_FILE_07xx13x, ZN
                           => n3944);
   U4362 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx13x,
                           B1 => n4129, B2 => fromRegsPortxREG_FILE_05xx13x, ZN
                           => n3943);
   U4363 : AND3_X1 port map( A1 => n3945, A2 => n3944, A3 => n3943, ZN => n3946
                           );
   U4364 : NAND4_X1 port map( A1 => n3949, A2 => n3948, A3 => n3947, A4 => 
                           n3946, ZN => ashr_25xAx13x);
   U4365 : AOI22_X1 port map( A1 => n4063, A2 => fromRegsPortxREG_FILE_17xx14x,
                           B1 => n4096, B2 => fromRegsPortxREG_FILE_24xx14x, ZN
                           => n3953);
   U4366 : AOI22_X1 port map( A1 => n3980, A2 => fromRegsPortxREG_FILE_08xx14x,
                           B1 => n4172, B2 => fromRegsPortxREG_FILE_27xx14x, ZN
                           => n3952);
   U4367 : NAND2_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_12xx14x,
                           ZN => n3951);
   U4368 : AOI22_X1 port map( A1 => n4151, A2 => fromRegsPortxREG_FILE_25xx14x,
                           B1 => n5336, B2 => fromRegsPortxREG_FILE_30xx14x, ZN
                           => n3950);
   U4369 : AND4_X1 port map( A1 => n3953, A2 => n3952, A3 => n3951, A4 => n3950
                           , ZN => n3969);
   U4370 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_26xx14x,
                           B1 => n4185, B2 => fromRegsPortxREG_FILE_14xx14x, ZN
                           => n3957);
   U4371 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_21xx14x,
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx14x, ZN
                           => n3956);
   U4372 : AOI22_X1 port map( A1 => n4128, A2 => fromRegsPortxREG_FILE_03xx14x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx14x, ZN
                           => n3955);
   U4373 : AOI22_X1 port map( A1 => n3999, A2 => fromRegsPortxREG_FILE_29xx14x,
                           B1 => n4091, B2 => fromRegsPortxREG_FILE_23xx14x, ZN
                           => n3954);
   U4374 : AND4_X1 port map( A1 => n3957, A2 => n3956, A3 => n3955, A4 => n3954
                           , ZN => n3968);
   U4375 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx14x,
                           B1 => n4114, B2 => fromRegsPortxREG_FILE_11xx14x, ZN
                           => n3961);
   U4376 : AOI22_X1 port map( A1 => n3986, A2 => fromRegsPortxREG_FILE_31xx14x,
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx14x, ZN
                           => n3960);
   U4377 : AOI22_X1 port map( A1 => n4119, A2 => fromRegsPortxREG_FILE_28xx14x,
                           B1 => n4186, B2 => fromRegsPortxREG_FILE_22xx14x, ZN
                           => n3959);
   U4378 : AOI22_X1 port map( A1 => n4058, A2 => fromRegsPortxREG_FILE_06xx14x,
                           B1 => n4281, B2 => fromRegsPortxREG_FILE_15xx14x, ZN
                           => n3958);
   U4379 : AND4_X1 port map( A1 => n3961, A2 => n3960, A3 => n3959, A4 => n3958
                           , ZN => n3967);
   U4380 : AOI22_X1 port map( A1 => n3970, A2 => fromRegsPortxREG_FILE_20xx14x,
                           B1 => n4129, B2 => fromRegsPortxREG_FILE_05xx14x, ZN
                           => n3965);
   U4381 : AOI22_X1 port map( A1 => n5364, A2 => fromRegsPortxREG_FILE_19xx14x,
                           B1 => n3985, B2 => fromRegsPortxREG_FILE_18xx14x, ZN
                           => n3964);
   U4382 : AOI22_X1 port map( A1 => n4024, A2 => fromRegsPortxREG_FILE_02xx14x,
                           B1 => n3971, B2 => fromRegsPortxREG_FILE_10xx14x, ZN
                           => n3963);
   U4383 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx14x,
                           B1 => n4090, B2 => fromRegsPortxREG_FILE_07xx14x, ZN
                           => n3962);
   U4384 : AND4_X1 port map( A1 => n3965, A2 => n3964, A3 => n3963, A4 => n3962
                           , ZN => n3966);
   U4385 : NAND4_X1 port map( A1 => n3969, A2 => n3968, A3 => n3967, A4 => 
                           n3966, ZN => ashr_25xAx14x);
   U4386 : AOI22_X1 port map( A1 => n4058, A2 => fromRegsPortxREG_FILE_06xx15x,
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx15x, ZN
                           => n3975);
   U4387 : AOI22_X1 port map( A1 => n3970, A2 => fromRegsPortxREG_FILE_20xx15x,
                           B1 => n4185, B2 => fromRegsPortxREG_FILE_14xx15x, ZN
                           => n3974);
   U4388 : AOI22_X1 port map( A1 => n5364, A2 => fromRegsPortxREG_FILE_19xx15x,
                           B1 => n3971, B2 => fromRegsPortxREG_FILE_10xx15x, ZN
                           => n3973);
   U4389 : AOI22_X1 port map( A1 => n4128, A2 => fromRegsPortxREG_FILE_03xx15x,
                           B1 => n4091, B2 => fromRegsPortxREG_FILE_23xx15x, ZN
                           => n3972);
   U4390 : AND4_X1 port map( A1 => n3975, A2 => n3974, A3 => n3973, A4 => n3972
                           , ZN => n3994);
   U4391 : AOI22_X1 port map( A1 => n4024, A2 => fromRegsPortxREG_FILE_02xx15x,
                           B1 => n4114, B2 => fromRegsPortxREG_FILE_11xx15x, ZN
                           => n3979);
   U4392 : AOI22_X1 port map( A1 => n4119, A2 => fromRegsPortxREG_FILE_28xx15x,
                           B1 => n4186, B2 => fromRegsPortxREG_FILE_22xx15x, ZN
                           => n3978);
   U4393 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_21xx15x,
                           B1 => n4109, B2 => fromRegsPortxREG_FILE_12xx15x, ZN
                           => n3977);
   U4394 : AOI22_X1 port map( A1 => n4063, A2 => fromRegsPortxREG_FILE_17xx15x,
                           B1 => n4142, B2 => fromRegsPortxREG_FILE_09xx15x, ZN
                           => n3976);
   U4395 : AND4_X1 port map( A1 => n3979, A2 => n3978, A3 => n3977, A4 => n3976
                           , ZN => n3993);
   U4396 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx15x,
                           B1 => n4172, B2 => fromRegsPortxREG_FILE_27xx15x, ZN
                           => n3984);
   U4397 : AOI22_X1 port map( A1 => n4129, A2 => fromRegsPortxREG_FILE_05xx15x,
                           B1 => n4195, B2 => fromRegsPortxREG_FILE_26xx15x, ZN
                           => n3983);
   U4398 : AOI22_X1 port map( A1 => n4151, A2 => fromRegsPortxREG_FILE_25xx15x,
                           B1 => n3999, B2 => fromRegsPortxREG_FILE_29xx15x, ZN
                           => n3982);
   U4399 : NAND2_X1 port map( A1 => n3980, A2 => fromRegsPortxREG_FILE_08xx15x,
                           ZN => n3981);
   U4400 : AND4_X1 port map( A1 => n3984, A2 => n3983, A3 => n3982, A4 => n3981
                           , ZN => n3992);
   U4401 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_04xx15x,
                           B1 => n3985, B2 => fromRegsPortxREG_FILE_18xx15x, ZN
                           => n3990);
   U4402 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx15x,
                           B1 => n4090, B2 => fromRegsPortxREG_FILE_07xx15x, ZN
                           => n3989);
   U4403 : AOI22_X1 port map( A1 => n4281, A2 => fromRegsPortxREG_FILE_15xx15x,
                           B1 => n4096, B2 => fromRegsPortxREG_FILE_24xx15x, ZN
                           => n3988);
   U4404 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx15x,
                           B1 => n3986, B2 => fromRegsPortxREG_FILE_31xx15x, ZN
                           => n3987);
   U4405 : AND4_X1 port map( A1 => n3990, A2 => n3989, A3 => n3988, A4 => n3987
                           , ZN => n3991);
   U4406 : NAND4_X1 port map( A1 => n3994, A2 => n3993, A3 => n3992, A4 => 
                           n3991, ZN => ashr_25xAx15x);
   U4407 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx16x,
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx16x, ZN
                           => n3998);
   U4408 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx16x,
                           B1 => n4109, B2 => fromRegsPortxREG_FILE_12xx16x, ZN
                           => n3997);
   U4409 : AOI22_X1 port map( A1 => n4281, A2 => fromRegsPortxREG_FILE_15xx16x,
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_28xx16x, ZN
                           => n3996);
   U4410 : AOI22_X1 port map( A1 => n4058, A2 => fromRegsPortxREG_FILE_06xx16x,
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx16x, ZN
                           => n3995);
   U4411 : AND4_X1 port map( A1 => n3998, A2 => n3997, A3 => n3996, A4 => n3995
                           , ZN => n4015);
   U4412 : AOI22_X1 port map( A1 => n4186, A2 => fromRegsPortxREG_FILE_22xx16x,
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx16x, ZN
                           => n4003);
   U4413 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_11xx16x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx16x, ZN
                           => n4002);
   U4414 : AOI22_X1 port map( A1 => n3999, A2 => fromRegsPortxREG_FILE_29xx16x,
                           B1 => n4041, B2 => fromRegsPortxREG_FILE_01xx16x, ZN
                           => n4001);
   U4415 : AOI22_X1 port map( A1 => n4129, A2 => fromRegsPortxREG_FILE_05xx16x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx16x, ZN
                           => n4000);
   U4416 : AND4_X1 port map( A1 => n4003, A2 => n4002, A3 => n4001, A4 => n4000
                           , ZN => n4014);
   U4417 : AOI22_X1 port map( A1 => n4128, A2 => fromRegsPortxREG_FILE_03xx16x,
                           B1 => n4024, B2 => fromRegsPortxREG_FILE_02xx16x, ZN
                           => n4007);
   U4418 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx16x,
                           B1 => n4089, B2 => fromRegsPortxREG_FILE_19xx16x, ZN
                           => n4006);
   U4419 : AOI22_X1 port map( A1 => n4063, A2 => fromRegsPortxREG_FILE_17xx16x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx16x, ZN
                           => n4005);
   U4420 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_31xx16x,
                           B1 => n4096, B2 => fromRegsPortxREG_FILE_24xx16x, ZN
                           => n4004);
   U4421 : AND4_X1 port map( A1 => n4007, A2 => n4006, A3 => n4005, A4 => n4004
                           , ZN => n4013);
   U4422 : AOI22_X1 port map( A1 => n4091, A2 => fromRegsPortxREG_FILE_23xx16x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx16x, ZN
                           => n4011);
   U4423 : AOI22_X1 port map( A1 => n4090, A2 => fromRegsPortxREG_FILE_07xx16x,
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx16x, ZN
                           => n4010);
   U4424 : AOI22_X1 port map( A1 => n4151, A2 => fromRegsPortxREG_FILE_25xx16x,
                           B1 => n4072, B2 => fromRegsPortxREG_FILE_30xx16x, ZN
                           => n4009);
   U4425 : NAND2_X1 port map( A1 => n5365, A2 => fromRegsPortxREG_FILE_14xx16x,
                           ZN => n4008);
   U4426 : AND4_X1 port map( A1 => n4011, A2 => n4010, A3 => n4009, A4 => n4008
                           , ZN => n4012);
   U4427 : NAND4_X1 port map( A1 => n4015, A2 => n4014, A3 => n4013, A4 => 
                           n4012, ZN => ashr_25xAx16x);
   U4428 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx17x,
                           B1 => n4089, B2 => fromRegsPortxREG_FILE_19xx17x, ZN
                           => n4019);
   U4429 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx17x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx17x, ZN
                           => n4018);
   U4430 : AOI22_X1 port map( A1 => n4195, A2 => fromRegsPortxREG_FILE_26xx17x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx17x, ZN
                           => n4017);
   U4431 : AOI22_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_12xx17x,
                           B1 => n4204, B2 => fromRegsPortxREG_FILE_13xx17x, ZN
                           => n4016);
   U4432 : AND4_X1 port map( A1 => n4019, A2 => n4018, A3 => n4017, A4 => n4016
                           , ZN => n4036);
   U4433 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx17x,
                           B1 => n4063, B2 => fromRegsPortxREG_FILE_17xx17x, ZN
                           => n4023);
   U4434 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_31xx17x,
                           B1 => n5354, B2 => fromRegsPortxREG_FILE_04xx17x, ZN
                           => n4022);
   U4435 : AOI22_X1 port map( A1 => n4041, A2 => fromRegsPortxREG_FILE_01xx17x,
                           B1 => n5351, B2 => fromRegsPortxREG_FILE_20xx17x, ZN
                           => n4021);
   U4436 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx17x,
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_28xx17x, ZN
                           => n4020);
   U4437 : AND4_X1 port map( A1 => n4023, A2 => n4022, A3 => n4021, A4 => n4020
                           , ZN => n4035);
   U4438 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx17x,
                           B1 => n4114, B2 => fromRegsPortxREG_FILE_11xx17x, ZN
                           => n4028);
   U4439 : AOI22_X1 port map( A1 => n4024, A2 => fromRegsPortxREG_FILE_02xx17x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_21xx17x, ZN
                           => n4027);
   U4440 : AOI22_X1 port map( A1 => n4172, A2 => fromRegsPortxREG_FILE_27xx17x,
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx17x, ZN
                           => n4026);
   U4441 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx17x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx17x, ZN
                           => n4025);
   U4442 : AND4_X1 port map( A1 => n4028, A2 => n4027, A3 => n4026, A4 => n4025
                           , ZN => n4034);
   U4443 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx17x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx17x, ZN
                           => n4032);
   U4444 : AOI22_X1 port map( A1 => n4151, A2 => fromRegsPortxREG_FILE_25xx17x,
                           B1 => n4096, B2 => fromRegsPortxREG_FILE_24xx17x, ZN
                           => n4031);
   U4445 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx17x,
                           B1 => n4072, B2 => fromRegsPortxREG_FILE_30xx17x, ZN
                           => n4030);
   U4446 : NAND2_X1 port map( A1 => n5366, A2 => fromRegsPortxREG_FILE_10xx17x,
                           ZN => n4029);
   U4447 : AND4_X1 port map( A1 => n4032, A2 => n4031, A3 => n4030, A4 => n4029
                           , ZN => n4033);
   U4448 : NAND4_X1 port map( A1 => n4036, A2 => n4035, A3 => n4034, A4 => 
                           n4033, ZN => ashr_25xAx17x);
   U4449 : AOI22_X1 port map( A1 => n4151, A2 => fromRegsPortxREG_FILE_25xx18x,
                           B1 => n4129, B2 => fromRegsPortxREG_FILE_05xx18x, ZN
                           => n4040);
   U4450 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_31xx18x,
                           B1 => n5372, B2 => fromRegsPortxREG_FILE_02xx18x, ZN
                           => n4039);
   U4451 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx18x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx18x, ZN
                           => n4038);
   U4452 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx18x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx18x, ZN
                           => n4037);
   U4453 : AND4_X1 port map( A1 => n4040, A2 => n4039, A3 => n4038, A4 => n4037
                           , ZN => n4057);
   U4454 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx18x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_12xx18x, ZN
                           => n4045);
   U4455 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx18x,
                           B1 => n4186, B2 => fromRegsPortxREG_FILE_22xx18x, ZN
                           => n4044);
   U4456 : AOI22_X1 port map( A1 => n4041, A2 => fromRegsPortxREG_FILE_01xx18x,
                           B1 => n5351, B2 => fromRegsPortxREG_FILE_20xx18x, ZN
                           => n4043);
   U4457 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx18x,
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_28xx18x, ZN
                           => n4042);
   U4458 : AND4_X1 port map( A1 => n4045, A2 => n4044, A3 => n4043, A4 => n4042
                           , ZN => n4056);
   U4459 : AOI22_X1 port map( A1 => n5364, A2 => fromRegsPortxREG_FILE_19xx18x,
                           B1 => n4204, B2 => fromRegsPortxREG_FILE_13xx18x, ZN
                           => n4049);
   U4460 : AOI22_X1 port map( A1 => n4072, A2 => fromRegsPortxREG_FILE_30xx18x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx18x, ZN
                           => n4048);
   U4461 : AOI22_X1 port map( A1 => n4090, A2 => fromRegsPortxREG_FILE_07xx18x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_21xx18x, ZN
                           => n4047);
   U4462 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx18x,
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_11xx18x, ZN
                           => n4046);
   U4463 : AND4_X1 port map( A1 => n4049, A2 => n4048, A3 => n4047, A4 => n4046
                           , ZN => n4055);
   U4464 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx18x,
                           B1 => n4096, B2 => fromRegsPortxREG_FILE_24xx18x, ZN
                           => n4053);
   U4465 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_04xx18x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx18x, ZN
                           => n4052);
   U4466 : AOI22_X1 port map( A1 => n4142, A2 => fromRegsPortxREG_FILE_09xx18x,
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx18x, ZN
                           => n4051);
   U4467 : NAND2_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx18x,
                           ZN => n4050);
   U4468 : AND4_X1 port map( A1 => n4053, A2 => n4052, A3 => n4051, A4 => n4050
                           , ZN => n4054);
   U4469 : NAND4_X1 port map( A1 => n4057, A2 => n4056, A3 => n4055, A4 => 
                           n4054, ZN => ashr_25xAx18x);
   U4470 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx19x,
                           B1 => n4058, B2 => fromRegsPortxREG_FILE_06xx19x, ZN
                           => n4062);
   U4471 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_31xx19x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx19x, ZN
                           => n4061);
   U4472 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_11xx19x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx19x, ZN
                           => n4060);
   U4473 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_28xx19x,
                           B1 => n4089, B2 => fromRegsPortxREG_FILE_19xx19x, ZN
                           => n4059);
   U4474 : AND4_X1 port map( A1 => n4062, A2 => n4061, A3 => n4060, A4 => n4059
                           , ZN => n4080);
   U4475 : AOI22_X1 port map( A1 => n4172, A2 => fromRegsPortxREG_FILE_27xx19x,
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx19x, ZN
                           => n4067);
   U4476 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx19x,
                           B1 => n4063, B2 => fromRegsPortxREG_FILE_17xx19x, ZN
                           => n4066);
   U4477 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx19x,
                           B1 => n5354, B2 => fromRegsPortxREG_FILE_04xx19x, ZN
                           => n4065);
   U4478 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx19x,
                           B1 => n4109, B2 => fromRegsPortxREG_FILE_12xx19x, ZN
                           => n4064);
   U4479 : AND4_X1 port map( A1 => n4067, A2 => n4066, A3 => n4065, A4 => n4064
                           , ZN => n4079);
   U4480 : AOI22_X1 port map( A1 => n5372, A2 => fromRegsPortxREG_FILE_02xx19x,
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx19x, ZN
                           => n4071);
   U4481 : AOI22_X1 port map( A1 => n4195, A2 => fromRegsPortxREG_FILE_26xx19x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx19x, ZN
                           => n4070);
   U4482 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx19x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_21xx19x, ZN
                           => n4069);
   U4483 : AOI22_X1 port map( A1 => n4151, A2 => fromRegsPortxREG_FILE_25xx19x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx19x, ZN
                           => n4068);
   U4484 : AND4_X1 port map( A1 => n4071, A2 => n4070, A3 => n4069, A4 => n4068
                           , ZN => n4078);
   U4485 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx19x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx19x, ZN
                           => n4076);
   U4486 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx19x,
                           B1 => n4096, B2 => fromRegsPortxREG_FILE_24xx19x, ZN
                           => n4075);
   U4487 : NAND2_X1 port map( A1 => n4091, A2 => fromRegsPortxREG_FILE_23xx19x,
                           ZN => n4074);
   U4488 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx19x,
                           B1 => n4072, B2 => fromRegsPortxREG_FILE_30xx19x, ZN
                           => n4073);
   U4489 : AND4_X1 port map( A1 => n4076, A2 => n4075, A3 => n4074, A4 => n4073
                           , ZN => n4077);
   U4490 : NAND4_X1 port map( A1 => n4080, A2 => n4079, A3 => n4078, A4 => 
                           n4077, ZN => ashr_25xAx19x);
   U4491 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx20x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx20x, ZN
                           => n4084);
   U4492 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx20x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx20x, ZN
                           => n4083);
   U4493 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx20x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx20x, ZN
                           => n4082);
   U4494 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx20x,
                           B1 => n4204, B2 => fromRegsPortxREG_FILE_13xx20x, ZN
                           => n4081);
   U4495 : AND4_X1 port map( A1 => n4084, A2 => n4083, A3 => n4082, A4 => n4081
                           , ZN => n4104);
   U4496 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx20x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_16xx20x, ZN
                           => n4088);
   U4497 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx20x,
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx20x, ZN
                           => n4087);
   U4498 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx20x,
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_28xx20x, ZN
                           => n4086);
   U4499 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx20x,
                           B1 => n4109, B2 => fromRegsPortxREG_FILE_12xx20x, ZN
                           => n4085);
   U4500 : AND4_X1 port map( A1 => n4088, A2 => n4087, A3 => n4086, A4 => n4085
                           , ZN => n4103);
   U4501 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx20x,
                           B1 => n4114, B2 => fromRegsPortxREG_FILE_11xx20x, ZN
                           => n4095);
   U4502 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx20x,
                           B1 => n4089, B2 => fromRegsPortxREG_FILE_19xx20x, ZN
                           => n4094);
   U4503 : AOI22_X1 port map( A1 => n4090, A2 => fromRegsPortxREG_FILE_07xx20x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_21xx20x, ZN
                           => n4093);
   U4504 : AOI22_X1 port map( A1 => n4151, A2 => fromRegsPortxREG_FILE_25xx20x,
                           B1 => n4091, B2 => fromRegsPortxREG_FILE_23xx20x, ZN
                           => n4092);
   U4505 : AND4_X1 port map( A1 => n4095, A2 => n4094, A3 => n4093, A4 => n4092
                           , ZN => n4102);
   U4506 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_31xx20x,
                           B1 => n4096, B2 => fromRegsPortxREG_FILE_24xx20x, ZN
                           => n4100);
   U4507 : AOI22_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_04xx20x,
                           B1 => n4195, B2 => fromRegsPortxREG_FILE_26xx20x, ZN
                           => n4099);
   U4508 : AOI22_X1 port map( A1 => n5372, A2 => fromRegsPortxREG_FILE_02xx20x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx20x, ZN
                           => n4098);
   U4509 : NAND2_X1 port map( A1 => n4142, A2 => fromRegsPortxREG_FILE_09xx20x,
                           ZN => n4097);
   U4510 : AND4_X1 port map( A1 => n4100, A2 => n4099, A3 => n4098, A4 => n4097
                           , ZN => n4101);
   U4511 : NAND4_X1 port map( A1 => n4104, A2 => n4103, A3 => n4102, A4 => 
                           n4101, ZN => ashr_25xAx20x);
   U4512 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx21x,
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_31xx21x, ZN
                           => n4108);
   U4513 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx21x,
                           B1 => n5336, B2 => fromRegsPortxREG_FILE_30xx21x, ZN
                           => n4107);
   U4514 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx21x,
                           B1 => n4195, B2 => fromRegsPortxREG_FILE_26xx21x, ZN
                           => n4106);
   U4515 : NAND2_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_27xx21x,
                           ZN => n4105);
   U4516 : AND4_X1 port map( A1 => n4108, A2 => n4107, A3 => n4106, A4 => n4105
                           , ZN => n4127);
   U4517 : AOI22_X1 port map( A1 => n5372, A2 => fromRegsPortxREG_FILE_02xx21x,
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx21x, ZN
                           => n4113);
   U4518 : AOI22_X1 port map( A1 => n5373, A2 => fromRegsPortxREG_FILE_24xx21x,
                           B1 => n4186, B2 => fromRegsPortxREG_FILE_22xx21x, ZN
                           => n4112);
   U4519 : AOI22_X1 port map( A1 => n4142, A2 => fromRegsPortxREG_FILE_09xx21x,
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx21x, ZN
                           => n4111);
   U4520 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx21x,
                           B1 => n4109, B2 => fromRegsPortxREG_FILE_12xx21x, ZN
                           => n4110);
   U4521 : AND4_X1 port map( A1 => n4113, A2 => n4112, A3 => n4111, A4 => n4110
                           , ZN => n4126);
   U4522 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx21x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_19xx21x, ZN
                           => n4118);
   U4523 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx21x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx21x, ZN
                           => n4117);
   U4524 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx21x,
                           B1 => n5335, B2 => fromRegsPortxREG_FILE_23xx21x, ZN
                           => n4116);
   U4525 : AOI22_X1 port map( A1 => n4151, A2 => fromRegsPortxREG_FILE_25xx21x,
                           B1 => n4114, B2 => fromRegsPortxREG_FILE_11xx21x, ZN
                           => n4115);
   U4526 : AND4_X1 port map( A1 => n4118, A2 => n4117, A3 => n4116, A4 => n4115
                           , ZN => n4125);
   U4527 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx21x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx21x, ZN
                           => n4123);
   U4528 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx21x,
                           B1 => n4204, B2 => fromRegsPortxREG_FILE_13xx21x, ZN
                           => n4122);
   U4529 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx21x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx21x, ZN
                           => n4121);
   U4530 : AOI22_X1 port map( A1 => n4119, A2 => fromRegsPortxREG_FILE_28xx21x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx21x, ZN
                           => n4120);
   U4531 : AND4_X1 port map( A1 => n4123, A2 => n4122, A3 => n4121, A4 => n4120
                           , ZN => n4124);
   U4532 : NAND4_X1 port map( A1 => n4127, A2 => n4126, A3 => n4125, A4 => 
                           n4124, ZN => ashr_25xAx21x);
   U4533 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx22x,
                           B1 => n4128, B2 => fromRegsPortxREG_FILE_03xx22x, ZN
                           => n4133);
   U4534 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx22x,
                           B1 => n4129, B2 => fromRegsPortxREG_FILE_05xx22x, ZN
                           => n4132);
   U4535 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx22x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_19xx22x, ZN
                           => n4131);
   U4536 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx22x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx22x, ZN
                           => n4130);
   U4537 : AND4_X1 port map( A1 => n4133, A2 => n4132, A3 => n4131, A4 => n4130
                           , ZN => n4150);
   U4538 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx22x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_16xx22x, ZN
                           => n4137);
   U4539 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx22x,
                           B1 => n5347, B2 => fromRegsPortxREG_FILE_17xx22x, ZN
                           => n4136);
   U4540 : AOI22_X1 port map( A1 => n4151, A2 => fromRegsPortxREG_FILE_25xx22x,
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_28xx22x, ZN
                           => n4135);
   U4541 : AOI22_X1 port map( A1 => n5372, A2 => fromRegsPortxREG_FILE_02xx22x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_12xx22x, ZN
                           => n4134);
   U4542 : AND4_X1 port map( A1 => n4137, A2 => n4136, A3 => n4135, A4 => n4134
                           , ZN => n4149);
   U4543 : AOI22_X1 port map( A1 => n4186, A2 => fromRegsPortxREG_FILE_22xx22x,
                           B1 => n4204, B2 => fromRegsPortxREG_FILE_13xx22x, ZN
                           => n4141);
   U4544 : AOI22_X1 port map( A1 => n5373, A2 => fromRegsPortxREG_FILE_24xx22x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx22x, ZN
                           => n4140);
   U4545 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx22x,
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx22x, ZN
                           => n4139);
   U4546 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_11xx22x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx22x, ZN
                           => n4138);
   U4547 : AND4_X1 port map( A1 => n4141, A2 => n4140, A3 => n4139, A4 => n4138
                           , ZN => n4148);
   U4548 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_31xx22x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx22x, ZN
                           => n4146);
   U4549 : AOI22_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_04xx22x,
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx22x, ZN
                           => n4145);
   U4550 : AOI22_X1 port map( A1 => n4142, A2 => fromRegsPortxREG_FILE_09xx22x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx22x, ZN
                           => n4144);
   U4551 : NAND2_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx22x,
                           ZN => n4143);
   U4552 : AND4_X1 port map( A1 => n4146, A2 => n4145, A3 => n4144, A4 => n4143
                           , ZN => n4147);
   U4553 : NAND4_X1 port map( A1 => n4150, A2 => n4149, A3 => n4148, A4 => 
                           n4147, ZN => ashr_25xAx22x);
   U4554 : AOI22_X1 port map( A1 => n4151, A2 => fromRegsPortxREG_FILE_25xx23x,
                           B1 => n5359, B2 => fromRegsPortxREG_FILE_06xx23x, ZN
                           => n4155);
   U4555 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx23x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx23x, ZN
                           => n4154);
   U4556 : AOI22_X1 port map( A1 => n5337, A2 => fromRegsPortxREG_FILE_09xx23x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_19xx23x, ZN
                           => n4153);
   U4557 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx23x,
                           B1 => n4204, B2 => fromRegsPortxREG_FILE_13xx23x, ZN
                           => n4152);
   U4558 : AND4_X1 port map( A1 => n4155, A2 => n4154, A3 => n4153, A4 => n4152
                           , ZN => n4171);
   U4559 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx23x,
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx23x, ZN
                           => n4159);
   U4560 : AOI22_X1 port map( A1 => n4172, A2 => fromRegsPortxREG_FILE_27xx23x,
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx23x, ZN
                           => n4158);
   U4561 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx23x,
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx23x, ZN
                           => n4157);
   U4562 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_31xx23x,
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_28xx23x, ZN
                           => n4156);
   U4563 : AND4_X1 port map( A1 => n4159, A2 => n4158, A3 => n4157, A4 => n4156
                           , ZN => n4170);
   U4564 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx23x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx23x, ZN
                           => n4163);
   U4565 : AOI22_X1 port map( A1 => n5372, A2 => fromRegsPortxREG_FILE_02xx23x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx23x, ZN
                           => n4162);
   U4566 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx23x,
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_01xx23x, ZN
                           => n4161);
   U4567 : AOI22_X1 port map( A1 => n5340, A2 => fromRegsPortxREG_FILE_07xx23x,
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_11xx23x, ZN
                           => n4160);
   U4568 : AND4_X1 port map( A1 => n4163, A2 => n4162, A3 => n4161, A4 => n4160
                           , ZN => n4169);
   U4569 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx23x,
                           B1 => n5373, B2 => fromRegsPortxREG_FILE_24xx23x, ZN
                           => n4167);
   U4570 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx23x,
                           B1 => n4195, B2 => fromRegsPortxREG_FILE_26xx23x, ZN
                           => n4166);
   U4571 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx23x,
                           B1 => n5348, B2 => fromRegsPortxREG_FILE_29xx23x, ZN
                           => n4165);
   U4572 : NAND2_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_12xx23x,
                           ZN => n4164);
   U4573 : AND4_X1 port map( A1 => n4167, A2 => n4166, A3 => n4165, A4 => n4164
                           , ZN => n4168);
   U4574 : NAND4_X1 port map( A1 => n4171, A2 => n4170, A3 => n4169, A4 => 
                           n4168, ZN => ashr_25xAx23x);
   U4575 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx24x,
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_31xx24x, ZN
                           => n4176);
   U4576 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_04xx24x,
                           B1 => n4195, B2 => fromRegsPortxREG_FILE_26xx24x, ZN
                           => n4175);
   U4577 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx24x,
                           B1 => n4172, B2 => fromRegsPortxREG_FILE_27xx24x, ZN
                           => n4174);
   U4578 : NAND2_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx24x,
                           ZN => n4173);
   U4579 : AND4_X1 port map( A1 => n4176, A2 => n4175, A3 => n4174, A4 => n4173
                           , ZN => n4194);
   U4580 : AOI22_X1 port map( A1 => n5361, A2 => fromRegsPortxREG_FILE_18xx24x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx24x, ZN
                           => n4180);
   U4581 : AOI22_X1 port map( A1 => n5372, A2 => fromRegsPortxREG_FILE_02xx24x,
                           B1 => n4204, B2 => fromRegsPortxREG_FILE_13xx24x, ZN
                           => n4179);
   U4582 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx24x,
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_01xx24x, ZN
                           => n4178);
   U4583 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx24x,
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_11xx24x, ZN
                           => n4177);
   U4584 : AND4_X1 port map( A1 => n4180, A2 => n4179, A3 => n4178, A4 => n4177
                           , ZN => n4193);
   U4585 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx24x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx24x, ZN
                           => n4184);
   U4586 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx24x,
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_28xx24x, ZN
                           => n4183);
   U4587 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx24x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_12xx24x, ZN
                           => n4182);
   U4588 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx24x,
                           B1 => n5335, B2 => fromRegsPortxREG_FILE_23xx24x, ZN
                           => n4181);
   U4589 : AND4_X1 port map( A1 => n4184, A2 => n4183, A3 => n4182, A4 => n4181
                           , ZN => n4192);
   U4590 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx24x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx24x, ZN
                           => n4190);
   U4591 : AOI22_X1 port map( A1 => n5258, A2 => fromRegsPortxREG_FILE_21xx24x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_19xx24x, ZN
                           => n4189);
   U4592 : AOI22_X1 port map( A1 => n4186, A2 => fromRegsPortxREG_FILE_22xx24x,
                           B1 => n4185, B2 => fromRegsPortxREG_FILE_14xx24x, ZN
                           => n4188);
   U4593 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx24x,
                           B1 => n5373, B2 => fromRegsPortxREG_FILE_24xx24x, ZN
                           => n4187);
   U4594 : AND4_X1 port map( A1 => n4190, A2 => n4189, A3 => n4188, A4 => n4187
                           , ZN => n4191);
   U4595 : NAND4_X1 port map( A1 => n4194, A2 => n4193, A3 => n4192, A4 => 
                           n4191, ZN => ashr_25xAx24x);
   U4596 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx25x,
                           B1 => n5373, B2 => fromRegsPortxREG_FILE_24xx25x, ZN
                           => n4199);
   U4597 : AOI22_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_12xx25x,
                           B1 => n4195, B2 => fromRegsPortxREG_FILE_26xx25x, ZN
                           => n4198);
   U4598 : NAND2_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx25x,
                           ZN => n4197);
   U4599 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_31xx25x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx25x, ZN
                           => n4196);
   U4600 : AND4_X1 port map( A1 => n4199, A2 => n4198, A3 => n4197, A4 => n4196
                           , ZN => n4216);
   U4601 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx25x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_21xx25x, ZN
                           => n4203);
   U4602 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx25x,
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx25x, ZN
                           => n4202);
   U4603 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx25x,
                           B1 => n5351, B2 => fromRegsPortxREG_FILE_20xx25x, ZN
                           => n4201);
   U4604 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx25x,
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx25x, ZN
                           => n4200);
   U4605 : AND4_X1 port map( A1 => n4203, A2 => n4202, A3 => n4201, A4 => n4200
                           , ZN => n4215);
   U4606 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx25x,
                           B1 => n4204, B2 => fromRegsPortxREG_FILE_13xx25x, ZN
                           => n4208);
   U4607 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx25x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx25x, ZN
                           => n4207);
   U4608 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx25x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx25x, ZN
                           => n4206);
   U4609 : AOI22_X1 port map( A1 => n5372, A2 => fromRegsPortxREG_FILE_02xx25x,
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_11xx25x, ZN
                           => n4205);
   U4610 : AND4_X1 port map( A1 => n4208, A2 => n4207, A3 => n4206, A4 => n4205
                           , ZN => n4214);
   U4611 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_28xx25x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx25x, ZN
                           => n4212);
   U4612 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx25x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_19xx25x, ZN
                           => n4211);
   U4613 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx25x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx25x, ZN
                           => n4210);
   U4614 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx25x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx25x, ZN
                           => n4209);
   U4615 : AND4_X1 port map( A1 => n4212, A2 => n4211, A3 => n4210, A4 => n4209
                           , ZN => n4213);
   U4616 : NAND4_X1 port map( A1 => n4216, A2 => n4215, A3 => n4214, A4 => 
                           n4213, ZN => ashr_25xAx25x);
   U4617 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx27x,
                           B1 => n5371, B2 => fromRegsPortxREG_FILE_05xx27x, ZN
                           => n4220);
   U4618 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx27x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_03xx27x, ZN
                           => n4219);
   U4619 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx27x,
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx27x, ZN
                           => n4218);
   U4620 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_28xx27x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx27x, ZN
                           => n4217);
   U4621 : AND4_X1 port map( A1 => n4220, A2 => n4219, A3 => n4218, A4 => n4217
                           , ZN => n4236);
   U4622 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx27x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_21xx27x, ZN
                           => n4224);
   U4623 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx27x,
                           B1 => n5347, B2 => fromRegsPortxREG_FILE_17xx27x, ZN
                           => n4223);
   U4624 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx27x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_12xx27x, ZN
                           => n4222);
   U4625 : AOI22_X1 port map( A1 => n5372, A2 => fromRegsPortxREG_FILE_02xx27x,
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx27x, ZN
                           => n4221);
   U4626 : AND4_X1 port map( A1 => n4224, A2 => n4223, A3 => n4222, A4 => n4221
                           , ZN => n4235);
   U4627 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx27x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx27x, ZN
                           => n4228);
   U4628 : AOI22_X1 port map( A1 => n5340, A2 => fromRegsPortxREG_FILE_07xx27x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx27x, ZN
                           => n4227);
   U4629 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_11xx27x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx27x, ZN
                           => n4226);
   U4630 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx27x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_19xx27x, ZN
                           => n4225);
   U4631 : AND4_X1 port map( A1 => n4228, A2 => n4227, A3 => n4226, A4 => n4225
                           , ZN => n4234);
   U4632 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx27x,
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_31xx27x, ZN
                           => n4232);
   U4633 : AOI22_X1 port map( A1 => n5349, A2 => fromRegsPortxREG_FILE_22xx27x,
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx27x, ZN
                           => n4231);
   U4634 : AOI22_X1 port map( A1 => n5373, A2 => fromRegsPortxREG_FILE_24xx27x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx27x, ZN
                           => n4230);
   U4635 : NAND2_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx27x,
                           ZN => n4229);
   U4636 : AND4_X1 port map( A1 => n4232, A2 => n4231, A3 => n4230, A4 => n4229
                           , ZN => n4233);
   U4637 : NAND4_X1 port map( A1 => n4236, A2 => n4235, A3 => n4234, A4 => 
                           n4233, ZN => ashr_25xAx27x);
   U4638 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx28x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_12xx28x, ZN
                           => n4240);
   U4639 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx28x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_21xx28x, ZN
                           => n4239);
   U4640 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx28x,
                           B1 => n5351, B2 => fromRegsPortxREG_FILE_20xx28x, ZN
                           => n4238);
   U4641 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx28x,
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_04xx28x, ZN
                           => n4237);
   U4642 : AND4_X1 port map( A1 => n4240, A2 => n4239, A3 => n4238, A4 => n4237
                           , ZN => n4256);
   U4643 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx28x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx28x, ZN
                           => n4244);
   U4644 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_13xx28x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx28x, ZN
                           => n4243);
   U4645 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx28x,
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_11xx28x, ZN
                           => n4242);
   U4646 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx28x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx28x, ZN
                           => n4241);
   U4647 : AND4_X1 port map( A1 => n4244, A2 => n4243, A3 => n4242, A4 => n4241
                           , ZN => n4255);
   U4648 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx28x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx28x, ZN
                           => n4248);
   U4649 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx28x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_19xx28x, ZN
                           => n4247);
   U4650 : AOI22_X1 port map( A1 => n5349, A2 => fromRegsPortxREG_FILE_22xx28x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx28x, ZN
                           => n4246);
   U4651 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx28x,
                           B1 => n5373, B2 => fromRegsPortxREG_FILE_24xx28x, ZN
                           => n4245);
   U4652 : AND4_X1 port map( A1 => n4248, A2 => n4247, A3 => n4246, A4 => n4245
                           , ZN => n4254);
   U4653 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx28x,
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_31xx28x, ZN
                           => n4252);
   U4654 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_28xx28x,
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx28x, ZN
                           => n4251);
   U4655 : AOI22_X1 port map( A1 => n5372, A2 => fromRegsPortxREG_FILE_02xx28x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx28x, ZN
                           => n4250);
   U4656 : NAND2_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx28x,
                           ZN => n4249);
   U4657 : AND4_X1 port map( A1 => n4252, A2 => n4251, A3 => n4250, A4 => n4249
                           , ZN => n4253);
   U4658 : NAND4_X1 port map( A1 => n4256, A2 => n4255, A3 => n4254, A4 => 
                           n4253, ZN => ashr_25xAx28x);
   U4659 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx29x,
                           B1 => n5373, B2 => fromRegsPortxREG_FILE_24xx29x, ZN
                           => n4260);
   U4660 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx29x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx29x, ZN
                           => n4259);
   U4661 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx29x,
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx29x, ZN
                           => n4258);
   U4662 : NAND2_X1 port map( A1 => n5337, A2 => fromRegsPortxREG_FILE_09xx29x,
                           ZN => n4257);
   U4663 : AND4_X1 port map( A1 => n4260, A2 => n4259, A3 => n4258, A4 => n4257
                           , ZN => n4276);
   U4664 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx29x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx29x, ZN
                           => n4264);
   U4665 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_31xx29x,
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx29x, ZN
                           => n4263);
   U4666 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx29x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx29x, ZN
                           => n4262);
   U4667 : AOI22_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_04xx29x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_19xx29x, ZN
                           => n4261);
   U4668 : AND4_X1 port map( A1 => n4264, A2 => n4263, A3 => n4262, A4 => n4261
                           , ZN => n4275);
   U4669 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx29x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_21xx29x, ZN
                           => n4268);
   U4670 : AOI22_X1 port map( A1 => n5340, A2 => fromRegsPortxREG_FILE_07xx29x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_12xx29x, ZN
                           => n4267);
   U4671 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx29x,
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_28xx29x, ZN
                           => n4266);
   U4672 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx29x,
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_11xx29x, ZN
                           => n4265);
   U4673 : AND4_X1 port map( A1 => n4268, A2 => n4267, A3 => n4266, A4 => n4265
                           , ZN => n4274);
   U4674 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx29x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_03xx29x, ZN
                           => n4272);
   U4675 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx29x,
                           B1 => n5372, B2 => fromRegsPortxREG_FILE_02xx29x, ZN
                           => n4271);
   U4676 : AOI22_X1 port map( A1 => n5349, A2 => fromRegsPortxREG_FILE_22xx29x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx29x, ZN
                           => n4270);
   U4677 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx29x,
                           B1 => n5371, B2 => fromRegsPortxREG_FILE_05xx29x, ZN
                           => n4269);
   U4678 : AND4_X1 port map( A1 => n4272, A2 => n4271, A3 => n4270, A4 => n4269
                           , ZN => n4273);
   U4679 : NAND4_X1 port map( A1 => n4276, A2 => n4275, A3 => n4274, A4 => 
                           n4273, ZN => ashr_25xAx29x);
   U4680 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_27xx30x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx30x, ZN
                           => n4280);
   U4681 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx30x,
                           B1 => n5371, B2 => fromRegsPortxREG_FILE_05xx30x, ZN
                           => n4279);
   U4682 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_28xx30x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_19xx30x, ZN
                           => n4278);
   U4683 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx30x,
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx30x, ZN
                           => n4277);
   U4684 : AND4_X1 port map( A1 => n4280, A2 => n4279, A3 => n4278, A4 => n4277
                           , ZN => n4297);
   U4685 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx30x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx30x, ZN
                           => n4285);
   U4686 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx30x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx30x, ZN
                           => n4284);
   U4687 : AOI22_X1 port map( A1 => n4281, A2 => fromRegsPortxREG_FILE_15xx30x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx30x, ZN
                           => n4283);
   U4688 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx30x,
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_01xx30x, ZN
                           => n4282);
   U4689 : AND4_X1 port map( A1 => n4285, A2 => n4284, A3 => n4283, A4 => n4282
                           , ZN => n4296);
   U4690 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx30x,
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx30x, ZN
                           => n4289);
   U4691 : AOI22_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_04xx30x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_12xx30x, ZN
                           => n4288);
   U4692 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx30x,
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx30x, ZN
                           => n4287);
   U4693 : AOI22_X1 port map( A1 => n5340, A2 => fromRegsPortxREG_FILE_07xx30x,
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_11xx30x, ZN
                           => n4286);
   U4694 : AND4_X1 port map( A1 => n4289, A2 => n4288, A3 => n4287, A4 => n4286
                           , ZN => n4295);
   U4695 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_31xx30x,
                           B1 => n5372, B2 => fromRegsPortxREG_FILE_02xx30x, ZN
                           => n4293);
   U4696 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx30x,
                           B1 => n5373, B2 => fromRegsPortxREG_FILE_24xx30x, ZN
                           => n4292);
   U4697 : NAND2_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx30x,
                           ZN => n4291);
   U4698 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx30x,
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx30x, ZN
                           => n4290);
   U4699 : AND4_X1 port map( A1 => n4293, A2 => n4292, A3 => n4291, A4 => n4290
                           , ZN => n4294);
   U4700 : NAND4_X1 port map( A1 => n4297, A2 => n4296, A3 => n4295, A4 => 
                           n4294, ZN => ashr_25xAx30x);
   U4701 : NOR2_X1 port map( A1 => toRegsPortxDSTxx0x, A2 => n7536, ZN => n4299
                           );
   U4702 : NAND3_X1 port map( A1 => n7530, A2 => n7533, A3 => 
                           toRegsPortxDSTxx3x, ZN => n7510);
   U4703 : OR2_X1 port map( A1 => n7535, A2 => n7510, ZN => n7495);
   U4704 : INV_X1 port map( A => n7495, ZN => n4298);
   U4705 : AOI21_X1 port map( B1 => n4299, B2 => n4298, A => rst, ZN => n4300);
   U4706 : INV_X1 port map( A => n4300, ZN => IF_RegsxN698);
   U4707 : NAND2_X1 port map( A1 => n5692, A2 => fromMemoryPortxLOADEDDATAx(30)
                           , ZN => n4301);
   U4708 : NAND2_X1 port map( A1 => n4611, A2 => n4301, ZN => add_x_26xBx30x);
   U4709 : INV_X1 port map( A => add_x_26xBx30x, ZN => intadd_3xBx2x);
   U4710 : OR2_X1 port map( A1 => n5629, A2 => n5631, ZN => n5687);
   U4711 : NOR2_X1 port map( A1 => n5687, A2 => n5713, ZN => n5691);
   U4712 : NAND2_X1 port map( A1 => n5691, A2 => n6045, ZN => n5673);
   U4713 : CLKBUF_X1 port map( A => n5673, Z => n5678);
   U4714 : AOI21_X1 port map( B1 => n5691, B2 => n6043, A => n7546, ZN => n5676
                           );
   U4715 : CLKBUF_X1 port map( A => n5676, Z => n5674);
   U4716 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(21), ZN => n5734);
   U4717 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(20), A2 => n5734
                           , ZN => n4306);
   U4718 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4306,
                           ZN => n5182);
   U4719 : CLKBUF_X1 port map( A => n5182, Z => n5276);
   U4720 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(20), ZN => n6982);
   U4721 : NAND2_X1 port map( A1 => n5734, A2 => n6982, ZN => n4315);
   U4722 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4315,
                           ZN => n5120);
   U4723 : CLKBUF_X1 port map( A => n5120, Z => n5280);
   U4724 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx30x,
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_24xx30x, ZN
                           => n4305);
   U4725 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(23), A2 => 
                           fromMemoryPortxLOADEDDATAx(22), ZN => n4326);
   U4726 : NOR2_X1 port map( A1 => n4326, A2 => n4306, ZN => n5053);
   U4727 : CLKBUF_X1 port map( A => n5053, Z => n5278);
   U4728 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(21), A2 => n6982
                           , ZN => n4307);
   U4729 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4307,
                           ZN => n5087);
   U4730 : CLKBUF_X1 port map( A => n5087, Z => n5277);
   U4731 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx30x,
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx30x, ZN
                           => n4304);
   U4732 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(21), A2 => 
                           fromMemoryPortxLOADEDDATAx(20), ZN => n4308);
   U4733 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4308,
                           ZN => n5119);
   U4734 : CLKBUF_X1 port map( A => n5119, Z => n5279);
   U4735 : NOR2_X1 port map( A1 => n4326, A2 => n4315, ZN => n5085);
   U4736 : CLKBUF_X1 port map( A => n5085, Z => n5281);
   U4737 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_27xx30x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx30x, ZN
                           => n4303);
   U4738 : NOR2_X1 port map( A1 => n4326, A2 => n4307, ZN => n5086);
   U4739 : CLKBUF_X1 port map( A => n5086, Z => n5275);
   U4740 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(22), ZN => n7027);
   U4741 : NOR3_X1 port map( A1 => n5275, A2 => n7027, A3 => n5734, ZN => n5054
                           );
   U4742 : CLKBUF_X1 port map( A => n5054, Z => n5282);
   U4743 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx30x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx30x, ZN
                           => n4302);
   U4744 : NAND4_X1 port map( A1 => n4305, A2 => n4304, A3 => n4303, A4 => 
                           n4302, ZN => n4314);
   U4745 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(23), ZN => n7065);
   U4746 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n7065
                           , ZN => n4335);
   U4747 : NOR2_X1 port map( A1 => n4306, A2 => n4335, ZN => n5158);
   U4748 : CLKBUF_X1 port map( A => n5158, Z => n5288);
   U4749 : NAND2_X1 port map( A1 => n7065, A2 => n7027, ZN => n4322);
   U4750 : NOR2_X1 port map( A1 => n4306, A2 => n4322, ZN => n5125);
   U4751 : CLKBUF_X1 port map( A => n5125, Z => n5292);
   U4752 : AOI22_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx30x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx30x, ZN
                           => n4312);
   U4753 : NOR2_X1 port map( A1 => n4308, A2 => n4335, ZN => n5126);
   U4754 : CLKBUF_X1 port map( A => n5126, Z => n5289);
   U4755 : NOR2_X1 port map( A1 => n4307, A2 => n4322, ZN => n5093);
   U4756 : CLKBUF_X1 port map( A => n5093, Z => n5293);
   U4757 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx30x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx30x, ZN
                           => n4311);
   U4758 : NOR2_X1 port map( A1 => n4315, A2 => n4335, ZN => n5092);
   U4759 : CLKBUF_X1 port map( A => n5092, Z => n5290);
   U4760 : NOR2_X1 port map( A1 => n4307, A2 => n4335, ZN => n5287);
   U4761 : CLKBUF_X1 port map( A => n5287, Z => n5224);
   U4762 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx30x,
                           B1 => n5224, B2 => fromRegsPortxREG_FILE_22xx30x, ZN
                           => n4310);
   U4763 : NOR2_X1 port map( A1 => n4308, A2 => n4322, ZN => n5187);
   U4764 : CLKBUF_X1 port map( A => n5187, Z => n5291);
   U4765 : NAND2_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_19xx30x,
                           ZN => n4309);
   U4766 : NAND4_X1 port map( A1 => n4312, A2 => n4311, A3 => n4310, A4 => 
                           n4309, ZN => n4313);
   U4767 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4314
                           , A => n4313, ZN => n4321);
   U4768 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(24), ZN => n5200);
   U4769 : CLKBUF_X1 port map( A => n5200, Z => n5758);
   U4770 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(21), A2 => n5758
                           , A3 => n6982, ZN => n4331);
   U4771 : NOR2_X1 port map( A1 => n4326, A2 => n4331, ZN => n5102);
   U4772 : CLKBUF_X1 port map( A => n5102, Z => n5302);
   U4773 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(21), A2 => 
                           fromMemoryPortxLOADEDDATAx(24), ZN => n4327);
   U4774 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(20), A2 => n4327
                           , ZN => n4334);
   U4775 : INV_X1 port map( A => n4334, ZN => n5194);
   U4776 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx30x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx30x, ZN
                           => n4320);
   U4777 : NAND2_X1 port map( A1 => n6982, A2 => n4327, ZN => n4332);
   U4778 : INV_X1 port map( A => n4332, ZN => n5301);
   U4779 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4331,
                           ZN => n5165);
   U4780 : CLKBUF_X1 port map( A => n5165, Z => n5300);
   U4781 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(21), A2 => 
                           fromMemoryPortxLOADEDDATAx(20), A3 => n5758, ZN => 
                           n4325);
   U4782 : NOR2_X1 port map( A1 => n4326, A2 => n4325, ZN => n5100);
   U4783 : CLKBUF_X1 port map( A => n5100, Z => n5305);
   U4784 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx30x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx30x, ZN
                           => n4317);
   U4785 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4325,
                           ZN => n5101);
   U4786 : CLKBUF_X1 port map( A => n5101, Z => n5303);
   U4787 : NOR2_X1 port map( A1 => n4315, A2 => n4322, ZN => n5065);
   U4788 : CLKBUF_X1 port map( A => n5065, Z => n5309);
   U4789 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_11xx30x,
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx30x, ZN
                           => n4316);
   U4790 : NAND2_X1 port map( A1 => n4317, A2 => n4316, ZN => n4318);
   U4791 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx30x, B2 => n5301,
                           A => n4318, ZN => n4319);
   U4792 : OAI211_X1 port map( C1 => n4321, C2 => n5758, A => n4320, B => n4319
                           , ZN => n4329);
   U4793 : NOR2_X1 port map( A1 => n4322, A2 => n4331, ZN => n4867);
   U4794 : CLKBUF_X1 port map( A => n4867, Z => n5326);
   U4795 : INV_X1 port map( A => n4322, ZN => n4323);
   U4796 : NAND2_X1 port map( A1 => n4323, A2 => n4327, ZN => n4340);
   U4797 : INV_X1 port map( A => n4340, ZN => n4324);
   U4798 : NOR2_X1 port map( A1 => n5326, A2 => n4324, ZN => n5047);
   U4799 : CLKBUF_X1 port map( A => n5047, Z => n5331);
   U4800 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(23), A2 => n4325,
                           ZN => n4330);
   U4801 : AOI21_X1 port map( B1 => n4327, B2 => n4326, A => n4330, ZN => n4328
                           );
   U4802 : AND2_X1 port map( A1 => n5331, A2 => n4328, ZN => n5238);
   U4803 : NAND2_X1 port map( A1 => n4329, A2 => n5238, ZN => n4346);
   U4804 : INV_X1 port map( A => n4330, ZN => n4333);
   U4805 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4333,
                           ZN => n5142);
   U4806 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4332,
                           ZN => n5039);
   U4807 : CLKBUF_X1 port map( A => n5039, Z => n5321);
   U4808 : AOI22_X1 port map( A1 => n5142, A2 => fromRegsPortxREG_FILE_03xx30x,
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx30x, ZN
                           => n4339);
   U4809 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4334,
                           ZN => n5203);
   U4810 : CLKBUF_X1 port map( A => n5203, Z => n5318);
   U4811 : NOR2_X1 port map( A1 => n4335, A2 => n4331, ZN => n5141);
   U4812 : CLKBUF_X1 port map( A => n5141, Z => n5316);
   U4813 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx30x,
                           B1 => n5316, B2 => fromRegsPortxREG_FILE_06xx30x, ZN
                           => n4338);
   U4814 : NOR2_X1 port map( A1 => n4335, A2 => n4332, ZN => n5073);
   U4815 : CLKBUF_X1 port map( A => n5073, Z => n5317);
   U4816 : NOR2_X1 port map( A1 => n7027, A2 => n4333, ZN => n5140);
   U4817 : CLKBUF_X1 port map( A => n5140, Z => n5319);
   U4818 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx30x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx30x, ZN
                           => n4337);
   U4819 : NOR2_X1 port map( A1 => n4335, A2 => n4334, ZN => n5010);
   U4820 : CLKBUF_X1 port map( A => n5010, Z => n5320);
   U4821 : NAND2_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_05xx30x,
                           ZN => n4336);
   U4822 : NAND4_X1 port map( A1 => n4339, A2 => n4338, A3 => n4337, A4 => 
                           n4336, ZN => n4344);
   U4823 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx30x,
                           ZN => n4342);
   U4824 : NOR2_X1 port map( A1 => n6982, A2 => n4340, ZN => n5327);
   U4825 : CLKBUF_X1 port map( A => n5327, Z => n5244);
   U4826 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx30x, A2 => n5244,
                           ZN => n4341);
   U4827 : NAND2_X1 port map( A1 => n4342, A2 => n4341, ZN => n4343);
   U4828 : AOI21_X1 port map( B1 => n4344, B2 => n5331, A => n4343, ZN => n4345
                           );
   U4829 : NAND2_X1 port map( A1 => n4346, A2 => n4345, ZN => n7317);
   U4830 : INV_X1 port map( A => n7317, ZN => n7483);
   U4831 : OAI22_X1 port map( A1 => n5678, A2 => intadd_3xBx2x, B1 => n5674, B2
                           => n7483, ZN => n4347);
   U4832 : XOR2_X1 port map( A => n7546, B => n4347, Z => 
                           DP_OP_719J1_125_1055xn38);
   U4833 : NAND2_X1 port map( A1 => n5692, A2 => fromMemoryPortxLOADEDDATAx(29)
                           , ZN => n4348);
   U4834 : NAND2_X1 port map( A1 => n4611, A2 => n4348, ZN => add_x_26xBx29x);
   U4835 : INV_X1 port map( A => add_x_26xBx29x, ZN => intadd_3xBx1x);
   U4836 : CLKBUF_X1 port map( A => n4349, Z => n5252);
   U4837 : CLKBUF_X1 port map( A => n5676, Z => n5677);
   U4838 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx29x,
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_24xx29x, ZN
                           => n4353);
   U4839 : AOI22_X1 port map( A1 => n5053, A2 => fromRegsPortxREG_FILE_29xx29x,
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx29x, ZN
                           => n4352);
   U4840 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_27xx29x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx29x, ZN
                           => n4351);
   U4841 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx29x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx29x, ZN
                           => n4350);
   U4842 : NAND4_X1 port map( A1 => n4353, A2 => n4352, A3 => n4351, A4 => 
                           n4350, ZN => n4359);
   U4843 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx29x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx29x, ZN
                           => n4357);
   U4844 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx29x,
                           B1 => n5288, B2 => fromRegsPortxREG_FILE_21xx29x, ZN
                           => n4356);
   U4845 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx29x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx29x, ZN
                           => n4355);
   U4846 : NAND2_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_19xx29x,
                           ZN => n4354);
   U4847 : NAND4_X1 port map( A1 => n4357, A2 => n4356, A3 => n4355, A4 => 
                           n4354, ZN => n4358);
   U4848 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4359
                           , A => n4358, ZN => n4365);
   U4849 : AOI22_X1 port map( A1 => n5301, A2 => fromRegsPortxREG_FILE_12xx29x,
                           B1 => n5302, B2 => fromRegsPortxREG_FILE_14xx29x, ZN
                           => n4364);
   U4850 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_11xx29x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx29x, ZN
                           => n4361);
   U4851 : CLKBUF_X1 port map( A => n5194, Z => n5304);
   U4852 : AOI22_X1 port map( A1 => n5309, A2 => fromRegsPortxREG_FILE_16xx29x,
                           B1 => n5304, B2 => fromRegsPortxREG_FILE_13xx29x, ZN
                           => n4360);
   U4853 : NAND2_X1 port map( A1 => n4361, A2 => n4360, ZN => n4362);
   U4854 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx29x, B2 => n5300,
                           A => n4362, ZN => n4363);
   U4855 : OAI211_X1 port map( C1 => n4365, C2 => n5758, A => n4364, B => n4363
                           , ZN => n4366);
   U4856 : NAND2_X1 port map( A1 => n4366, A2 => n5238, ZN => n4376);
   U4857 : AOI22_X1 port map( A1 => n5142, A2 => fromRegsPortxREG_FILE_03xx29x,
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx29x, ZN
                           => n4370);
   U4858 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx29x,
                           B1 => n5316, B2 => fromRegsPortxREG_FILE_06xx29x, ZN
                           => n4369);
   U4859 : AOI22_X1 port map( A1 => n5203, A2 => fromRegsPortxREG_FILE_09xx29x,
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx29x, ZN
                           => n4368);
   U4860 : NAND2_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_07xx29x,
                           ZN => n4367);
   U4861 : NAND4_X1 port map( A1 => n4370, A2 => n4369, A3 => n4368, A4 => 
                           n4367, ZN => n4374);
   U4862 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx29x,
                           ZN => n4372);
   U4863 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx29x, A2 => n5244,
                           ZN => n4371);
   U4864 : NAND2_X1 port map( A1 => n4372, A2 => n4371, ZN => n4373);
   U4865 : AOI21_X1 port map( B1 => n4374, B2 => n5331, A => n4373, ZN => n4375
                           );
   U4866 : NAND2_X1 port map( A1 => n4376, A2 => n4375, ZN => n7247);
   U4867 : INV_X1 port map( A => n7247, ZN => n7481);
   U4868 : OAI22_X1 port map( A1 => n5678, A2 => intadd_3xBx1x, B1 => n5677, B2
                           => n7481, ZN => n4377);
   U4869 : XOR2_X1 port map( A => n5252, B => n4377, Z => 
                           DP_OP_719J1_125_1055xn39);
   U4870 : NAND2_X1 port map( A1 => n5692, A2 => fromMemoryPortxLOADEDDATAx(28)
                           , ZN => n4378);
   U4871 : NAND2_X1 port map( A1 => n4611, A2 => n4378, ZN => add_x_26xBx28x);
   U4872 : INV_X1 port map( A => add_x_26xBx28x, ZN => intadd_3xBx0x);
   U4873 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx28x,
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx28x, ZN
                           => n4382);
   U4874 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_24xx28x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx28x, ZN
                           => n4381);
   U4875 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx28x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_27xx28x, ZN
                           => n4380);
   U4876 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx28x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx28x, ZN
                           => n4379);
   U4877 : NAND4_X1 port map( A1 => n4382, A2 => n4381, A3 => n4380, A4 => 
                           n4379, ZN => n4388);
   U4878 : AOI22_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx28x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx28x, ZN
                           => n4386);
   U4879 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx28x,
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_19xx28x, ZN
                           => n4385);
   U4880 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx28x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx28x, ZN
                           => n4384);
   U4881 : NAND2_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx28x,
                           ZN => n4383);
   U4882 : NAND4_X1 port map( A1 => n4386, A2 => n4385, A3 => n4384, A4 => 
                           n4383, ZN => n4387);
   U4883 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4388
                           , A => n4387, ZN => n4394);
   U4884 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_13xx28x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx28x, ZN
                           => n4393);
   U4885 : CLKBUF_X1 port map( A => n5301, Z => n5234);
   U4886 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx28x,
                           B1 => n5303, B2 => fromRegsPortxREG_FILE_11xx28x, ZN
                           => n4390);
   U4887 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx28x,
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx28x, ZN
                           => n4389);
   U4888 : NAND2_X1 port map( A1 => n4390, A2 => n4389, ZN => n4391);
   U4889 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx28x, B2 => n5234,
                           A => n4391, ZN => n4392);
   U4890 : OAI211_X1 port map( C1 => n4394, C2 => n5758, A => n4393, B => n4392
                           , ZN => n4395);
   U4891 : NAND2_X1 port map( A1 => n4395, A2 => n5238, ZN => n4405);
   U4892 : CLKBUF_X1 port map( A => n5142, Z => n5315);
   U4893 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx28x,
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx28x, ZN
                           => n4399);
   U4894 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx28x,
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx28x, ZN
                           => n4398);
   U4895 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx28x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx28x, ZN
                           => n4397);
   U4896 : NAND2_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx28x,
                           ZN => n4396);
   U4897 : NAND4_X1 port map( A1 => n4399, A2 => n4398, A3 => n4397, A4 => 
                           n4396, ZN => n4403);
   U4898 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx28x,
                           ZN => n4401);
   U4899 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx28x, A2 => n5244,
                           ZN => n4400);
   U4900 : NAND2_X1 port map( A1 => n4401, A2 => n4400, ZN => n4402);
   U4901 : AOI21_X1 port map( B1 => n4403, B2 => n5331, A => n4402, ZN => n4404
                           );
   U4902 : NAND2_X1 port map( A1 => n4405, A2 => n4404, ZN => n7237);
   U4903 : INV_X1 port map( A => n7237, ZN => n7480);
   U4904 : OAI22_X1 port map( A1 => n5678, A2 => intadd_3xBx0x, B1 => n5677, B2
                           => n7480, ZN => n4406);
   U4905 : XOR2_X1 port map( A => n7546, B => n4406, Z => 
                           DP_OP_719J1_125_1055xn40);
   U4906 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx27x,
                           B1 => n5278, B2 => fromRegsPortxREG_FILE_29xx27x, ZN
                           => n4410);
   U4907 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx27x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx27x, ZN
                           => n4409);
   U4908 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_26xx27x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_27xx27x, ZN
                           => n4408);
   U4909 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_24xx27x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx27x, ZN
                           => n4407);
   U4910 : NAND4_X1 port map( A1 => n4410, A2 => n4409, A3 => n4408, A4 => 
                           n4407, ZN => n4416);
   U4911 : AOI22_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_18xx27x,
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_19xx27x, ZN
                           => n4414);
   U4912 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx27x,
                           B1 => n5287, B2 => fromRegsPortxREG_FILE_22xx27x, ZN
                           => n4413);
   U4913 : AOI22_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx27x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx27x, ZN
                           => n4412);
   U4914 : NAND2_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx27x,
                           ZN => n4411);
   U4915 : NAND4_X1 port map( A1 => n4414, A2 => n4413, A3 => n4412, A4 => 
                           n4411, ZN => n4415);
   U4916 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4416
                           , A => n4415, ZN => n4422);
   U4917 : AOI22_X1 port map( A1 => n5102, A2 => fromRegsPortxREG_FILE_14xx27x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx27x, ZN
                           => n4421);
   U4918 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx27x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx27x, ZN
                           => n4418);
   U4919 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_11xx27x,
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx27x, ZN
                           => n4417);
   U4920 : NAND2_X1 port map( A1 => n4418, A2 => n4417, ZN => n4419);
   U4921 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx27x, B2 => n5301,
                           A => n4419, ZN => n4420);
   U4922 : OAI211_X1 port map( C1 => n4422, C2 => n5758, A => n4421, B => n4420
                           , ZN => n4423);
   U4923 : NAND2_X1 port map( A1 => n4423, A2 => n5238, ZN => n4433);
   U4924 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx27x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx27x, ZN
                           => n4427);
   U4925 : AOI22_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx27x,
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx27x, ZN
                           => n4426);
   U4926 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx27x,
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx27x, ZN
                           => n4425);
   U4927 : NAND2_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx27x,
                           ZN => n4424);
   U4928 : NAND4_X1 port map( A1 => n4427, A2 => n4426, A3 => n4425, A4 => 
                           n4424, ZN => n4431);
   U4929 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx27x,
                           ZN => n4429);
   U4930 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx27x, A2 => n5244,
                           ZN => n4428);
   U4931 : NAND2_X1 port map( A1 => n4429, A2 => n4428, ZN => n4430);
   U4932 : AOI21_X1 port map( B1 => n4431, B2 => n5331, A => n4430, ZN => n4432
                           );
   U4933 : NAND2_X1 port map( A1 => n4433, A2 => n4432, ZN => n7179);
   U4934 : INV_X1 port map( A => n7179, ZN => n7479);
   U4935 : CLKBUF_X1 port map( A => n5676, Z => n7360);
   U4936 : CLKBUF_X1 port map( A => n5673, Z => n5675);
   U4937 : INV_X1 port map( A => add_x_26xBx27x, ZN => n5462);
   U4938 : OAI22_X1 port map( A1 => n7479, A2 => n7360, B1 => n5675, B2 => 
                           n5462, ZN => n4434);
   U4939 : XOR2_X1 port map( A => n7546, B => n4434, Z => 
                           DP_OP_719J1_125_1055xn41);
   U4940 : NAND2_X1 port map( A1 => n5692, A2 => fromMemoryPortxLOADEDDATAx(26)
                           , ZN => n4435);
   U4941 : NAND2_X1 port map( A1 => n4611, A2 => n4435, ZN => add_x_26xBx26x);
   U4942 : INV_X1 port map( A => add_x_26xBx26x, ZN => n7120);
   U4943 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx26x,
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx26x, ZN
                           => n4439);
   U4944 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx26x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx26x, ZN
                           => n4438);
   U4945 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_24xx26x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_27xx26x, ZN
                           => n4437);
   U4946 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx26x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx26x, ZN
                           => n4436);
   U4947 : NAND4_X1 port map( A1 => n4439, A2 => n4438, A3 => n4437, A4 => 
                           n4436, ZN => n4445);
   U4948 : AOI22_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx26x,
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_19xx26x, ZN
                           => n4443);
   U4949 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx26x,
                           B1 => n5289, B2 => fromRegsPortxREG_FILE_23xx26x, ZN
                           => n4442);
   U4950 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx26x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx26x, ZN
                           => n4441);
   U4951 : NAND2_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_17xx26x,
                           ZN => n4440);
   U4952 : NAND4_X1 port map( A1 => n4443, A2 => n4442, A3 => n4441, A4 => 
                           n4440, ZN => n4444);
   U4953 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4445
                           , A => n4444, ZN => n4451);
   U4954 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_11xx26x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx26x, ZN
                           => n4450);
   U4955 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx26x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx26x, ZN
                           => n4447);
   U4956 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx26x,
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx26x, ZN
                           => n4446);
   U4957 : NAND2_X1 port map( A1 => n4447, A2 => n4446, ZN => n4448);
   U4958 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx26x, B2 => n5301,
                           A => n4448, ZN => n4449);
   U4959 : OAI211_X1 port map( C1 => n4451, C2 => n5758, A => n4450, B => n4449
                           , ZN => n4452);
   U4960 : NAND2_X1 port map( A1 => n4452, A2 => n5238, ZN => n4462);
   U4961 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx26x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx26x, ZN
                           => n4456);
   U4962 : AOI22_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx26x,
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx26x, ZN
                           => n4455);
   U4963 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx26x,
                           B1 => n5315, B2 => fromRegsPortxREG_FILE_03xx26x, ZN
                           => n4454);
   U4964 : NAND2_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_05xx26x,
                           ZN => n4453);
   U4965 : NAND4_X1 port map( A1 => n4456, A2 => n4455, A3 => n4454, A4 => 
                           n4453, ZN => n4460);
   U4966 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx26x,
                           ZN => n4458);
   U4967 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx26x, A2 => n5244,
                           ZN => n4457);
   U4968 : NAND2_X1 port map( A1 => n4458, A2 => n4457, ZN => n4459);
   U4969 : AOI21_X1 port map( B1 => n4460, B2 => n5331, A => n4459, ZN => n4461
                           );
   U4970 : NAND2_X1 port map( A1 => n4462, A2 => n4461, ZN => n7114);
   U4971 : INV_X1 port map( A => n7114, ZN => n7478);
   U4972 : OAI22_X1 port map( A1 => n5678, A2 => n7120, B1 => n7360, B2 => 
                           n7478, ZN => n4463);
   U4973 : XOR2_X1 port map( A => n5252, B => n4463, Z => 
                           DP_OP_719J1_125_1055xn42);
   U4974 : NAND2_X1 port map( A1 => n5692, A2 => fromMemoryPortxLOADEDDATAx(25)
                           , ZN => n4464);
   U4975 : NAND2_X1 port map( A1 => n4611, A2 => n4464, ZN => add_x_26xBx25x);
   U4976 : INV_X1 port map( A => add_x_26xBx25x, ZN => n7076);
   U4977 : AOI22_X1 port map( A1 => n5053, A2 => fromRegsPortxREG_FILE_29xx25x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx25x, ZN
                           => n4468);
   U4978 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx25x,
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_24xx25x, ZN
                           => n4467);
   U4979 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx25x,
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx25x, ZN
                           => n4466);
   U4980 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_27xx25x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx25x, ZN
                           => n4465);
   U4981 : NAND4_X1 port map( A1 => n4468, A2 => n4467, A3 => n4466, A4 => 
                           n4465, ZN => n4474);
   U4982 : AOI22_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx25x,
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_19xx25x, ZN
                           => n4472);
   U4983 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx25x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx25x, ZN
                           => n4471);
   U4984 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx25x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx25x, ZN
                           => n4470);
   U4985 : NAND2_X1 port map( A1 => n5287, A2 => fromRegsPortxREG_FILE_22xx25x,
                           ZN => n4469);
   U4986 : NAND4_X1 port map( A1 => n4472, A2 => n4471, A3 => n4470, A4 => 
                           n4469, ZN => n4473);
   U4987 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4474
                           , A => n4473, ZN => n4480);
   U4988 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx25x,
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx25x, ZN
                           => n4479);
   U4989 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx25x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx25x, ZN
                           => n4476);
   U4990 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_11xx25x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx25x, ZN
                           => n4475);
   U4991 : NAND2_X1 port map( A1 => n4476, A2 => n4475, ZN => n4477);
   U4992 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx25x, B2 => n5301,
                           A => n4477, ZN => n4478);
   U4993 : OAI211_X1 port map( C1 => n4480, C2 => n5758, A => n4479, B => n4478
                           , ZN => n4481);
   U4994 : NAND2_X1 port map( A1 => n4481, A2 => n5238, ZN => n4491);
   U4995 : AOI22_X1 port map( A1 => n5142, A2 => fromRegsPortxREG_FILE_03xx25x,
                           B1 => n5316, B2 => fromRegsPortxREG_FILE_06xx25x, ZN
                           => n4485);
   U4996 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx25x,
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx25x, ZN
                           => n4484);
   U4997 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_05xx25x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx25x, ZN
                           => n4483);
   U4998 : NAND2_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx25x,
                           ZN => n4482);
   U4999 : NAND4_X1 port map( A1 => n4485, A2 => n4484, A3 => n4483, A4 => 
                           n4482, ZN => n4489);
   U5000 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx25x,
                           ZN => n4487);
   U5001 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx25x, A2 => n5244,
                           ZN => n4486);
   U5002 : NAND2_X1 port map( A1 => n4487, A2 => n4486, ZN => n4488);
   U5003 : AOI21_X1 port map( B1 => n4489, B2 => n5331, A => n4488, ZN => n4490
                           );
   U5004 : NAND2_X1 port map( A1 => n4491, A2 => n4490, ZN => n7093);
   U5005 : INV_X1 port map( A => n7093, ZN => n7477);
   U5006 : OAI22_X1 port map( A1 => n5678, A2 => n7076, B1 => n5674, B2 => 
                           n7477, ZN => n4492);
   U5007 : XOR2_X1 port map( A => n7546, B => n4492, Z => 
                           DP_OP_719J1_125_1055xn43);
   U5008 : NAND2_X1 port map( A1 => n5692, A2 => fromMemoryPortxLOADEDDATAx(24)
                           , ZN => n4493);
   U5009 : NAND2_X1 port map( A1 => n4611, A2 => n4493, ZN => add_x_26xBx24x);
   U5010 : INV_X1 port map( A => add_x_26xBx24x, ZN => intadd_1xBx7x);
   U5011 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_26xx24x,
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_24xx24x, ZN
                           => n4497);
   U5012 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx24x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx24x, ZN
                           => n4496);
   U5013 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx24x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_27xx24x, ZN
                           => n4495);
   U5014 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx24x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx24x, ZN
                           => n4494);
   U5015 : NAND4_X1 port map( A1 => n4497, A2 => n4496, A3 => n4495, A4 => 
                           n4494, ZN => n4503);
   U5016 : AOI22_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx24x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx24x, ZN
                           => n4501);
   U5017 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx24x,
                           B1 => n5289, B2 => fromRegsPortxREG_FILE_23xx24x, ZN
                           => n4500);
   U5018 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx24x,
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_19xx24x, ZN
                           => n4499);
   U5019 : NAND2_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_18xx24x,
                           ZN => n4498);
   U5020 : NAND4_X1 port map( A1 => n4501, A2 => n4500, A3 => n4499, A4 => 
                           n4498, ZN => n4502);
   U5021 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4503
                           , A => n4502, ZN => n4509);
   U5022 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx24x,
                           B1 => n5301, B2 => fromRegsPortxREG_FILE_12xx24x, ZN
                           => n4508);
   U5023 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx24x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx24x, ZN
                           => n4505);
   U5024 : AOI22_X1 port map( A1 => n5309, A2 => fromRegsPortxREG_FILE_16xx24x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx24x, ZN
                           => n4504);
   U5025 : NAND2_X1 port map( A1 => n4505, A2 => n4504, ZN => n4506);
   U5026 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_11xx24x, B2 => n5303,
                           A => n4506, ZN => n4507);
   U5027 : OAI211_X1 port map( C1 => n4509, C2 => n5758, A => n4508, B => n4507
                           , ZN => n4510);
   U5028 : NAND2_X1 port map( A1 => n4510, A2 => n5238, ZN => n4520);
   U5029 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_08xx24x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx24x, ZN
                           => n4514);
   U5030 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx24x,
                           B1 => n5316, B2 => fromRegsPortxREG_FILE_06xx24x, ZN
                           => n4513);
   U5031 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx24x,
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx24x, ZN
                           => n4512);
   U5032 : NAND2_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx24x,
                           ZN => n4511);
   U5033 : NAND4_X1 port map( A1 => n4514, A2 => n4513, A3 => n4512, A4 => 
                           n4511, ZN => n4518);
   U5034 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx24x,
                           ZN => n4516);
   U5035 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx24x, A2 => n5244,
                           ZN => n4515);
   U5036 : NAND2_X1 port map( A1 => n4516, A2 => n4515, ZN => n4517);
   U5037 : AOI21_X1 port map( B1 => n4518, B2 => n5331, A => n4517, ZN => n4519
                           );
   U5038 : NAND2_X1 port map( A1 => n4520, A2 => n4519, ZN => n5744);
   U5039 : INV_X1 port map( A => n5744, ZN => n7476);
   U5040 : OAI22_X1 port map( A1 => n5673, A2 => intadd_1xBx7x, B1 => n5674, B2
                           => n7476, ZN => n4521);
   U5041 : XOR2_X1 port map( A => n7546, B => n4521, Z => 
                           DP_OP_719J1_125_1055xn44);
   U5042 : NAND2_X1 port map( A1 => n4611, A2 => n7065, ZN => n4522);
   U5043 : AND2_X1 port map( A1 => n4552, A2 => n4522, ZN => add_x_26xBx23x);
   U5044 : INV_X1 port map( A => add_x_26xBx23x, ZN => intadd_1xBx6x);
   U5045 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx23x,
                           B1 => n5278, B2 => fromRegsPortxREG_FILE_29xx23x, ZN
                           => n4526);
   U5046 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_24xx23x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_27xx23x, ZN
                           => n4525);
   U5047 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx23x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx23x, ZN
                           => n4524);
   U5048 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_26xx23x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx23x, ZN
                           => n4523);
   U5049 : NAND4_X1 port map( A1 => n4526, A2 => n4525, A3 => n4524, A4 => 
                           n4523, ZN => n4532);
   U5050 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx23x,
                           B1 => n5126, B2 => fromRegsPortxREG_FILE_23xx23x, ZN
                           => n4530);
   U5051 : AOI22_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx23x,
                           B1 => n5224, B2 => fromRegsPortxREG_FILE_22xx23x, ZN
                           => n4529);
   U5052 : AOI22_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_18xx23x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx23x, ZN
                           => n4528);
   U5053 : NAND2_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_19xx23x,
                           ZN => n4527);
   U5054 : NAND4_X1 port map( A1 => n4530, A2 => n4529, A3 => n4528, A4 => 
                           n4527, ZN => n4531);
   U5055 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4532
                           , A => n4531, ZN => n4538);
   U5056 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx23x,
                           B1 => n5065, B2 => fromRegsPortxREG_FILE_16xx23x, ZN
                           => n4537);
   U5057 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx23x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx23x, ZN
                           => n4534);
   U5058 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_11xx23x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx23x, ZN
                           => n4533);
   U5059 : NAND2_X1 port map( A1 => n4534, A2 => n4533, ZN => n4535);
   U5060 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx23x, B2 => n5234,
                           A => n4535, ZN => n4536);
   U5061 : OAI211_X1 port map( C1 => n4538, C2 => n5200, A => n4537, B => n4536
                           , ZN => n4539);
   U5062 : NAND2_X1 port map( A1 => n4539, A2 => n5238, ZN => n4549);
   U5063 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx23x,
                           B1 => n5316, B2 => fromRegsPortxREG_FILE_06xx23x, ZN
                           => n4543);
   U5064 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx23x,
                           B1 => n5010, B2 => fromRegsPortxREG_FILE_05xx23x, ZN
                           => n4542);
   U5065 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx23x,
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx23x, ZN
                           => n4541);
   U5066 : NAND2_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_07xx23x,
                           ZN => n4540);
   U5067 : NAND4_X1 port map( A1 => n4543, A2 => n4542, A3 => n4541, A4 => 
                           n4540, ZN => n4547);
   U5068 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx23x,
                           ZN => n4545);
   U5069 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx23x, A2 => n5244,
                           ZN => n4544);
   U5070 : NAND2_X1 port map( A1 => n4545, A2 => n4544, ZN => n4546);
   U5071 : AOI21_X1 port map( B1 => n4547, B2 => n5331, A => n4546, ZN => n4548
                           );
   U5072 : NAND2_X1 port map( A1 => n4549, A2 => n4548, ZN => n7028);
   U5073 : INV_X1 port map( A => n7028, ZN => n7475);
   U5074 : OAI22_X1 port map( A1 => n7475, A2 => n5674, B1 => n5675, B2 => 
                           intadd_1xBx6x, ZN => n4550);
   U5075 : XOR2_X1 port map( A => n5252, B => n4550, Z => 
                           DP_OP_719J1_125_1055xn45);
   U5076 : NAND2_X1 port map( A1 => n4611, A2 => n7027, ZN => n4551);
   U5077 : AND2_X1 port map( A1 => n4552, A2 => n4551, ZN => add_x_26xBx22x);
   U5078 : INV_X1 port map( A => add_x_26xBx22x, ZN => intadd_1xBx5x);
   U5079 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_26xx22x,
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_24xx22x, ZN
                           => n4556);
   U5080 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx22x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_27xx22x, ZN
                           => n4555);
   U5081 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx22x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx22x, ZN
                           => n4554);
   U5082 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx22x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx22x, ZN
                           => n4553);
   U5083 : NAND4_X1 port map( A1 => n4556, A2 => n4555, A3 => n4554, A4 => 
                           n4553, ZN => n4562);
   U5084 : AOI22_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_18xx22x,
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_19xx22x, ZN
                           => n4560);
   U5085 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx22x,
                           B1 => n5288, B2 => fromRegsPortxREG_FILE_21xx22x, ZN
                           => n4559);
   U5086 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx22x,
                           B1 => n5224, B2 => fromRegsPortxREG_FILE_22xx22x, ZN
                           => n4558);
   U5087 : NAND2_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_17xx22x,
                           ZN => n4557);
   U5088 : NAND4_X1 port map( A1 => n4560, A2 => n4559, A3 => n4558, A4 => 
                           n4557, ZN => n4561);
   U5089 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4562
                           , A => n4561, ZN => n4568);
   U5090 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx22x,
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx22x, ZN
                           => n4567);
   U5091 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx22x,
                           B1 => n5303, B2 => fromRegsPortxREG_FILE_11xx22x, ZN
                           => n4564);
   U5092 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_13xx22x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx22x, ZN
                           => n4563);
   U5093 : NAND2_X1 port map( A1 => n4564, A2 => n4563, ZN => n4565);
   U5094 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx22x, B2 => n5234,
                           A => n4565, ZN => n4566);
   U5095 : OAI211_X1 port map( C1 => n4568, C2 => n5200, A => n4567, B => n4566
                           , ZN => n4569);
   U5096 : NAND2_X1 port map( A1 => n4569, A2 => n5238, ZN => n4579);
   U5097 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx22x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx22x, ZN
                           => n4573);
   U5098 : AOI22_X1 port map( A1 => n5039, A2 => fromRegsPortxREG_FILE_08xx22x,
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx22x, ZN
                           => n4572);
   U5099 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx22x,
                           B1 => n5315, B2 => fromRegsPortxREG_FILE_03xx22x, ZN
                           => n4571);
   U5100 : NAND2_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx22x,
                           ZN => n4570);
   U5101 : NAND4_X1 port map( A1 => n4573, A2 => n4572, A3 => n4571, A4 => 
                           n4570, ZN => n4577);
   U5102 : NAND2_X1 port map( A1 => n4867, A2 => fromRegsPortxREG_FILE_02xx22x,
                           ZN => n4575);
   U5103 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx22x, A2 => n5244,
                           ZN => n4574);
   U5104 : NAND2_X1 port map( A1 => n4575, A2 => n4574, ZN => n4576);
   U5105 : AOI21_X1 port map( B1 => n4577, B2 => n5331, A => n4576, ZN => n4578
                           );
   U5106 : NAND2_X1 port map( A1 => n4579, A2 => n4578, ZN => n6986);
   U5107 : INV_X1 port map( A => n6986, ZN => n7474);
   U5108 : OAI22_X1 port map( A1 => n5673, A2 => intadd_1xBx5x, B1 => n5677, B2
                           => n7474, ZN => n4580);
   U5109 : XOR2_X1 port map( A => n5252, B => n4580, Z => 
                           DP_OP_719J1_125_1055xn46);
   U5110 : NAND2_X1 port map( A1 => n5692, A2 => fromMemoryPortxLOADEDDATAx(21)
                           , ZN => n4581);
   U5111 : NAND2_X1 port map( A1 => n4611, A2 => n4581, ZN => add_x_26xBx21x);
   U5112 : INV_X1 port map( A => add_x_26xBx21x, ZN => intadd_1xBx4x);
   U5113 : AOI22_X1 port map( A1 => n5120, A2 => fromRegsPortxREG_FILE_24xx21x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx21x, ZN
                           => n4585);
   U5114 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx21x,
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx21x, ZN
                           => n4584);
   U5115 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx21x,
                           B1 => n5278, B2 => fromRegsPortxREG_FILE_29xx21x, ZN
                           => n4583);
   U5116 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_27xx21x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx21x, ZN
                           => n4582);
   U5117 : NAND4_X1 port map( A1 => n4585, A2 => n4584, A3 => n4583, A4 => 
                           n4582, ZN => n4591);
   U5118 : AOI22_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx21x,
                           B1 => n5224, B2 => fromRegsPortxREG_FILE_22xx21x, ZN
                           => n4589);
   U5119 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx21x,
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_19xx21x, ZN
                           => n4588);
   U5120 : AOI22_X1 port map( A1 => n5093, A2 => fromRegsPortxREG_FILE_18xx21x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx21x, ZN
                           => n4587);
   U5121 : NAND2_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx21x,
                           ZN => n4586);
   U5122 : NAND4_X1 port map( A1 => n4589, A2 => n4588, A3 => n4587, A4 => 
                           n4586, ZN => n4590);
   U5123 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4591
                           , A => n4590, ZN => n4597);
   U5124 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_11xx21x,
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx21x, ZN
                           => n4596);
   U5125 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx21x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx21x, ZN
                           => n4593);
   U5126 : AOI22_X1 port map( A1 => n5301, A2 => fromRegsPortxREG_FILE_12xx21x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx21x, ZN
                           => n4592);
   U5127 : NAND2_X1 port map( A1 => n4593, A2 => n4592, ZN => n4594);
   U5128 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx21x, B2 => n5300,
                           A => n4594, ZN => n4595);
   U5129 : OAI211_X1 port map( C1 => n4597, C2 => n5200, A => n4596, B => n4595
                           , ZN => n4598);
   U5130 : NAND2_X1 port map( A1 => n4598, A2 => n5238, ZN => n4608);
   U5131 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx21x,
                           B1 => n5316, B2 => fromRegsPortxREG_FILE_06xx21x, ZN
                           => n4602);
   U5132 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx21x,
                           B1 => n5010, B2 => fromRegsPortxREG_FILE_05xx21x, ZN
                           => n4601);
   U5133 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx21x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx21x, ZN
                           => n4600);
   U5134 : NAND2_X1 port map( A1 => n5039, A2 => fromRegsPortxREG_FILE_08xx21x,
                           ZN => n4599);
   U5135 : NAND4_X1 port map( A1 => n4602, A2 => n4601, A3 => n4600, A4 => 
                           n4599, ZN => n4606);
   U5136 : NAND2_X1 port map( A1 => n4867, A2 => fromRegsPortxREG_FILE_02xx21x,
                           ZN => n4604);
   U5137 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx21x, A2 => n5244,
                           ZN => n4603);
   U5138 : NAND2_X1 port map( A1 => n4604, A2 => n4603, ZN => n4605);
   U5139 : AOI21_X1 port map( B1 => n4606, B2 => n5331, A => n4605, ZN => n4607
                           );
   U5140 : NAND2_X1 port map( A1 => n4608, A2 => n4607, ZN => n5717);
   U5141 : INV_X1 port map( A => n5717, ZN => n7473);
   U5142 : OAI22_X1 port map( A1 => n5673, A2 => intadd_1xBx4x, B1 => n5676, B2
                           => n7473, ZN => n4609);
   U5143 : XOR2_X1 port map( A => n5252, B => n4609, Z => 
                           DP_OP_719J1_125_1055xn47);
   U5144 : NAND2_X1 port map( A1 => n5692, A2 => fromMemoryPortxLOADEDDATAx(20)
                           , ZN => n4610);
   U5145 : NAND2_X1 port map( A1 => n4611, A2 => n4610, ZN => add_x_26xBx20x);
   U5146 : INV_X1 port map( A => add_x_26xBx20x, ZN => intadd_1xBx3x);
   U5147 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx20x,
                           B1 => n5120, B2 => fromRegsPortxREG_FILE_24xx20x, ZN
                           => n4615);
   U5148 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx20x,
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx20x, ZN
                           => n4614);
   U5149 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx20x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_27xx20x, ZN
                           => n4613);
   U5150 : AOI22_X1 port map( A1 => n5282, A2 => fromRegsPortxREG_FILE_31xx20x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx20x, ZN
                           => n4612);
   U5151 : NAND4_X1 port map( A1 => n4615, A2 => n4614, A3 => n4613, A4 => 
                           n4612, ZN => n4621);
   U5152 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx20x,
                           B1 => n5224, B2 => fromRegsPortxREG_FILE_22xx20x, ZN
                           => n4619);
   U5153 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx20x,
                           B1 => n5093, B2 => fromRegsPortxREG_FILE_18xx20x, ZN
                           => n4618);
   U5154 : AOI22_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx20x,
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_19xx20x, ZN
                           => n4617);
   U5155 : NAND2_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_17xx20x,
                           ZN => n4616);
   U5156 : NAND4_X1 port map( A1 => n4619, A2 => n4618, A3 => n4617, A4 => 
                           n4616, ZN => n4620);
   U5157 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4621
                           , A => n4620, ZN => n4627);
   U5158 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx20x,
                           B1 => n5065, B2 => fromRegsPortxREG_FILE_16xx20x, ZN
                           => n4626);
   U5159 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx20x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx20x, ZN
                           => n4623);
   U5160 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_11xx20x,
                           B1 => n5304, B2 => fromRegsPortxREG_FILE_13xx20x, ZN
                           => n4622);
   U5161 : NAND2_X1 port map( A1 => n4623, A2 => n4622, ZN => n4624);
   U5162 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx20x, B2 => n5234,
                           A => n4624, ZN => n4625);
   U5163 : OAI211_X1 port map( C1 => n4627, C2 => n5200, A => n4626, B => n4625
                           , ZN => n4628);
   U5164 : NAND2_X1 port map( A1 => n4628, A2 => n5238, ZN => n4638);
   U5165 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx20x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx20x, ZN
                           => n4632);
   U5166 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx20x,
                           B1 => n5010, B2 => fromRegsPortxREG_FILE_05xx20x, ZN
                           => n4631);
   U5167 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx20x,
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx20x, ZN
                           => n4630);
   U5168 : NAND2_X1 port map( A1 => n5141, A2 => fromRegsPortxREG_FILE_06xx20x,
                           ZN => n4629);
   U5169 : NAND4_X1 port map( A1 => n4632, A2 => n4631, A3 => n4630, A4 => 
                           n4629, ZN => n4636);
   U5170 : NAND2_X1 port map( A1 => n4867, A2 => fromRegsPortxREG_FILE_02xx20x,
                           ZN => n4634);
   U5171 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx20x, A2 => n5244,
                           ZN => n4633);
   U5172 : NAND2_X1 port map( A1 => n4634, A2 => n4633, ZN => n4635);
   U5173 : AOI21_X1 port map( B1 => n4636, B2 => n5331, A => n4635, ZN => n4637
                           );
   U5174 : NAND2_X1 port map( A1 => n4638, A2 => n4637, ZN => n6962);
   U5175 : INV_X1 port map( A => n6962, ZN => n7472);
   U5176 : OAI22_X1 port map( A1 => n5673, A2 => intadd_1xBx3x, B1 => n5674, B2
                           => n7472, ZN => n4639);
   U5177 : XOR2_X1 port map( A => n5252, B => n4639, Z => 
                           DP_OP_719J1_125_1055xn48);
   U5178 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(31), A2 => n4640,
                           ZN => n4876);
   U5179 : AOI21_X1 port map( B1 => n4875, B2 => fromMemoryPortxLOADEDDATAx(31)
                           , A => n4876, ZN => n5652);
   U5180 : NAND2_X1 port map( A1 => n7441, A2 => fromMemoryPortxLOADEDDATAx(3),
                           ZN => n5641);
   U5181 : NAND2_X1 port map( A1 => n5641, A2 => n4641, ZN => n5650);
   U5182 : NAND2_X1 port map( A1 => n5650, A2 => fromMemoryPortxLOADEDDATAx(19)
                           , ZN => n4642);
   U5183 : NAND2_X1 port map( A1 => n5652, A2 => n4642, ZN => add_x_26xBx19x);
   U5184 : INV_X1 port map( A => add_x_26xBx19x, ZN => intadd_1xBx2x);
   U5185 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_26xx19x,
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_24xx19x, ZN
                           => n4646);
   U5186 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx19x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_27xx19x, ZN
                           => n4645);
   U5187 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx19x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx19x, ZN
                           => n4644);
   U5188 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx19x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx19x, ZN
                           => n4643);
   U5189 : NAND4_X1 port map( A1 => n4646, A2 => n4645, A3 => n4644, A4 => 
                           n4643, ZN => n4652);
   U5190 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx19x,
                           B1 => n5288, B2 => fromRegsPortxREG_FILE_21xx19x, ZN
                           => n4650);
   U5191 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx19x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx19x, ZN
                           => n4649);
   U5192 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx19x,
                           B1 => n5093, B2 => fromRegsPortxREG_FILE_18xx19x, ZN
                           => n4648);
   U5193 : NAND2_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_19xx19x,
                           ZN => n4647);
   U5194 : NAND4_X1 port map( A1 => n4650, A2 => n4649, A3 => n4648, A4 => 
                           n4647, ZN => n4651);
   U5195 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4652
                           , A => n4651, ZN => n4658);
   U5196 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_13xx19x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx19x, ZN
                           => n4657);
   U5197 : AOI22_X1 port map( A1 => n5102, A2 => fromRegsPortxREG_FILE_14xx19x,
                           B1 => n5303, B2 => fromRegsPortxREG_FILE_11xx19x, ZN
                           => n4654);
   U5198 : AOI22_X1 port map( A1 => n5301, A2 => fromRegsPortxREG_FILE_12xx19x,
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx19x, ZN
                           => n4653);
   U5199 : NAND2_X1 port map( A1 => n4654, A2 => n4653, ZN => n4655);
   U5200 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx19x, B2 => n5300,
                           A => n4655, ZN => n4656);
   U5201 : OAI211_X1 port map( C1 => n4658, C2 => n5200, A => n4657, B => n4656
                           , ZN => n4659);
   U5202 : NAND2_X1 port map( A1 => n4659, A2 => n5238, ZN => n4669);
   U5203 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx19x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx19x, ZN
                           => n4663);
   U5204 : AOI22_X1 port map( A1 => n5141, A2 => fromRegsPortxREG_FILE_06xx19x,
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx19x, ZN
                           => n4662);
   U5205 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx19x,
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx19x, ZN
                           => n4661);
   U5206 : NAND2_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx19x,
                           ZN => n4660);
   U5207 : NAND4_X1 port map( A1 => n4663, A2 => n4662, A3 => n4661, A4 => 
                           n4660, ZN => n4667);
   U5208 : NAND2_X1 port map( A1 => n4867, A2 => fromRegsPortxREG_FILE_02xx19x,
                           ZN => n4665);
   U5209 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx19x, A2 => n5244,
                           ZN => n4664);
   U5210 : NAND2_X1 port map( A1 => n4665, A2 => n4664, ZN => n4666);
   U5211 : AOI21_X1 port map( B1 => n4667, B2 => n5331, A => n4666, ZN => n4668
                           );
   U5212 : NAND2_X1 port map( A1 => n4669, A2 => n4668, ZN => n6918);
   U5213 : INV_X1 port map( A => n6918, ZN => n7471);
   U5214 : OAI22_X1 port map( A1 => n5673, A2 => intadd_1xBx2x, B1 => n5676, B2
                           => n7471, ZN => n4670);
   U5215 : XOR2_X1 port map( A => n7546, B => n4670, Z => 
                           DP_OP_719J1_125_1055xn49);
   U5216 : NAND2_X1 port map( A1 => n5650, A2 => fromMemoryPortxLOADEDDATAx(18)
                           , ZN => n4671);
   U5217 : NAND2_X1 port map( A1 => n5652, A2 => n4671, ZN => add_x_26xBx18x);
   U5218 : INV_X1 port map( A => add_x_26xBx18x, ZN => intadd_1xBx1x);
   U5219 : AOI22_X1 port map( A1 => n5120, A2 => fromRegsPortxREG_FILE_24xx18x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx18x, ZN
                           => n4675);
   U5220 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx18x,
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx18x, ZN
                           => n4674);
   U5221 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx18x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_27xx18x, ZN
                           => n4673);
   U5222 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx18x,
                           B1 => n5054, B2 => fromRegsPortxREG_FILE_31xx18x, ZN
                           => n4672);
   U5223 : NAND4_X1 port map( A1 => n4675, A2 => n4674, A3 => n4673, A4 => 
                           n4672, ZN => n4681);
   U5224 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx18x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx18x, ZN
                           => n4679);
   U5225 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx18x,
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_19xx18x, ZN
                           => n4678);
   U5226 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx18x,
                           B1 => n5093, B2 => fromRegsPortxREG_FILE_18xx18x, ZN
                           => n4677);
   U5227 : NAND2_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx18x,
                           ZN => n4676);
   U5228 : NAND4_X1 port map( A1 => n4679, A2 => n4678, A3 => n4677, A4 => 
                           n4676, ZN => n4680);
   U5229 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4681
                           , A => n4680, ZN => n4687);
   U5230 : AOI22_X1 port map( A1 => n5301, A2 => fromRegsPortxREG_FILE_12xx18x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx18x, ZN
                           => n4686);
   U5231 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx18x,
                           B1 => n5303, B2 => fromRegsPortxREG_FILE_11xx18x, ZN
                           => n4683);
   U5232 : AOI22_X1 port map( A1 => n5065, A2 => fromRegsPortxREG_FILE_16xx18x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx18x, ZN
                           => n4682);
   U5233 : NAND2_X1 port map( A1 => n4683, A2 => n4682, ZN => n4684);
   U5234 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx18x, B2 => n5165,
                           A => n4684, ZN => n4685);
   U5235 : OAI211_X1 port map( C1 => n4687, C2 => n5200, A => n4686, B => n4685
                           , ZN => n4688);
   U5236 : NAND2_X1 port map( A1 => n4688, A2 => n5238, ZN => n4698);
   U5237 : AOI22_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx18x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx18x, ZN
                           => n4692);
   U5238 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx18x,
                           B1 => n5039, B2 => fromRegsPortxREG_FILE_08xx18x, ZN
                           => n4691);
   U5239 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx18x,
                           B1 => n5315, B2 => fromRegsPortxREG_FILE_03xx18x, ZN
                           => n4690);
   U5240 : NAND2_X1 port map( A1 => n5010, A2 => fromRegsPortxREG_FILE_05xx18x,
                           ZN => n4689);
   U5241 : NAND4_X1 port map( A1 => n4692, A2 => n4691, A3 => n4690, A4 => 
                           n4689, ZN => n4696);
   U5242 : NAND2_X1 port map( A1 => n4867, A2 => fromRegsPortxREG_FILE_02xx18x,
                           ZN => n4694);
   U5243 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx18x, A2 => n5244,
                           ZN => n4693);
   U5244 : NAND2_X1 port map( A1 => n4694, A2 => n4693, ZN => n4695);
   U5245 : AOI21_X1 port map( B1 => n4696, B2 => n5331, A => n4695, ZN => n4697
                           );
   U5246 : NAND2_X1 port map( A1 => n4698, A2 => n4697, ZN => n6891);
   U5247 : INV_X1 port map( A => n6891, ZN => n7470);
   U5248 : OAI22_X1 port map( A1 => n7470, A2 => n5676, B1 => n5675, B2 => 
                           intadd_1xBx1x, ZN => n4699);
   U5249 : XOR2_X1 port map( A => n5252, B => n4699, Z => 
                           DP_OP_719J1_125_1055xn50);
   U5250 : NAND2_X1 port map( A1 => n5650, A2 => fromMemoryPortxLOADEDDATAx(17)
                           , ZN => n4700);
   U5251 : NAND2_X1 port map( A1 => n5652, A2 => n4700, ZN => add_x_26xBx17x);
   U5252 : INV_X1 port map( A => add_x_26xBx17x, ZN => intadd_1xBx0x);
   U5253 : AOI22_X1 port map( A1 => n5087, A2 => fromRegsPortxREG_FILE_26xx17x,
                           B1 => n5120, B2 => fromRegsPortxREG_FILE_24xx17x, ZN
                           => n4704);
   U5254 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx17x,
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_27xx17x, ZN
                           => n4703);
   U5255 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx17x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx17x, ZN
                           => n4702);
   U5256 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx17x,
                           B1 => n5054, B2 => fromRegsPortxREG_FILE_31xx17x, ZN
                           => n4701);
   U5257 : NAND4_X1 port map( A1 => n4704, A2 => n4703, A3 => n4702, A4 => 
                           n4701, ZN => n4710);
   U5258 : AOI22_X1 port map( A1 => n5093, A2 => fromRegsPortxREG_FILE_18xx17x,
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_19xx17x, ZN
                           => n4708);
   U5259 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx17x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx17x, ZN
                           => n4707);
   U5260 : AOI22_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx17x,
                           B1 => n5287, B2 => fromRegsPortxREG_FILE_22xx17x, ZN
                           => n4706);
   U5261 : NAND2_X1 port map( A1 => n5092, A2 => fromRegsPortxREG_FILE_20xx17x,
                           ZN => n4705);
   U5262 : NAND4_X1 port map( A1 => n4708, A2 => n4707, A3 => n4706, A4 => 
                           n4705, ZN => n4709);
   U5263 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4710
                           , A => n4709, ZN => n4716);
   U5264 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_13xx17x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx17x, ZN
                           => n4715);
   U5265 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx17x,
                           B1 => n5303, B2 => fromRegsPortxREG_FILE_11xx17x, ZN
                           => n4712);
   U5266 : AOI22_X1 port map( A1 => n5301, A2 => fromRegsPortxREG_FILE_12xx17x,
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx17x, ZN
                           => n4711);
   U5267 : NAND2_X1 port map( A1 => n4712, A2 => n4711, ZN => n4713);
   U5268 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx17x, B2 => n5165,
                           A => n4713, ZN => n4714);
   U5269 : OAI211_X1 port map( C1 => n4716, C2 => n5200, A => n4715, B => n4714
                           , ZN => n4717);
   U5270 : NAND2_X1 port map( A1 => n4717, A2 => n5238, ZN => n4727);
   U5271 : AOI22_X1 port map( A1 => n5039, A2 => fromRegsPortxREG_FILE_08xx17x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx17x, ZN
                           => n4721);
   U5272 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx17x,
                           B1 => n5141, B2 => fromRegsPortxREG_FILE_06xx17x, ZN
                           => n4720);
   U5273 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx17x,
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx17x, ZN
                           => n4719);
   U5274 : NAND2_X1 port map( A1 => n5073, A2 => fromRegsPortxREG_FILE_04xx17x,
                           ZN => n4718);
   U5275 : NAND4_X1 port map( A1 => n4721, A2 => n4720, A3 => n4719, A4 => 
                           n4718, ZN => n4725);
   U5276 : NAND2_X1 port map( A1 => n4867, A2 => fromRegsPortxREG_FILE_02xx17x,
                           ZN => n4723);
   U5277 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx17x, A2 => n5244,
                           ZN => n4722);
   U5278 : NAND2_X1 port map( A1 => n4723, A2 => n4722, ZN => n4724);
   U5279 : AOI21_X1 port map( B1 => n4725, B2 => n5331, A => n4724, ZN => n4726
                           );
   U5280 : NAND2_X1 port map( A1 => n4727, A2 => n4726, ZN => n6835);
   U5281 : INV_X1 port map( A => n6835, ZN => n7469);
   U5282 : OAI22_X1 port map( A1 => n5678, A2 => intadd_1xBx0x, B1 => n5674, B2
                           => n7469, ZN => n4728);
   U5283 : XOR2_X1 port map( A => n5252, B => n4728, Z => 
                           DP_OP_719J1_125_1055xn51);
   U5284 : NAND2_X1 port map( A1 => n5650, A2 => fromMemoryPortxLOADEDDATAx(16)
                           , ZN => n4729);
   U5285 : NAND2_X1 port map( A1 => n5652, A2 => n4729, ZN => add_x_26xBx16x);
   U5286 : INV_X1 port map( A => add_x_26xBx16x, ZN => n6811);
   U5287 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx16x,
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_27xx16x, ZN
                           => n4733);
   U5288 : AOI22_X1 port map( A1 => n5087, A2 => fromRegsPortxREG_FILE_26xx16x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx16x, ZN
                           => n4732);
   U5289 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx16x,
                           B1 => n5120, B2 => fromRegsPortxREG_FILE_24xx16x, ZN
                           => n4731);
   U5290 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx16x,
                           B1 => n5054, B2 => fromRegsPortxREG_FILE_31xx16x, ZN
                           => n4730);
   U5291 : NAND4_X1 port map( A1 => n4733, A2 => n4732, A3 => n4731, A4 => 
                           n4730, ZN => n4739);
   U5292 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx16x,
                           B1 => n5126, B2 => fromRegsPortxREG_FILE_23xx16x, ZN
                           => n4737);
   U5293 : AOI22_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx16x,
                           B1 => n5187, B2 => fromRegsPortxREG_FILE_19xx16x, ZN
                           => n4736);
   U5294 : AOI22_X1 port map( A1 => n5093, A2 => fromRegsPortxREG_FILE_18xx16x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx16x, ZN
                           => n4735);
   U5295 : NAND2_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx16x,
                           ZN => n4734);
   U5296 : NAND4_X1 port map( A1 => n4737, A2 => n4736, A3 => n4735, A4 => 
                           n4734, ZN => n4738);
   U5297 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4739
                           , A => n4738, ZN => n4745);
   U5298 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx16x,
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx16x, ZN
                           => n4744);
   U5299 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_11xx16x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx16x, ZN
                           => n4741);
   U5300 : AOI22_X1 port map( A1 => n5301, A2 => fromRegsPortxREG_FILE_12xx16x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx16x, ZN
                           => n4740);
   U5301 : NAND2_X1 port map( A1 => n4741, A2 => n4740, ZN => n4742);
   U5302 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx16x, B2 => n5165,
                           A => n4742, ZN => n4743);
   U5303 : OAI211_X1 port map( C1 => n4745, C2 => n5200, A => n4744, B => n4743
                           , ZN => n4746);
   U5304 : NAND2_X1 port map( A1 => n4746, A2 => n5238, ZN => n4756);
   U5305 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx16x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx16x, ZN
                           => n4750);
   U5306 : AOI22_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx16x,
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx16x, ZN
                           => n4749);
   U5307 : AOI22_X1 port map( A1 => n5203, A2 => fromRegsPortxREG_FILE_09xx16x,
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx16x, ZN
                           => n4748);
   U5308 : NAND2_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx16x,
                           ZN => n4747);
   U5309 : NAND4_X1 port map( A1 => n4750, A2 => n4749, A3 => n4748, A4 => 
                           n4747, ZN => n4754);
   U5310 : NAND2_X1 port map( A1 => n4867, A2 => fromRegsPortxREG_FILE_02xx16x,
                           ZN => n4752);
   U5311 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx16x, A2 => n5244,
                           ZN => n4751);
   U5312 : NAND2_X1 port map( A1 => n4752, A2 => n4751, ZN => n4753);
   U5313 : AOI21_X1 port map( B1 => n4754, B2 => n5047, A => n4753, ZN => n4755
                           );
   U5314 : NAND2_X1 port map( A1 => n4756, A2 => n4755, ZN => n6805);
   U5315 : INV_X1 port map( A => n6805, ZN => n7468);
   U5316 : OAI22_X1 port map( A1 => n5673, A2 => n6811, B1 => n5674, B2 => 
                           n7468, ZN => n4757);
   U5317 : XOR2_X1 port map( A => n7546, B => n4757, Z => 
                           DP_OP_719J1_125_1055xn52);
   U5318 : NAND2_X1 port map( A1 => n5650, A2 => fromMemoryPortxLOADEDDATAx(15)
                           , ZN => n4758);
   U5319 : NAND2_X1 port map( A1 => n5652, A2 => n4758, ZN => add_x_26xBx15x);
   U5320 : INV_X1 port map( A => add_x_26xBx15x, ZN => n6778);
   U5321 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx15x,
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_27xx15x, ZN
                           => n4762);
   U5322 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx15x,
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_24xx15x, ZN
                           => n4761);
   U5323 : AOI22_X1 port map( A1 => n5087, A2 => fromRegsPortxREG_FILE_26xx15x,
                           B1 => n5085, B2 => fromRegsPortxREG_FILE_28xx15x, ZN
                           => n4760);
   U5324 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx15x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx15x, ZN
                           => n4759);
   U5325 : NAND4_X1 port map( A1 => n4762, A2 => n4761, A3 => n4760, A4 => 
                           n4759, ZN => n4768);
   U5326 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx15x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx15x, ZN
                           => n4766);
   U5327 : AOI22_X1 port map( A1 => n5092, A2 => fromRegsPortxREG_FILE_20xx15x,
                           B1 => n5126, B2 => fromRegsPortxREG_FILE_23xx15x, ZN
                           => n4765);
   U5328 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_19xx15x,
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx15x, ZN
                           => n4764);
   U5329 : NAND2_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx15x,
                           ZN => n4763);
   U5330 : NAND4_X1 port map( A1 => n4766, A2 => n4765, A3 => n4764, A4 => 
                           n4763, ZN => n4767);
   U5331 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4768
                           , A => n4767, ZN => n4774);
   U5332 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx15x,
                           B1 => n5065, B2 => fromRegsPortxREG_FILE_16xx15x, ZN
                           => n4773);
   U5333 : AOI22_X1 port map( A1 => n5102, A2 => fromRegsPortxREG_FILE_14xx15x,
                           B1 => n5303, B2 => fromRegsPortxREG_FILE_11xx15x, ZN
                           => n4770);
   U5334 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_13xx15x,
                           B1 => n5100, B2 => fromRegsPortxREG_FILE_15xx15x, ZN
                           => n4769);
   U5335 : NAND2_X1 port map( A1 => n4770, A2 => n4769, ZN => n4771);
   U5336 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx15x, B2 => n5301,
                           A => n4771, ZN => n4772);
   U5337 : OAI211_X1 port map( C1 => n4774, C2 => n5758, A => n4773, B => n4772
                           , ZN => n4775);
   U5338 : NAND2_X1 port map( A1 => n4775, A2 => n5238, ZN => n4785);
   U5339 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx15x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx15x, ZN
                           => n4779);
   U5340 : AOI22_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx15x,
                           B1 => n5039, B2 => fromRegsPortxREG_FILE_08xx15x, ZN
                           => n4778);
   U5341 : AOI22_X1 port map( A1 => n5073, A2 => fromRegsPortxREG_FILE_04xx15x,
                           B1 => n5010, B2 => fromRegsPortxREG_FILE_05xx15x, ZN
                           => n4777);
   U5342 : NAND2_X1 port map( A1 => n5142, A2 => fromRegsPortxREG_FILE_03xx15x,
                           ZN => n4776);
   U5343 : NAND4_X1 port map( A1 => n4779, A2 => n4778, A3 => n4777, A4 => 
                           n4776, ZN => n4783);
   U5344 : NAND2_X1 port map( A1 => n4867, A2 => fromRegsPortxREG_FILE_02xx15x,
                           ZN => n4781);
   U5345 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx15x, A2 => n5244,
                           ZN => n4780);
   U5346 : NAND2_X1 port map( A1 => n4781, A2 => n4780, ZN => n4782);
   U5347 : AOI21_X1 port map( B1 => n4783, B2 => n5047, A => n4782, ZN => n4784
                           );
   U5348 : NAND2_X1 port map( A1 => n4785, A2 => n4784, ZN => n6774);
   U5349 : INV_X1 port map( A => n6774, ZN => n7467);
   U5350 : OAI22_X1 port map( A1 => n5673, A2 => n6778, B1 => n5674, B2 => 
                           n7467, ZN => n4786);
   U5351 : XOR2_X1 port map( A => n5252, B => n4786, Z => 
                           DP_OP_719J1_125_1055xn53);
   U5352 : NAND2_X1 port map( A1 => n5650, A2 => fromMemoryPortxLOADEDDATAx(14)
                           , ZN => n4787);
   U5353 : NAND2_X1 port map( A1 => n5652, A2 => n4787, ZN => add_x_26xBx14x);
   U5354 : INV_X1 port map( A => add_x_26xBx14x, ZN => intadd_2xBx3x);
   U5355 : AOI22_X1 port map( A1 => n5086, A2 => fromRegsPortxREG_FILE_30xx14x,
                           B1 => n5276, B2 => fromRegsPortxREG_FILE_25xx14x, ZN
                           => n4791);
   U5356 : AOI22_X1 port map( A1 => n5087, A2 => fromRegsPortxREG_FILE_26xx14x,
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_24xx14x, ZN
                           => n4790);
   U5357 : AOI22_X1 port map( A1 => n5053, A2 => fromRegsPortxREG_FILE_29xx14x,
                           B1 => n5085, B2 => fromRegsPortxREG_FILE_28xx14x, ZN
                           => n4789);
   U5358 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_27xx14x,
                           B1 => n5054, B2 => fromRegsPortxREG_FILE_31xx14x, ZN
                           => n4788);
   U5359 : NAND4_X1 port map( A1 => n4791, A2 => n4790, A3 => n4789, A4 => 
                           n4788, ZN => n4797);
   U5360 : AOI22_X1 port map( A1 => n5093, A2 => fromRegsPortxREG_FILE_18xx14x,
                           B1 => n5187, B2 => fromRegsPortxREG_FILE_19xx14x, ZN
                           => n4795);
   U5361 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_21xx14x,
                           B1 => n5125, B2 => fromRegsPortxREG_FILE_17xx14x, ZN
                           => n4794);
   U5362 : AOI22_X1 port map( A1 => n5126, A2 => fromRegsPortxREG_FILE_23xx14x,
                           B1 => n5287, B2 => fromRegsPortxREG_FILE_22xx14x, ZN
                           => n4793);
   U5363 : NAND2_X1 port map( A1 => n5092, A2 => fromRegsPortxREG_FILE_20xx14x,
                           ZN => n4792);
   U5364 : NAND4_X1 port map( A1 => n4795, A2 => n4794, A3 => n4793, A4 => 
                           n4792, ZN => n4796);
   U5365 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4797
                           , A => n4796, ZN => n4803);
   U5366 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx14x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx14x, ZN
                           => n4802);
   U5367 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx14x,
                           B1 => n5100, B2 => fromRegsPortxREG_FILE_15xx14x, ZN
                           => n4799);
   U5368 : AOI22_X1 port map( A1 => n5101, A2 => fromRegsPortxREG_FILE_11xx14x,
                           B1 => n5065, B2 => fromRegsPortxREG_FILE_16xx14x, ZN
                           => n4798);
   U5369 : NAND2_X1 port map( A1 => n4799, A2 => n4798, ZN => n4800);
   U5370 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx14x, B2 => n5301,
                           A => n4800, ZN => n4801);
   U5371 : OAI211_X1 port map( C1 => n4803, C2 => n5758, A => n4802, B => n4801
                           , ZN => n4804);
   U5372 : NAND2_X1 port map( A1 => n4804, A2 => n5238, ZN => n4814);
   U5373 : AOI22_X1 port map( A1 => n5010, A2 => fromRegsPortxREG_FILE_05xx14x,
                           B1 => n5140, B2 => fromRegsPortxREG_FILE_07xx14x, ZN
                           => n4808);
   U5374 : AOI22_X1 port map( A1 => n5073, A2 => fromRegsPortxREG_FILE_04xx14x,
                           B1 => n5141, B2 => fromRegsPortxREG_FILE_06xx14x, ZN
                           => n4807);
   U5375 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx14x,
                           B1 => n5039, B2 => fromRegsPortxREG_FILE_08xx14x, ZN
                           => n4806);
   U5376 : NAND2_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx14x,
                           ZN => n4805);
   U5377 : NAND4_X1 port map( A1 => n4808, A2 => n4807, A3 => n4806, A4 => 
                           n4805, ZN => n4812);
   U5378 : NAND2_X1 port map( A1 => n4867, A2 => fromRegsPortxREG_FILE_02xx14x,
                           ZN => n4810);
   U5379 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx14x, A2 => n5244,
                           ZN => n4809);
   U5380 : NAND2_X1 port map( A1 => n4810, A2 => n4809, ZN => n4811);
   U5381 : AOI21_X1 port map( B1 => n4812, B2 => n5047, A => n4811, ZN => n4813
                           );
   U5382 : NAND2_X1 port map( A1 => n4814, A2 => n4813, ZN => n6726);
   U5383 : INV_X1 port map( A => n6726, ZN => n7466);
   U5384 : OAI22_X1 port map( A1 => n5673, A2 => intadd_2xBx3x, B1 => n5674, B2
                           => n7466, ZN => n4815);
   U5385 : XOR2_X1 port map( A => n5252, B => n4815, Z => 
                           DP_OP_719J1_125_1055xn54);
   U5386 : NAND2_X1 port map( A1 => n5650, A2 => fromMemoryPortxLOADEDDATAx(13)
                           , ZN => n4816);
   U5387 : NAND2_X1 port map( A1 => n5652, A2 => n4816, ZN => add_x_26xBx13x);
   U5388 : INV_X1 port map( A => add_x_26xBx13x, ZN => intadd_2xBx2x);
   U5389 : AOI22_X1 port map( A1 => n5276, A2 => fromRegsPortxREG_FILE_25xx13x,
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_27xx13x, ZN
                           => n4820);
   U5390 : AOI22_X1 port map( A1 => n5086, A2 => fromRegsPortxREG_FILE_30xx13x,
                           B1 => n5087, B2 => fromRegsPortxREG_FILE_26xx13x, ZN
                           => n4819);
   U5391 : AOI22_X1 port map( A1 => n5053, A2 => fromRegsPortxREG_FILE_29xx13x,
                           B1 => n5085, B2 => fromRegsPortxREG_FILE_28xx13x, ZN
                           => n4818);
   U5392 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_24xx13x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx13x, ZN
                           => n4817);
   U5393 : NAND4_X1 port map( A1 => n4820, A2 => n4819, A3 => n4818, A4 => 
                           n4817, ZN => n4826);
   U5394 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx13x,
                           B1 => n5125, B2 => fromRegsPortxREG_FILE_17xx13x, ZN
                           => n4824);
   U5395 : AOI22_X1 port map( A1 => n5092, A2 => fromRegsPortxREG_FILE_20xx13x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx13x, ZN
                           => n4823);
   U5396 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_21xx13x,
                           B1 => n5187, B2 => fromRegsPortxREG_FILE_19xx13x, ZN
                           => n4822);
   U5397 : NAND2_X1 port map( A1 => n5126, A2 => fromRegsPortxREG_FILE_23xx13x,
                           ZN => n4821);
   U5398 : NAND4_X1 port map( A1 => n4824, A2 => n4823, A3 => n4822, A4 => 
                           n4821, ZN => n4825);
   U5399 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4826
                           , A => n4825, ZN => n4832);
   U5400 : AOI22_X1 port map( A1 => n5065, A2 => fromRegsPortxREG_FILE_16xx13x,
                           B1 => n5100, B2 => fromRegsPortxREG_FILE_15xx13x, ZN
                           => n4831);
   U5401 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx13x,
                           B1 => n5101, B2 => fromRegsPortxREG_FILE_11xx13x, ZN
                           => n4828);
   U5402 : AOI22_X1 port map( A1 => n5301, A2 => fromRegsPortxREG_FILE_12xx13x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx13x, ZN
                           => n4827);
   U5403 : NAND2_X1 port map( A1 => n4828, A2 => n4827, ZN => n4829);
   U5404 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx13x, B2 => n5300,
                           A => n4829, ZN => n4830);
   U5405 : OAI211_X1 port map( C1 => n4832, C2 => n5758, A => n4831, B => n4830
                           , ZN => n4833);
   U5406 : NAND2_X1 port map( A1 => n4833, A2 => n5238, ZN => n4843);
   U5407 : AOI22_X1 port map( A1 => n5073, A2 => fromRegsPortxREG_FILE_04xx13x,
                           B1 => n5140, B2 => fromRegsPortxREG_FILE_07xx13x, ZN
                           => n4837);
   U5408 : AOI22_X1 port map( A1 => n5203, A2 => fromRegsPortxREG_FILE_09xx13x,
                           B1 => n5039, B2 => fromRegsPortxREG_FILE_08xx13x, ZN
                           => n4836);
   U5409 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx13x,
                           B1 => n5010, B2 => fromRegsPortxREG_FILE_05xx13x, ZN
                           => n4835);
   U5410 : NAND2_X1 port map( A1 => n5141, A2 => fromRegsPortxREG_FILE_06xx13x,
                           ZN => n4834);
   U5411 : NAND4_X1 port map( A1 => n4837, A2 => n4836, A3 => n4835, A4 => 
                           n4834, ZN => n4841);
   U5412 : NAND2_X1 port map( A1 => n4867, A2 => fromRegsPortxREG_FILE_02xx13x,
                           ZN => n4839);
   U5413 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx13x, A2 => n5244,
                           ZN => n4838);
   U5414 : NAND2_X1 port map( A1 => n4839, A2 => n4838, ZN => n4840);
   U5415 : AOI21_X1 port map( B1 => n4841, B2 => n5047, A => n4840, ZN => n4842
                           );
   U5416 : NAND2_X1 port map( A1 => n4843, A2 => n4842, ZN => n6702);
   U5417 : INV_X1 port map( A => n6702, ZN => n7465);
   U5418 : OAI22_X1 port map( A1 => n5673, A2 => intadd_2xBx2x, B1 => n5674, B2
                           => n7465, ZN => n4844);
   U5419 : XOR2_X1 port map( A => n7546, B => n4844, Z => 
                           DP_OP_719J1_125_1055xn55);
   U5420 : NAND2_X1 port map( A1 => n5650, A2 => fromMemoryPortxLOADEDDATAx(12)
                           , ZN => n4845);
   U5421 : NAND2_X1 port map( A1 => n5652, A2 => n4845, ZN => add_x_26xBx12x);
   U5422 : INV_X1 port map( A => add_x_26xBx12x, ZN => intadd_2xBx1x);
   U5423 : AOI22_X1 port map( A1 => n5086, A2 => fromRegsPortxREG_FILE_30xx12x,
                           B1 => n5087, B2 => fromRegsPortxREG_FILE_26xx12x, ZN
                           => n4849);
   U5424 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_27xx12x,
                           B1 => n5085, B2 => fromRegsPortxREG_FILE_28xx12x, ZN
                           => n4848);
   U5425 : AOI22_X1 port map( A1 => n5182, A2 => fromRegsPortxREG_FILE_25xx12x,
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_29xx12x, ZN
                           => n4847);
   U5426 : AOI22_X1 port map( A1 => n5120, A2 => fromRegsPortxREG_FILE_24xx12x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx12x, ZN
                           => n4846);
   U5427 : NAND4_X1 port map( A1 => n4849, A2 => n4848, A3 => n4847, A4 => 
                           n4846, ZN => n4855);
   U5428 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_19xx12x,
                           B1 => n5125, B2 => fromRegsPortxREG_FILE_17xx12x, ZN
                           => n4853);
   U5429 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx12x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx12x, ZN
                           => n4852);
   U5430 : AOI22_X1 port map( A1 => n5092, A2 => fromRegsPortxREG_FILE_20xx12x,
                           B1 => n5126, B2 => fromRegsPortxREG_FILE_23xx12x, ZN
                           => n4851);
   U5431 : NAND2_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_21xx12x,
                           ZN => n4850);
   U5432 : NAND4_X1 port map( A1 => n4853, A2 => n4852, A3 => n4851, A4 => 
                           n4850, ZN => n4854);
   U5433 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4855
                           , A => n4854, ZN => n4861);
   U5434 : AOI22_X1 port map( A1 => n5101, A2 => fromRegsPortxREG_FILE_11xx12x,
                           B1 => n5065, B2 => fromRegsPortxREG_FILE_16xx12x, ZN
                           => n4860);
   U5435 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_10xx12x,
                           B1 => n5100, B2 => fromRegsPortxREG_FILE_15xx12x, ZN
                           => n4857);
   U5436 : AOI22_X1 port map( A1 => n5102, A2 => fromRegsPortxREG_FILE_14xx12x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx12x, ZN
                           => n4856);
   U5437 : NAND2_X1 port map( A1 => n4857, A2 => n4856, ZN => n4858);
   U5438 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx12x, B2 => n5234,
                           A => n4858, ZN => n4859);
   U5439 : OAI211_X1 port map( C1 => n4861, C2 => n5758, A => n4860, B => n4859
                           , ZN => n4862);
   U5440 : NAND2_X1 port map( A1 => n4862, A2 => n5238, ZN => n4873);
   U5441 : AOI22_X1 port map( A1 => n5203, A2 => fromRegsPortxREG_FILE_09xx12x,
                           B1 => n5140, B2 => fromRegsPortxREG_FILE_07xx12x, ZN
                           => n4866);
   U5442 : AOI22_X1 port map( A1 => n5073, A2 => fromRegsPortxREG_FILE_04xx12x,
                           B1 => n5141, B2 => fromRegsPortxREG_FILE_06xx12x, ZN
                           => n4865);
   U5443 : AOI22_X1 port map( A1 => n5039, A2 => fromRegsPortxREG_FILE_08xx12x,
                           B1 => n5010, B2 => fromRegsPortxREG_FILE_05xx12x, ZN
                           => n4864);
   U5444 : NAND2_X1 port map( A1 => n5142, A2 => fromRegsPortxREG_FILE_03xx12x,
                           ZN => n4863);
   U5445 : NAND4_X1 port map( A1 => n4866, A2 => n4865, A3 => n4864, A4 => 
                           n4863, ZN => n4871);
   U5446 : NAND2_X1 port map( A1 => n4867, A2 => fromRegsPortxREG_FILE_02xx12x,
                           ZN => n4869);
   U5447 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx12x, A2 => n5327,
                           ZN => n4868);
   U5448 : NAND2_X1 port map( A1 => n4869, A2 => n4868, ZN => n4870);
   U5449 : AOI21_X1 port map( B1 => n4871, B2 => n5047, A => n4870, ZN => n4872
                           );
   U5450 : NAND2_X1 port map( A1 => n4873, A2 => n4872, ZN => n6658);
   U5451 : INV_X1 port map( A => n6658, ZN => n7464);
   U5452 : OAI22_X1 port map( A1 => n7464, A2 => n5676, B1 => n5675, B2 => 
                           intadd_2xBx1x, ZN => n4874);
   U5453 : XOR2_X1 port map( A => n5252, B => n4874, Z => 
                           DP_OP_719J1_125_1055xn56);
   U5454 : NAND2_X1 port map( A1 => n4875, A2 => fromMemoryPortxLOADEDDATAx(7),
                           ZN => n4880);
   U5455 : INV_X1 port map( A => n4876, ZN => n4877);
   U5456 : OAI21_X1 port map( B1 => n5641, B2 => n6982, A => n4877, ZN => n4878
                           );
   U5457 : INV_X1 port map( A => n4878, ZN => n4879);
   U5458 : NAND2_X1 port map( A1 => n4880, A2 => n4879, ZN => add_x_26xBx11x);
   U5459 : INV_X1 port map( A => add_x_26xBx11x, ZN => intadd_2xBx0x);
   U5460 : AOI22_X1 port map( A1 => n5182, A2 => fromRegsPortxREG_FILE_25xx11x,
                           B1 => n5085, B2 => fromRegsPortxREG_FILE_28xx11x, ZN
                           => n4884);
   U5461 : AOI22_X1 port map( A1 => n5086, A2 => fromRegsPortxREG_FILE_30xx11x,
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx11x, ZN
                           => n4883);
   U5462 : AOI22_X1 port map( A1 => n5053, A2 => fromRegsPortxREG_FILE_29xx11x,
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_24xx11x, ZN
                           => n4882);
   U5463 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_27xx11x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx11x, ZN
                           => n4881);
   U5464 : NAND4_X1 port map( A1 => n4884, A2 => n4883, A3 => n4882, A4 => 
                           n4881, ZN => n4890);
   U5465 : AOI22_X1 port map( A1 => n5093, A2 => fromRegsPortxREG_FILE_18xx11x,
                           B1 => n5125, B2 => fromRegsPortxREG_FILE_17xx11x, ZN
                           => n4888);
   U5466 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_21xx11x,
                           B1 => n5187, B2 => fromRegsPortxREG_FILE_19xx11x, ZN
                           => n4887);
   U5467 : AOI22_X1 port map( A1 => n5126, A2 => fromRegsPortxREG_FILE_23xx11x,
                           B1 => n5287, B2 => fromRegsPortxREG_FILE_22xx11x, ZN
                           => n4886);
   U5468 : NAND2_X1 port map( A1 => n5092, A2 => fromRegsPortxREG_FILE_20xx11x,
                           ZN => n4885);
   U5469 : NAND4_X1 port map( A1 => n4888, A2 => n4887, A3 => n4886, A4 => 
                           n4885, ZN => n4889);
   U5470 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4890
                           , A => n4889, ZN => n4896);
   U5471 : AOI22_X1 port map( A1 => n5065, A2 => fromRegsPortxREG_FILE_16xx11x,
                           B1 => n5100, B2 => fromRegsPortxREG_FILE_15xx11x, ZN
                           => n4895);
   U5472 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_10xx11x,
                           B1 => n5101, B2 => fromRegsPortxREG_FILE_11xx11x, ZN
                           => n4892);
   U5473 : AOI22_X1 port map( A1 => n5102, A2 => fromRegsPortxREG_FILE_14xx11x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx11x, ZN
                           => n4891);
   U5474 : NAND2_X1 port map( A1 => n4892, A2 => n4891, ZN => n4893);
   U5475 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx11x, B2 => n5234,
                           A => n4893, ZN => n4894);
   U5476 : OAI211_X1 port map( C1 => n4896, C2 => n5758, A => n4895, B => n4894
                           , ZN => n4897);
   U5477 : CLKBUF_X1 port map( A => n5238, Z => n5313);
   U5478 : NAND2_X1 port map( A1 => n4897, A2 => n5313, ZN => n4907);
   U5479 : AOI22_X1 port map( A1 => n5073, A2 => fromRegsPortxREG_FILE_04xx11x,
                           B1 => n5142, B2 => fromRegsPortxREG_FILE_03xx11x, ZN
                           => n4901);
   U5480 : AOI22_X1 port map( A1 => n5203, A2 => fromRegsPortxREG_FILE_09xx11x,
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx11x, ZN
                           => n4900);
   U5481 : AOI22_X1 port map( A1 => n5039, A2 => fromRegsPortxREG_FILE_08xx11x,
                           B1 => n5140, B2 => fromRegsPortxREG_FILE_07xx11x, ZN
                           => n4899);
   U5482 : NAND2_X1 port map( A1 => n5141, A2 => fromRegsPortxREG_FILE_06xx11x,
                           ZN => n4898);
   U5483 : NAND4_X1 port map( A1 => n4901, A2 => n4900, A3 => n4899, A4 => 
                           n4898, ZN => n4905);
   U5484 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx11x,
                           ZN => n4903);
   U5485 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx11x, A2 => n5244,
                           ZN => n4902);
   U5486 : NAND2_X1 port map( A1 => n4903, A2 => n4902, ZN => n4904);
   U5487 : AOI21_X1 port map( B1 => n4905, B2 => n5047, A => n4904, ZN => n4906
                           );
   U5488 : NAND2_X1 port map( A1 => n4907, A2 => n4906, ZN => n6616);
   U5489 : INV_X1 port map( A => n6616, ZN => n7463);
   U5490 : OAI22_X1 port map( A1 => n5673, A2 => intadd_2xBx0x, B1 => n5674, B2
                           => n7463, ZN => n4908);
   U5491 : XOR2_X1 port map( A => n5252, B => n4908, Z => 
                           DP_OP_719J1_125_1055xn57);
   U5492 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(30), A2 => n5052,
                           ZN => add_x_26xBx10x);
   U5493 : INV_X1 port map( A => add_x_26xBx10x, ZN => n5835);
   U5494 : AOI22_X1 port map( A1 => n5182, A2 => fromRegsPortxREG_FILE_25xx10x,
                           B1 => n5087, B2 => fromRegsPortxREG_FILE_26xx10x, ZN
                           => n4912);
   U5495 : AOI22_X1 port map( A1 => n5086, A2 => fromRegsPortxREG_FILE_30xx10x,
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_27xx10x, ZN
                           => n4911);
   U5496 : AOI22_X1 port map( A1 => n5120, A2 => fromRegsPortxREG_FILE_24xx10x,
                           B1 => n5085, B2 => fromRegsPortxREG_FILE_28xx10x, ZN
                           => n4910);
   U5497 : AOI22_X1 port map( A1 => n5053, A2 => fromRegsPortxREG_FILE_29xx10x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx10x, ZN
                           => n4909);
   U5498 : NAND4_X1 port map( A1 => n4912, A2 => n4911, A3 => n4910, A4 => 
                           n4909, ZN => n4918);
   U5499 : AOI22_X1 port map( A1 => n5092, A2 => fromRegsPortxREG_FILE_20xx10x,
                           B1 => n5287, B2 => fromRegsPortxREG_FILE_22xx10x, ZN
                           => n4916);
   U5500 : AOI22_X1 port map( A1 => n5126, A2 => fromRegsPortxREG_FILE_23xx10x,
                           B1 => n5187, B2 => fromRegsPortxREG_FILE_19xx10x, ZN
                           => n4915);
   U5501 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_21xx10x,
                           B1 => n5125, B2 => fromRegsPortxREG_FILE_17xx10x, ZN
                           => n4914);
   U5502 : NAND2_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_18xx10x,
                           ZN => n4913);
   U5503 : NAND4_X1 port map( A1 => n4916, A2 => n4915, A3 => n4914, A4 => 
                           n4913, ZN => n4917);
   U5504 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4918
                           , A => n4917, ZN => n4924);
   U5505 : AOI22_X1 port map( A1 => n5101, A2 => fromRegsPortxREG_FILE_11xx10x,
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx10x, ZN
                           => n4923);
   U5506 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_10xx10x,
                           B1 => n5100, B2 => fromRegsPortxREG_FILE_15xx10x, ZN
                           => n4920);
   U5507 : AOI22_X1 port map( A1 => n5102, A2 => fromRegsPortxREG_FILE_14xx10x,
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx10x, ZN
                           => n4919);
   U5508 : NAND2_X1 port map( A1 => n4920, A2 => n4919, ZN => n4921);
   U5509 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx10x, B2 => n5234,
                           A => n4921, ZN => n4922);
   U5510 : OAI211_X1 port map( C1 => n4924, C2 => n5758, A => n4923, B => n4922
                           , ZN => n4925);
   U5511 : NAND2_X1 port map( A1 => n4925, A2 => n5313, ZN => n4935);
   U5512 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx10x,
                           B1 => n5010, B2 => fromRegsPortxREG_FILE_05xx10x, ZN
                           => n4929);
   U5513 : AOI22_X1 port map( A1 => n5141, A2 => fromRegsPortxREG_FILE_06xx10x,
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx10x, ZN
                           => n4928);
   U5514 : AOI22_X1 port map( A1 => n5073, A2 => fromRegsPortxREG_FILE_04xx10x,
                           B1 => n5140, B2 => fromRegsPortxREG_FILE_07xx10x, ZN
                           => n4927);
   U5515 : NAND2_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx10x,
                           ZN => n4926);
   U5516 : NAND4_X1 port map( A1 => n4929, A2 => n4928, A3 => n4927, A4 => 
                           n4926, ZN => n4933);
   U5517 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx10x,
                           ZN => n4931);
   U5518 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx10x, A2 => n5327,
                           ZN => n4930);
   U5519 : NAND2_X1 port map( A1 => n4931, A2 => n4930, ZN => n4932);
   U5520 : AOI21_X1 port map( B1 => n4933, B2 => n5047, A => n4932, ZN => n4934
                           );
   U5521 : NAND2_X1 port map( A1 => n4935, A2 => n4934, ZN => n6555);
   U5522 : INV_X1 port map( A => n6555, ZN => n7462);
   U5523 : OAI22_X1 port map( A1 => n5673, A2 => n5835, B1 => n5674, B2 => 
                           n7462, ZN => n4936);
   U5524 : XOR2_X1 port map( A => n7546, B => n4936, Z => 
                           DP_OP_719J1_125_1055xn58);
   U5525 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(29), A2 => n5052,
                           ZN => add_x_26xBx9x);
   U5526 : AOI22_X1 port map( A1 => n5053, A2 => fromRegsPortxREG_FILE_29xx9x, 
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_27xx9x, ZN 
                           => n4940);
   U5527 : AOI22_X1 port map( A1 => n5182, A2 => fromRegsPortxREG_FILE_25xx9x, 
                           B1 => n5085, B2 => fromRegsPortxREG_FILE_28xx9x, ZN 
                           => n4939);
   U5528 : AOI22_X1 port map( A1 => n5086, A2 => fromRegsPortxREG_FILE_30xx9x, 
                           B1 => n5087, B2 => fromRegsPortxREG_FILE_26xx9x, ZN 
                           => n4938);
   U5529 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_24xx9x, 
                           B1 => n5054, B2 => fromRegsPortxREG_FILE_31xx9x, ZN 
                           => n4937);
   U5530 : NAND4_X1 port map( A1 => n4940, A2 => n4939, A3 => n4938, A4 => 
                           n4937, ZN => n4946);
   U5531 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_21xx9x, 
                           B1 => n5125, B2 => fromRegsPortxREG_FILE_17xx9x, ZN 
                           => n4944);
   U5532 : AOI22_X1 port map( A1 => n5093, A2 => fromRegsPortxREG_FILE_18xx9x, 
                           B1 => n5187, B2 => fromRegsPortxREG_FILE_19xx9x, ZN 
                           => n4943);
   U5533 : AOI22_X1 port map( A1 => n5126, A2 => fromRegsPortxREG_FILE_23xx9x, 
                           B1 => n5287, B2 => fromRegsPortxREG_FILE_22xx9x, ZN 
                           => n4942);
   U5534 : NAND2_X1 port map( A1 => n5092, A2 => fromRegsPortxREG_FILE_20xx9x, 
                           ZN => n4941);
   U5535 : NAND4_X1 port map( A1 => n4944, A2 => n4943, A3 => n4942, A4 => 
                           n4941, ZN => n4945);
   U5536 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4946
                           , A => n4945, ZN => n4952);
   U5537 : AOI22_X1 port map( A1 => n5102, A2 => fromRegsPortxREG_FILE_14xx9x, 
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx9x, ZN 
                           => n4951);
   U5538 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx9x, 
                           B1 => n5100, B2 => fromRegsPortxREG_FILE_15xx9x, ZN 
                           => n4948);
   U5539 : AOI22_X1 port map( A1 => n5101, A2 => fromRegsPortxREG_FILE_11xx9x, 
                           B1 => n5065, B2 => fromRegsPortxREG_FILE_16xx9x, ZN 
                           => n4947);
   U5540 : NAND2_X1 port map( A1 => n4948, A2 => n4947, ZN => n4949);
   U5541 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx9x, B2 => n5301, 
                           A => n4949, ZN => n4950);
   U5542 : OAI211_X1 port map( C1 => n4952, C2 => n5758, A => n4951, B => n4950
                           , ZN => n4953);
   U5543 : NAND2_X1 port map( A1 => n4953, A2 => n5313, ZN => n4963);
   U5544 : AOI22_X1 port map( A1 => n5039, A2 => fromRegsPortxREG_FILE_08xx9x, 
                           B1 => n5140, B2 => fromRegsPortxREG_FILE_07xx9x, ZN 
                           => n4957);
   U5545 : AOI22_X1 port map( A1 => n5073, A2 => fromRegsPortxREG_FILE_04xx9x, 
                           B1 => n5010, B2 => fromRegsPortxREG_FILE_05xx9x, ZN 
                           => n4956);
   U5546 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx9x, 
                           B1 => n5141, B2 => fromRegsPortxREG_FILE_06xx9x, ZN 
                           => n4955);
   U5547 : NAND2_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx9x, 
                           ZN => n4954);
   U5548 : NAND4_X1 port map( A1 => n4957, A2 => n4956, A3 => n4955, A4 => 
                           n4954, ZN => n4961);
   U5549 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx9x, 
                           ZN => n4959);
   U5550 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx9x, A2 => n5327, 
                           ZN => n4958);
   U5551 : NAND2_X1 port map( A1 => n4959, A2 => n4958, ZN => n4960);
   U5552 : AOI21_X1 port map( B1 => n4961, B2 => n5047, A => n4960, ZN => n4962
                           );
   U5553 : NAND2_X1 port map( A1 => n4963, A2 => n4962, ZN => n6504);
   U5554 : INV_X1 port map( A => n6504, ZN => n7461);
   U5555 : INV_X1 port map( A => add_x_26xBx9x, ZN => n6500);
   U5556 : OAI22_X1 port map( A1 => n7461, A2 => n5674, B1 => n5675, B2 => 
                           n6500, ZN => n4964);
   U5557 : XOR2_X1 port map( A => n5252, B => n4964, Z => 
                           DP_OP_719J1_125_1055xn59);
   U5558 : INV_X1 port map( A => add_x_26xBx8x, ZN => n5586);
   U5559 : AOI22_X1 port map( A1 => n5120, A2 => fromRegsPortxREG_FILE_24xx8x, 
                           B1 => n5085, B2 => fromRegsPortxREG_FILE_28xx8x, ZN 
                           => n4968);
   U5560 : AOI22_X1 port map( A1 => n5086, A2 => fromRegsPortxREG_FILE_30xx8x, 
                           B1 => n5087, B2 => fromRegsPortxREG_FILE_26xx8x, ZN 
                           => n4967);
   U5561 : AOI22_X1 port map( A1 => n5053, A2 => fromRegsPortxREG_FILE_29xx8x, 
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_27xx8x, ZN 
                           => n4966);
   U5562 : AOI22_X1 port map( A1 => n5182, A2 => fromRegsPortxREG_FILE_25xx8x, 
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx8x, ZN 
                           => n4965);
   U5563 : NAND4_X1 port map( A1 => n4968, A2 => n4967, A3 => n4966, A4 => 
                           n4965, ZN => n4974);
   U5564 : AOI22_X1 port map( A1 => n5092, A2 => fromRegsPortxREG_FILE_20xx8x, 
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx8x, ZN 
                           => n4972);
   U5565 : AOI22_X1 port map( A1 => n5126, A2 => fromRegsPortxREG_FILE_23xx8x, 
                           B1 => n5125, B2 => fromRegsPortxREG_FILE_17xx8x, ZN 
                           => n4971);
   U5566 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx8x, 
                           B1 => n5187, B2 => fromRegsPortxREG_FILE_19xx8x, ZN 
                           => n4970);
   U5567 : NAND2_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_21xx8x, 
                           ZN => n4969);
   U5568 : NAND4_X1 port map( A1 => n4972, A2 => n4971, A3 => n4970, A4 => 
                           n4969, ZN => n4973);
   U5569 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4974
                           , A => n4973, ZN => n4980);
   U5570 : AOI22_X1 port map( A1 => n5102, A2 => fromRegsPortxREG_FILE_14xx8x, 
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx8x, ZN 
                           => n4979);
   U5571 : AOI22_X1 port map( A1 => n5101, A2 => fromRegsPortxREG_FILE_11xx8x, 
                           B1 => n5100, B2 => fromRegsPortxREG_FILE_15xx8x, ZN 
                           => n4976);
   U5572 : AOI22_X1 port map( A1 => n5301, A2 => fromRegsPortxREG_FILE_12xx8x, 
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx8x, ZN 
                           => n4975);
   U5573 : NAND2_X1 port map( A1 => n4976, A2 => n4975, ZN => n4977);
   U5574 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx8x, B2 => n5300, 
                           A => n4977, ZN => n4978);
   U5575 : OAI211_X1 port map( C1 => n4980, C2 => n5758, A => n4979, B => n4978
                           , ZN => n4981);
   U5576 : NAND2_X1 port map( A1 => n4981, A2 => n5313, ZN => n4991);
   U5577 : AOI22_X1 port map( A1 => n5203, A2 => fromRegsPortxREG_FILE_09xx8x, 
                           B1 => n5142, B2 => fromRegsPortxREG_FILE_03xx8x, ZN 
                           => n4985);
   U5578 : AOI22_X1 port map( A1 => n5073, A2 => fromRegsPortxREG_FILE_04xx8x, 
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx8x, ZN 
                           => n4984);
   U5579 : AOI22_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx8x, 
                           B1 => n5140, B2 => fromRegsPortxREG_FILE_07xx8x, ZN 
                           => n4983);
   U5580 : NAND2_X1 port map( A1 => n5010, A2 => fromRegsPortxREG_FILE_05xx8x, 
                           ZN => n4982);
   U5581 : NAND4_X1 port map( A1 => n4985, A2 => n4984, A3 => n4983, A4 => 
                           n4982, ZN => n4989);
   U5582 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx8x, 
                           ZN => n4987);
   U5583 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx8x, A2 => n5327, 
                           ZN => n4986);
   U5584 : NAND2_X1 port map( A1 => n4987, A2 => n4986, ZN => n4988);
   U5585 : AOI21_X1 port map( B1 => n4989, B2 => n5047, A => n4988, ZN => n4990
                           );
   U5586 : NAND2_X1 port map( A1 => n4991, A2 => n4990, ZN => n6445);
   U5587 : INV_X1 port map( A => n6445, ZN => n7460);
   U5588 : OAI22_X1 port map( A1 => n5675, A2 => n5586, B1 => n5674, B2 => 
                           n7460, ZN => n4992);
   U5589 : XOR2_X1 port map( A => n5252, B => n4992, Z => 
                           DP_OP_719J1_125_1055xn60);
   U5590 : INV_X1 port map( A => add_x_26xBx7x, ZN => n6420);
   U5591 : AOI22_X1 port map( A1 => n5182, A2 => fromRegsPortxREG_FILE_25xx7x, 
                           B1 => n5085, B2 => fromRegsPortxREG_FILE_28xx7x, ZN 
                           => n4996);
   U5592 : AOI22_X1 port map( A1 => n5087, A2 => fromRegsPortxREG_FILE_26xx7x, 
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_27xx7x, ZN 
                           => n4995);
   U5593 : AOI22_X1 port map( A1 => n5086, A2 => fromRegsPortxREG_FILE_30xx7x, 
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_29xx7x, ZN 
                           => n4994);
   U5594 : AOI22_X1 port map( A1 => n5120, A2 => fromRegsPortxREG_FILE_24xx7x, 
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx7x, ZN 
                           => n4993);
   U5595 : NAND4_X1 port map( A1 => n4996, A2 => n4995, A3 => n4994, A4 => 
                           n4993, ZN => n5002);
   U5596 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx7x, 
                           B1 => n5288, B2 => fromRegsPortxREG_FILE_21xx7x, ZN 
                           => n5000);
   U5597 : AOI22_X1 port map( A1 => n5093, A2 => fromRegsPortxREG_FILE_18xx7x, 
                           B1 => n5125, B2 => fromRegsPortxREG_FILE_17xx7x, ZN 
                           => n4999);
   U5598 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx7x, 
                           B1 => n5187, B2 => fromRegsPortxREG_FILE_19xx7x, ZN 
                           => n4998);
   U5599 : NAND2_X1 port map( A1 => n5287, A2 => fromRegsPortxREG_FILE_22xx7x, 
                           ZN => n4997);
   U5600 : NAND4_X1 port map( A1 => n5000, A2 => n4999, A3 => n4998, A4 => 
                           n4997, ZN => n5001);
   U5601 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5002
                           , A => n5001, ZN => n5008);
   U5602 : AOI22_X1 port map( A1 => n5301, A2 => fromRegsPortxREG_FILE_12xx7x, 
                           B1 => n5100, B2 => fromRegsPortxREG_FILE_15xx7x, ZN 
                           => n5007);
   U5603 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_10xx7x, 
                           B1 => n5101, B2 => fromRegsPortxREG_FILE_11xx7x, ZN 
                           => n5004);
   U5604 : AOI22_X1 port map( A1 => n5065, A2 => fromRegsPortxREG_FILE_16xx7x, 
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx7x, ZN 
                           => n5003);
   U5605 : NAND2_X1 port map( A1 => n5004, A2 => n5003, ZN => n5005);
   U5606 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_14xx7x, B2 => n5102, 
                           A => n5005, ZN => n5006);
   U5607 : OAI211_X1 port map( C1 => n5008, C2 => n5200, A => n5007, B => n5006
                           , ZN => n5009);
   U5608 : NAND2_X1 port map( A1 => n5009, A2 => n5313, ZN => n5020);
   U5609 : AOI22_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx7x, 
                           B1 => n5140, B2 => fromRegsPortxREG_FILE_07xx7x, ZN 
                           => n5014);
   U5610 : AOI22_X1 port map( A1 => n5203, A2 => fromRegsPortxREG_FILE_09xx7x, 
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx7x, ZN 
                           => n5013);
   U5611 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx7x, 
                           B1 => n5142, B2 => fromRegsPortxREG_FILE_03xx7x, ZN 
                           => n5012);
   U5612 : NAND2_X1 port map( A1 => n5010, A2 => fromRegsPortxREG_FILE_05xx7x, 
                           ZN => n5011);
   U5613 : NAND4_X1 port map( A1 => n5014, A2 => n5013, A3 => n5012, A4 => 
                           n5011, ZN => n5018);
   U5614 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx7x, 
                           ZN => n5016);
   U5615 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx7x, A2 => n5327, 
                           ZN => n5015);
   U5616 : NAND2_X1 port map( A1 => n5016, A2 => n5015, ZN => n5017);
   U5617 : AOI21_X1 port map( B1 => n5018, B2 => n5047, A => n5017, ZN => n5019
                           );
   U5618 : NAND2_X1 port map( A1 => n5020, A2 => n5019, ZN => n6406);
   U5619 : INV_X1 port map( A => n6406, ZN => n7459);
   U5620 : OAI22_X1 port map( A1 => n5675, A2 => n6420, B1 => n5674, B2 => 
                           n7459, ZN => n5021);
   U5621 : XOR2_X1 port map( A => n7546, B => n5021, Z => 
                           DP_OP_719J1_125_1055xn61);
   U5622 : AOI22_X1 port map( A1 => n5086, A2 => fromRegsPortxREG_FILE_30xx6x, 
                           B1 => n5085, B2 => fromRegsPortxREG_FILE_28xx6x, ZN 
                           => n5025);
   U5623 : AOI22_X1 port map( A1 => n5120, A2 => fromRegsPortxREG_FILE_24xx6x, 
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_27xx6x, ZN 
                           => n5024);
   U5624 : AOI22_X1 port map( A1 => n5182, A2 => fromRegsPortxREG_FILE_25xx6x, 
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx6x, ZN 
                           => n5023);
   U5625 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx6x, 
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx6x, ZN 
                           => n5022);
   U5626 : NAND4_X1 port map( A1 => n5025, A2 => n5024, A3 => n5023, A4 => 
                           n5022, ZN => n5031);
   U5627 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx6x, 
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx6x, ZN 
                           => n5029);
   U5628 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx6x, 
                           B1 => n5288, B2 => fromRegsPortxREG_FILE_21xx6x, ZN 
                           => n5028);
   U5629 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_19xx6x, 
                           B1 => n5125, B2 => fromRegsPortxREG_FILE_17xx6x, ZN 
                           => n5027);
   U5630 : NAND2_X1 port map( A1 => n5287, A2 => fromRegsPortxREG_FILE_22xx6x, 
                           ZN => n5026);
   U5631 : NAND4_X1 port map( A1 => n5029, A2 => n5028, A3 => n5027, A4 => 
                           n5026, ZN => n5030);
   U5632 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5031
                           , A => n5030, ZN => n5037);
   U5633 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx6x, 
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx6x, ZN 
                           => n5036);
   U5634 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_10xx6x, 
                           B1 => n5101, B2 => fromRegsPortxREG_FILE_11xx6x, ZN 
                           => n5033);
   U5635 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_13xx6x, 
                           B1 => n5100, B2 => fromRegsPortxREG_FILE_15xx6x, ZN 
                           => n5032);
   U5636 : NAND2_X1 port map( A1 => n5033, A2 => n5032, ZN => n5034);
   U5637 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx6x, B2 => n5234, 
                           A => n5034, ZN => n5035);
   U5638 : OAI211_X1 port map( C1 => n5037, C2 => n5200, A => n5036, B => n5035
                           , ZN => n5038);
   U5639 : NAND2_X1 port map( A1 => n5038, A2 => n5313, ZN => n5050);
   U5640 : AOI22_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx6x, 
                           B1 => n5140, B2 => fromRegsPortxREG_FILE_07xx6x, ZN 
                           => n5043);
   U5641 : AOI22_X1 port map( A1 => n5203, A2 => fromRegsPortxREG_FILE_09xx6x, 
                           B1 => n5073, B2 => fromRegsPortxREG_FILE_04xx6x, ZN 
                           => n5042);
   U5642 : AOI22_X1 port map( A1 => n5039, A2 => fromRegsPortxREG_FILE_08xx6x, 
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx6x, ZN 
                           => n5041);
   U5643 : NAND2_X1 port map( A1 => n5142, A2 => fromRegsPortxREG_FILE_03xx6x, 
                           ZN => n5040);
   U5644 : NAND4_X1 port map( A1 => n5043, A2 => n5042, A3 => n5041, A4 => 
                           n5040, ZN => n5048);
   U5645 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx6x, 
                           ZN => n5045);
   U5646 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx6x, A2 => n5327, 
                           ZN => n5044);
   U5647 : NAND2_X1 port map( A1 => n5045, A2 => n5044, ZN => n5046);
   U5648 : AOI21_X1 port map( B1 => n5048, B2 => n5047, A => n5046, ZN => n5049
                           );
   U5649 : NAND2_X1 port map( A1 => n5050, A2 => n5049, ZN => n6353);
   U5650 : INV_X1 port map( A => n6353, ZN => n7458);
   U5651 : INV_X1 port map( A => add_x_26xBx6x, ZN => n6359);
   U5652 : OAI22_X1 port map( A1 => n5677, A2 => n7458, B1 => n5675, B2 => 
                           n6359, ZN => n5051);
   U5653 : XOR2_X1 port map( A => n5252, B => n5051, Z => 
                           DP_OP_719J1_125_1055xn62);
   U5654 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(25), A2 => n5052,
                           ZN => add_x_26xBx5x);
   U5655 : AOI22_X1 port map( A1 => n5086, A2 => fromRegsPortxREG_FILE_30xx5x, 
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_27xx5x, ZN 
                           => n5058);
   U5656 : AOI22_X1 port map( A1 => n5182, A2 => fromRegsPortxREG_FILE_25xx5x, 
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_24xx5x, ZN 
                           => n5057);
   U5657 : AOI22_X1 port map( A1 => n5053, A2 => fromRegsPortxREG_FILE_29xx5x, 
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx5x, ZN 
                           => n5056);
   U5658 : AOI22_X1 port map( A1 => n5054, A2 => fromRegsPortxREG_FILE_31xx5x, 
                           B1 => n5085, B2 => fromRegsPortxREG_FILE_28xx5x, ZN 
                           => n5055);
   U5659 : NAND4_X1 port map( A1 => n5058, A2 => n5057, A3 => n5056, A4 => 
                           n5055, ZN => n5064);
   U5660 : AOI22_X1 port map( A1 => n5092, A2 => fromRegsPortxREG_FILE_20xx5x, 
                           B1 => n5187, B2 => fromRegsPortxREG_FILE_19xx5x, ZN 
                           => n5062);
   U5661 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_21xx5x, 
                           B1 => n5125, B2 => fromRegsPortxREG_FILE_17xx5x, ZN 
                           => n5061);
   U5662 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx5x, 
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx5x, ZN 
                           => n5060);
   U5663 : NAND2_X1 port map( A1 => n5287, A2 => fromRegsPortxREG_FILE_22xx5x, 
                           ZN => n5059);
   U5664 : NAND4_X1 port map( A1 => n5062, A2 => n5061, A3 => n5060, A4 => 
                           n5059, ZN => n5063);
   U5665 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5064
                           , A => n5063, ZN => n5071);
   U5666 : AOI22_X1 port map( A1 => n5065, A2 => fromRegsPortxREG_FILE_16xx5x, 
                           B1 => n5100, B2 => fromRegsPortxREG_FILE_15xx5x, ZN 
                           => n5070);
   U5667 : AOI22_X1 port map( A1 => n5102, A2 => fromRegsPortxREG_FILE_14xx5x, 
                           B1 => n5101, B2 => fromRegsPortxREG_FILE_11xx5x, ZN 
                           => n5067);
   U5668 : AOI22_X1 port map( A1 => n5301, A2 => fromRegsPortxREG_FILE_12xx5x, 
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx5x, ZN 
                           => n5066);
   U5669 : NAND2_X1 port map( A1 => n5067, A2 => n5066, ZN => n5068);
   U5670 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx5x, B2 => n5165, 
                           A => n5068, ZN => n5069);
   U5671 : OAI211_X1 port map( C1 => n5071, C2 => n5200, A => n5070, B => n5069
                           , ZN => n5072);
   U5672 : NAND2_X1 port map( A1 => n5072, A2 => n5313, ZN => n5083);
   U5673 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx5x, 
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx5x, ZN 
                           => n5077);
   U5674 : AOI22_X1 port map( A1 => n5141, A2 => fromRegsPortxREG_FILE_06xx5x, 
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx5x, ZN 
                           => n5076);
   U5675 : AOI22_X1 port map( A1 => n5073, A2 => fromRegsPortxREG_FILE_04xx5x, 
                           B1 => n5140, B2 => fromRegsPortxREG_FILE_07xx5x, ZN 
                           => n5075);
   U5676 : NAND2_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx5x, 
                           ZN => n5074);
   U5677 : NAND4_X1 port map( A1 => n5077, A2 => n5076, A3 => n5075, A4 => 
                           n5074, ZN => n5081);
   U5678 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx5x, 
                           ZN => n5079);
   U5679 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx5x, A2 => n5327, 
                           ZN => n5078);
   U5680 : NAND2_X1 port map( A1 => n5079, A2 => n5078, ZN => n5080);
   U5681 : AOI21_X1 port map( B1 => n5081, B2 => n5331, A => n5080, ZN => n5082
                           );
   U5682 : NAND2_X1 port map( A1 => n5083, A2 => n5082, ZN => n5399);
   U5683 : INV_X1 port map( A => n5399, ZN => n7457);
   U5684 : INV_X1 port map( A => add_x_26xBx5x, ZN => n6307);
   U5685 : OAI22_X1 port map( A1 => n7457, A2 => n7360, B1 => n5675, B2 => 
                           n6307, ZN => n5084);
   U5686 : XOR2_X1 port map( A => n5252, B => n5084, Z => 
                           DP_OP_719J1_125_1055xn63);
   U5687 : AOI22_X1 port map( A1 => n5086, A2 => fromRegsPortxREG_FILE_30xx4x, 
                           B1 => n5085, B2 => fromRegsPortxREG_FILE_28xx4x, ZN 
                           => n5091);
   U5688 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx4x, 
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_24xx4x, ZN 
                           => n5090);
   U5689 : AOI22_X1 port map( A1 => n5182, A2 => fromRegsPortxREG_FILE_25xx4x, 
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_27xx4x, ZN 
                           => n5089);
   U5690 : AOI22_X1 port map( A1 => n5087, A2 => fromRegsPortxREG_FILE_26xx4x, 
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx4x, ZN 
                           => n5088);
   U5691 : NAND4_X1 port map( A1 => n5091, A2 => n5090, A3 => n5089, A4 => 
                           n5088, ZN => n5099);
   U5692 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx4x, 
                           B1 => n5125, B2 => fromRegsPortxREG_FILE_17xx4x, ZN 
                           => n5097);
   U5693 : AOI22_X1 port map( A1 => n5092, A2 => fromRegsPortxREG_FILE_20xx4x, 
                           B1 => n5289, B2 => fromRegsPortxREG_FILE_23xx4x, ZN 
                           => n5096);
   U5694 : AOI22_X1 port map( A1 => n5093, A2 => fromRegsPortxREG_FILE_18xx4x, 
                           B1 => n5187, B2 => fromRegsPortxREG_FILE_19xx4x, ZN 
                           => n5095);
   U5695 : NAND2_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_21xx4x, 
                           ZN => n5094);
   U5696 : NAND4_X1 port map( A1 => n5097, A2 => n5096, A3 => n5095, A4 => 
                           n5094, ZN => n5098);
   U5697 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5099
                           , A => n5098, ZN => n5108);
   U5698 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_13xx4x, 
                           B1 => n5100, B2 => fromRegsPortxREG_FILE_15xx4x, ZN 
                           => n5107);
   U5699 : AOI22_X1 port map( A1 => n5102, A2 => fromRegsPortxREG_FILE_14xx4x, 
                           B1 => n5101, B2 => fromRegsPortxREG_FILE_11xx4x, ZN 
                           => n5104);
   U5700 : AOI22_X1 port map( A1 => n5234, A2 => fromRegsPortxREG_FILE_12xx4x, 
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx4x, ZN 
                           => n5103);
   U5701 : NAND2_X1 port map( A1 => n5104, A2 => n5103, ZN => n5105);
   U5702 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx4x, B2 => n5300, 
                           A => n5105, ZN => n5106);
   U5703 : OAI211_X1 port map( C1 => n5108, C2 => n5200, A => n5107, B => n5106
                           , ZN => n5117);
   U5704 : AOI22_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx4x, 
                           B1 => n5140, B2 => fromRegsPortxREG_FILE_07xx4x, ZN 
                           => n5112);
   U5705 : AOI22_X1 port map( A1 => n5203, A2 => fromRegsPortxREG_FILE_09xx4x, 
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx4x, ZN 
                           => n5111);
   U5706 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx4x, 
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx4x, ZN 
                           => n5110);
   U5707 : NAND2_X1 port map( A1 => n5142, A2 => fromRegsPortxREG_FILE_03xx4x, 
                           ZN => n5109);
   U5708 : NAND4_X1 port map( A1 => n5112, A2 => n5111, A3 => n5110, A4 => 
                           n5109, ZN => n5113);
   U5709 : NAND2_X1 port map( A1 => n5113, A2 => n5331, ZN => n5115);
   U5710 : AOI22_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx4x, 
                           B1 => n5327, B2 => fromRegsPortxREG_FILE_01xx4x, ZN 
                           => n5114);
   U5711 : NAND2_X1 port map( A1 => n5115, A2 => n5114, ZN => n5116);
   U5712 : INV_X1 port map( A => ashr_25xSHx4x, ZN => n7327);
   U5713 : OAI22_X1 port map( A1 => n7081, A2 => n5674, B1 => n5675, B2 => 
                           n7327, ZN => n5118);
   U5714 : XOR2_X1 port map( A => n7546, B => n5118, Z => 
                           DP_OP_719J1_125_1055xn64);
   U5715 : AOI22_X1 port map( A1 => n5120, A2 => fromRegsPortxREG_FILE_24xx3x, 
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_27xx3x, ZN 
                           => n5124);
   U5716 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx3x, 
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx3x, ZN 
                           => n5123);
   U5717 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx3x, 
                           B1 => n5276, B2 => fromRegsPortxREG_FILE_25xx3x, ZN 
                           => n5122);
   U5718 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_26xx3x, 
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx3x, ZN 
                           => n5121);
   U5719 : NAND4_X1 port map( A1 => n5124, A2 => n5123, A3 => n5122, A4 => 
                           n5121, ZN => n5132);
   U5720 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx3x, 
                           B1 => n5187, B2 => fromRegsPortxREG_FILE_19xx3x, ZN 
                           => n5130);
   U5721 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_21xx3x, 
                           B1 => n5125, B2 => fromRegsPortxREG_FILE_17xx3x, ZN 
                           => n5129);
   U5722 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx3x, 
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx3x, ZN 
                           => n5128);
   U5723 : NAND2_X1 port map( A1 => n5126, A2 => fromRegsPortxREG_FILE_23xx3x, 
                           ZN => n5127);
   U5724 : NAND4_X1 port map( A1 => n5130, A2 => n5129, A3 => n5128, A4 => 
                           n5127, ZN => n5131);
   U5725 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5132
                           , A => n5131, ZN => n5138);
   U5726 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_13xx3x, 
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx3x, ZN 
                           => n5137);
   U5727 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_10xx3x, 
                           B1 => n5303, B2 => fromRegsPortxREG_FILE_11xx3x, ZN 
                           => n5134);
   U5728 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx3x, 
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx3x, ZN 
                           => n5133);
   U5729 : NAND2_X1 port map( A1 => n5134, A2 => n5133, ZN => n5135);
   U5730 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx3x, B2 => n5234, 
                           A => n5135, ZN => n5136);
   U5731 : OAI211_X1 port map( C1 => n5138, C2 => n5200, A => n5137, B => n5136
                           , ZN => n5139);
   U5732 : NAND2_X1 port map( A1 => n5139, A2 => n5313, ZN => n5152);
   U5733 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_08xx3x, 
                           B1 => n5140, B2 => fromRegsPortxREG_FILE_07xx3x, ZN 
                           => n5146);
   U5734 : AOI22_X1 port map( A1 => n5203, A2 => fromRegsPortxREG_FILE_09xx3x, 
                           B1 => n5141, B2 => fromRegsPortxREG_FILE_06xx3x, ZN 
                           => n5145);
   U5735 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx3x, 
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx3x, ZN 
                           => n5144);
   U5736 : NAND2_X1 port map( A1 => n5142, A2 => fromRegsPortxREG_FILE_03xx3x, 
                           ZN => n5143);
   U5737 : NAND4_X1 port map( A1 => n5146, A2 => n5145, A3 => n5144, A4 => 
                           n5143, ZN => n5150);
   U5738 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx3x, 
                           ZN => n5148);
   U5739 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx3x, A2 => n5327, 
                           ZN => n5147);
   U5740 : NAND2_X1 port map( A1 => n5148, A2 => n5147, ZN => n5149);
   U5741 : AOI21_X1 port map( B1 => n5150, B2 => n5331, A => n5149, ZN => n5151
                           );
   U5742 : NAND2_X2 port map( A1 => n5152, A2 => n5151, ZN => n7203);
   U5743 : INV_X2 port map( A => n7203, ZN => n7372);
   U5744 : OAI22_X1 port map( A1 => n7372, A2 => n5677, B1 => n5675, B2 => 
                           intadd_4xBx2x, ZN => n5153);
   U5745 : XOR2_X1 port map( A => n5252, B => n5153, Z => 
                           DP_OP_719J1_125_1055xn65);
   U5746 : AOI22_X1 port map( A1 => n5182, A2 => fromRegsPortxREG_FILE_25xx2x, 
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx2x, ZN 
                           => n5157);
   U5747 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx2x, 
                           B1 => n5278, B2 => fromRegsPortxREG_FILE_29xx2x, ZN 
                           => n5156);
   U5748 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_24xx2x, 
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx2x, ZN 
                           => n5155);
   U5749 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_27xx2x, 
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx2x, ZN 
                           => n5154);
   U5750 : NAND4_X1 port map( A1 => n5157, A2 => n5156, A3 => n5155, A4 => 
                           n5154, ZN => n5164);
   U5751 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_21xx2x, 
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx2x, ZN 
                           => n5162);
   U5752 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx2x, 
                           B1 => n5224, B2 => fromRegsPortxREG_FILE_22xx2x, ZN 
                           => n5161);
   U5753 : AOI22_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_18xx2x, 
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_19xx2x, ZN 
                           => n5160);
   U5754 : NAND2_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx2x, 
                           ZN => n5159);
   U5755 : NAND4_X1 port map( A1 => n5162, A2 => n5161, A3 => n5160, A4 => 
                           n5159, ZN => n5163);
   U5756 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5164
                           , A => n5163, ZN => n5171);
   U5757 : AOI22_X1 port map( A1 => n5301, A2 => fromRegsPortxREG_FILE_12xx2x, 
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx2x, ZN 
                           => n5170);
   U5758 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_10xx2x, 
                           B1 => n5302, B2 => fromRegsPortxREG_FILE_14xx2x, ZN 
                           => n5167);
   U5759 : AOI22_X1 port map( A1 => n5309, A2 => fromRegsPortxREG_FILE_16xx2x, 
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx2x, ZN 
                           => n5166);
   U5760 : NAND2_X1 port map( A1 => n5167, A2 => n5166, ZN => n5168);
   U5761 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_11xx2x, B2 => n5303, 
                           A => n5168, ZN => n5169);
   U5762 : OAI211_X1 port map( C1 => n5171, C2 => n5200, A => n5170, B => n5169
                           , ZN => n5180);
   U5763 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx2x, 
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx2x, ZN 
                           => n5175);
   U5764 : AOI22_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx2x, 
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx2x, ZN 
                           => n5174);
   U5765 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx2x, 
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx2x, ZN 
                           => n5173);
   U5766 : NAND2_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx2x, 
                           ZN => n5172);
   U5767 : NAND4_X1 port map( A1 => n5175, A2 => n5174, A3 => n5173, A4 => 
                           n5172, ZN => n5176);
   U5768 : NAND2_X1 port map( A1 => n5176, A2 => n5331, ZN => n5178);
   U5769 : AOI22_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx2x, 
                           B1 => n5327, B2 => fromRegsPortxREG_FILE_01xx2x, ZN 
                           => n5177);
   U5770 : NAND2_X1 port map( A1 => n5178, A2 => n5177, ZN => n5179);
   U5771 : AOI21_X1 port map( B1 => n5180, B2 => n5313, A => n5179, ZN => n6600
                           );
   U5772 : CLKBUF_X1 port map( A => n6600, Z => n7038);
   U5773 : OAI22_X1 port map( A1 => intadd_4xBx1x, A2 => n5675, B1 => n5674, B2
                           => n7038, ZN => n5181);
   U5774 : XOR2_X1 port map( A => n7546, B => n5181, Z => 
                           DP_OP_719J1_125_1055xn66);
   U5775 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx1x, 
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_27xx1x, ZN 
                           => n5186);
   U5776 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_26xx1x, 
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx1x, ZN 
                           => n5185);
   U5777 : AOI22_X1 port map( A1 => n5182, A2 => fromRegsPortxREG_FILE_25xx1x, 
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_24xx1x, ZN 
                           => n5184);
   U5778 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx1x, 
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx1x, ZN 
                           => n5183);
   U5779 : NAND4_X1 port map( A1 => n5186, A2 => n5185, A3 => n5184, A4 => 
                           n5183, ZN => n5193);
   U5780 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx1x, 
                           B1 => n5187, B2 => fromRegsPortxREG_FILE_19xx1x, ZN 
                           => n5191);
   U5781 : AOI22_X1 port map( A1 => n5288, A2 => fromRegsPortxREG_FILE_21xx1x, 
                           B1 => n5287, B2 => fromRegsPortxREG_FILE_22xx1x, ZN 
                           => n5190);
   U5782 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx1x, 
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx1x, ZN 
                           => n5189);
   U5783 : NAND2_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_18xx1x, 
                           ZN => n5188);
   U5784 : NAND4_X1 port map( A1 => n5191, A2 => n5190, A3 => n5189, A4 => 
                           n5188, ZN => n5192);
   U5785 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5193
                           , A => n5192, ZN => n5201);
   U5786 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_11xx1x, 
                           B1 => n5194, B2 => fromRegsPortxREG_FILE_13xx1x, ZN 
                           => n5199);
   U5787 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx1x, 
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx1x, ZN 
                           => n5196);
   U5788 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx1x, 
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx1x, ZN 
                           => n5195);
   U5789 : NAND2_X1 port map( A1 => n5196, A2 => n5195, ZN => n5197);
   U5790 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx1x, B2 => n5234, 
                           A => n5197, ZN => n5198);
   U5791 : OAI211_X1 port map( C1 => n5201, C2 => n5200, A => n5199, B => n5198
                           , ZN => n5202);
   U5792 : NAND2_X1 port map( A1 => n5202, A2 => n5313, ZN => n5213);
   U5793 : AOI22_X1 port map( A1 => n5203, A2 => fromRegsPortxREG_FILE_09xx1x, 
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx1x, ZN 
                           => n5207);
   U5794 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx1x, 
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx1x, ZN 
                           => n5206);
   U5795 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx1x, 
                           B1 => n5316, B2 => fromRegsPortxREG_FILE_06xx1x, ZN 
                           => n5205);
   U5796 : NAND2_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_05xx1x, 
                           ZN => n5204);
   U5797 : NAND4_X1 port map( A1 => n5207, A2 => n5206, A3 => n5205, A4 => 
                           n5204, ZN => n5211);
   U5798 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx1x, 
                           ZN => n5209);
   U5799 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx1x, A2 => n5244, 
                           ZN => n5208);
   U5800 : NAND2_X1 port map( A1 => n5209, A2 => n5208, ZN => n5210);
   U5801 : AOI21_X1 port map( B1 => n5211, B2 => n5331, A => n5210, ZN => n5212
                           );
   U5802 : NAND2_X1 port map( A1 => n5213, A2 => n5212, ZN => n7082);
   U5803 : CLKBUF_X1 port map( A => n7082, Z => n7399);
   U5804 : INV_X1 port map( A => n7399, ZN => n6144);
   U5805 : OAI22_X1 port map( A1 => intadd_4xBx0x, A2 => n5675, B1 => n5674, B2
                           => n6144, ZN => n5214);
   U5806 : XOR2_X1 port map( A => n7546, B => n5214, Z => 
                           DP_OP_719J1_125_1055xn67);
   U5807 : NAND2_X1 port map( A1 => n7456, A2 => fromMemoryPortxLOADEDDATAx(7),
                           ZN => n5219);
   U5808 : AND2_X1 port map( A1 => n7448, A2 => n5215, ZN => n5216);
   U5809 : NAND2_X1 port map( A1 => n5712, A2 => n5216, ZN => n5217);
   U5810 : NAND2_X1 port map( A1 => n5217, A2 => fromMemoryPortxLOADEDDATAx(20)
                           , ZN => n5218);
   U5811 : NAND2_X2 port map( A1 => n5219, A2 => n5218, ZN => n7408);
   U5812 : INV_X1 port map( A => n7408, ZN => n7329);
   U5813 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_27xx0x, 
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_28xx0x, ZN 
                           => n5223);
   U5814 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_29xx0x, 
                           B1 => n5277, B2 => fromRegsPortxREG_FILE_26xx0x, ZN 
                           => n5222);
   U5815 : AOI22_X1 port map( A1 => n5275, A2 => fromRegsPortxREG_FILE_30xx0x, 
                           B1 => n5276, B2 => fromRegsPortxREG_FILE_25xx0x, ZN 
                           => n5221);
   U5816 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_24xx0x, 
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_31xx0x, ZN 
                           => n5220);
   U5817 : NAND4_X1 port map( A1 => n5223, A2 => n5222, A3 => n5221, A4 => 
                           n5220, ZN => n5230);
   U5818 : AOI22_X1 port map( A1 => n5224, A2 => fromRegsPortxREG_FILE_22xx0x, 
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_18xx0x, ZN 
                           => n5228);
   U5819 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_23xx0x, 
                           B1 => n5288, B2 => fromRegsPortxREG_FILE_21xx0x, ZN 
                           => n5227);
   U5820 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_20xx0x, 
                           B1 => n5292, B2 => fromRegsPortxREG_FILE_17xx0x, ZN 
                           => n5226);
   U5821 : NAND2_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_19xx0x, 
                           ZN => n5225);
   U5822 : NAND4_X1 port map( A1 => n5228, A2 => n5227, A3 => n5226, A4 => 
                           n5225, ZN => n5229);
   U5823 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5230
                           , A => n5229, ZN => n5237);
   U5824 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_13xx0x, 
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_15xx0x, ZN 
                           => n5236);
   U5825 : AOI22_X1 port map( A1 => n5300, A2 => fromRegsPortxREG_FILE_10xx0x, 
                           B1 => n5303, B2 => fromRegsPortxREG_FILE_11xx0x, ZN 
                           => n5232);
   U5826 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_14xx0x, 
                           B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx0x, ZN 
                           => n5231);
   U5827 : NAND2_X1 port map( A1 => n5232, A2 => n5231, ZN => n5233);
   U5828 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx0x, B2 => n5234, 
                           A => n5233, ZN => n5235);
   U5829 : OAI211_X1 port map( C1 => n5237, C2 => n5758, A => n5236, B => n5235
                           , ZN => n5239);
   U5830 : NAND2_X1 port map( A1 => n5239, A2 => n5238, ZN => n5250);
   U5831 : AOI22_X1 port map( A1 => n5315, A2 => fromRegsPortxREG_FILE_03xx0x, 
                           B1 => n5321, B2 => fromRegsPortxREG_FILE_08xx0x, ZN 
                           => n5243);
   U5832 : AOI22_X1 port map( A1 => n5316, A2 => fromRegsPortxREG_FILE_06xx0x, 
                           B1 => n5320, B2 => fromRegsPortxREG_FILE_05xx0x, ZN 
                           => n5242);
   U5833 : AOI22_X1 port map( A1 => n5317, A2 => fromRegsPortxREG_FILE_04xx0x, 
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_07xx0x, ZN 
                           => n5241);
   U5834 : NAND2_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_09xx0x, 
                           ZN => n5240);
   U5835 : NAND4_X1 port map( A1 => n5243, A2 => n5242, A3 => n5241, A4 => 
                           n5240, ZN => n5248);
   U5836 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx0x, 
                           ZN => n5246);
   U5837 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx0x, A2 => n5244, 
                           ZN => n5245);
   U5838 : NAND2_X1 port map( A1 => n5246, A2 => n5245, ZN => n5247);
   U5839 : AOI21_X1 port map( B1 => n5248, B2 => n5331, A => n5247, ZN => n5249
                           );
   U5840 : NAND2_X1 port map( A1 => n5250, A2 => n5249, ZN => n7395);
   U5841 : CLKBUF_X1 port map( A => n7395, Z => n7161);
   U5842 : INV_X1 port map( A => n7161, ZN => n7396);
   U5843 : OAI22_X1 port map( A1 => n5673, A2 => n7329, B1 => n5677, B2 => 
                           n7396, ZN => n5251);
   U5844 : XOR2_X1 port map( A => n5252, B => n5251, Z => 
                           DP_OP_719J1_125_1055xn68);
   U5845 : XOR2_X1 port map( A => n7547, B => n7317, Z => 
                           DP_OP_679J1_122_3096xn38);
   U5846 : XOR2_X1 port map( A => n7547, B => n7247, Z => 
                           DP_OP_679J1_122_3096xn39);
   U5847 : XOR2_X1 port map( A => n7547, B => n7237, Z => 
                           DP_OP_679J1_122_3096xn40);
   U5848 : XOR2_X1 port map( A => n7547, B => n7179, Z => 
                           DP_OP_679J1_122_3096xn41);
   U5849 : XOR2_X1 port map( A => n7547, B => n7114, Z => 
                           DP_OP_679J1_122_3096xn42);
   U5850 : XOR2_X1 port map( A => n7547, B => n7093, Z => 
                           DP_OP_679J1_122_3096xn43);
   U5851 : XOR2_X1 port map( A => n7547, B => n5744, Z => 
                           DP_OP_679J1_122_3096xn44);
   U5852 : XOR2_X1 port map( A => n5679, B => n7028, Z => 
                           DP_OP_679J1_122_3096xn45);
   U5853 : XOR2_X1 port map( A => n5679, B => n6986, Z => 
                           DP_OP_679J1_122_3096xn46);
   U5854 : XOR2_X1 port map( A => n5679, B => n5717, Z => 
                           DP_OP_679J1_122_3096xn47);
   U5855 : XOR2_X1 port map( A => n5679, B => n6962, Z => 
                           DP_OP_679J1_122_3096xn48);
   U5856 : XOR2_X1 port map( A => n5679, B => n6918, Z => 
                           DP_OP_679J1_122_3096xn49);
   U5857 : XOR2_X1 port map( A => n5679, B => n6891, Z => 
                           DP_OP_679J1_122_3096xn50);
   U5858 : XOR2_X1 port map( A => n7547, B => n6835, Z => 
                           DP_OP_679J1_122_3096xn51);
   U5859 : XOR2_X1 port map( A => n7547, B => n6805, Z => 
                           DP_OP_679J1_122_3096xn52);
   U5860 : XOR2_X1 port map( A => n7547, B => n6774, Z => 
                           DP_OP_679J1_122_3096xn53);
   U5861 : XOR2_X1 port map( A => n7547, B => n6726, Z => 
                           DP_OP_679J1_122_3096xn54);
   U5862 : XOR2_X1 port map( A => n7547, B => n6702, Z => 
                           DP_OP_679J1_122_3096xn55);
   U5863 : XOR2_X1 port map( A => n7547, B => n6658, Z => 
                           DP_OP_679J1_122_3096xn56);
   U5864 : XOR2_X1 port map( A => n7547, B => n6616, Z => 
                           DP_OP_679J1_122_3096xn57);
   U5865 : XOR2_X1 port map( A => n7547, B => n6555, Z => 
                           DP_OP_679J1_122_3096xn58);
   U5866 : XOR2_X1 port map( A => n7547, B => n6504, Z => 
                           DP_OP_679J1_122_3096xn59);
   U5867 : XOR2_X1 port map( A => n7547, B => n6445, Z => 
                           DP_OP_679J1_122_3096xn60);
   U5868 : XOR2_X1 port map( A => n7547, B => n6406, Z => 
                           DP_OP_679J1_122_3096xn61);
   U5869 : XOR2_X1 port map( A => n7547, B => n6353, Z => 
                           DP_OP_679J1_122_3096xn62);
   U5870 : XOR2_X1 port map( A => n7547, B => n5399, Z => 
                           DP_OP_679J1_122_3096xn63);
   U5871 : INV_X1 port map( A => n7081, ZN => n7345);
   U5872 : XOR2_X1 port map( A => n7547, B => n7345, Z => 
                           DP_OP_679J1_122_3096xn64);
   U5873 : XOR2_X1 port map( A => n7547, B => n7203, Z => 
                           DP_OP_679J1_122_3096xn65);
   U5874 : CLKBUF_X1 port map( A => n6600, Z => n7305);
   U5875 : INV_X1 port map( A => n7305, ZN => n7036);
   U5876 : XOR2_X1 port map( A => n7547, B => n7036, Z => 
                           DP_OP_679J1_122_3096xn66);
   U5877 : CLKBUF_X1 port map( A => n7082, Z => n7263);
   U5878 : XOR2_X1 port map( A => n7547, B => n7263, Z => 
                           DP_OP_679J1_122_3096xn67);
   U5879 : CLKBUF_X1 port map( A => n7395, Z => n7296);
   U5880 : XOR2_X1 port map( A => n7547, B => n7296, Z => 
                           DP_OP_679J1_122_3096xn68);
   U5881 : INV_X1 port map( A => ashr_25xAx1x, ZN => intadd_4xAx0x);
   U5882 : INV_X1 port map( A => ashr_25xAx30x, ZN => intadd_3xAx2x);
   U5883 : INV_X1 port map( A => ashr_25xAx29x, ZN => intadd_3xAx1x);
   U5884 : INV_X1 port map( A => ashr_25xAx28x, ZN => intadd_3xAx0x);
   U5885 : INV_X1 port map( A => ashr_25xAx14x, ZN => intadd_2xAx3x);
   U5886 : INV_X1 port map( A => ashr_25xAx13x, ZN => intadd_2xAx2x);
   U5887 : INV_X1 port map( A => ashr_25xAx11x, ZN => intadd_2xAx0x);
   U5888 : INV_X1 port map( A => ashr_25xAx24x, ZN => intadd_1xAx7x);
   U5889 : INV_X1 port map( A => ashr_25xAx23x, ZN => intadd_1xAx6x);
   U5890 : INV_X1 port map( A => ashr_25xAx22x, ZN => intadd_1xAx5x);
   U5891 : INV_X1 port map( A => ashr_25xAx21x, ZN => intadd_1xAx4x);
   U5892 : INV_X1 port map( A => ashr_25xAx20x, ZN => intadd_1xAx3x);
   U5893 : INV_X1 port map( A => ashr_25xAx19x, ZN => intadd_1xAx2x);
   U5894 : INV_X1 port map( A => ashr_25xAx18x, ZN => intadd_1xAx1x);
   U5895 : INV_X1 port map( A => ashr_25xAx17x, ZN => intadd_1xAx0x);
   U5896 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_28xx26x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_27xx26x, ZN
                           => n5257);
   U5897 : AOI22_X1 port map( A1 => n5359, A2 => fromRegsPortxREG_FILE_06xx26x,
                           B1 => n5348, B2 => fromRegsPortxREG_FILE_29xx26x, ZN
                           => n5256);
   U5898 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx26x,
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_26xx26x, ZN
                           => n5255);
   U5899 : NAND2_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_04xx26x,
                           ZN => n5254);
   U5900 : AND4_X1 port map( A1 => n5257, A2 => n5256, A3 => n5255, A4 => n5254
                           , ZN => n5274);
   U5901 : AOI22_X1 port map( A1 => n5373, A2 => fromRegsPortxREG_FILE_24xx26x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_21xx26x, ZN
                           => n5262);
   U5902 : AOI22_X1 port map( A1 => n5337, A2 => fromRegsPortxREG_FILE_09xx26x,
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx26x, ZN
                           => n5261);
   U5903 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx26x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_16xx26x, ZN
                           => n5260);
   U5904 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx26x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_12xx26x, ZN
                           => n5259);
   U5905 : AND4_X1 port map( A1 => n5262, A2 => n5261, A3 => n5260, A4 => n5259
                           , ZN => n5273);
   U5906 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_15xx26x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_10xx26x, ZN
                           => n5266);
   U5907 : AOI22_X1 port map( A1 => n5364, A2 => fromRegsPortxREG_FILE_19xx26x,
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx26x, ZN
                           => n5265);
   U5908 : AOI22_X1 port map( A1 => n5335, A2 => fromRegsPortxREG_FILE_23xx26x,
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_11xx26x, ZN
                           => n5264);
   U5909 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_20xx26x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx26x, ZN
                           => n5263);
   U5910 : AND4_X1 port map( A1 => n5266, A2 => n5265, A3 => n5264, A4 => n5263
                           , ZN => n5272);
   U5911 : AOI22_X1 port map( A1 => n5347, A2 => fromRegsPortxREG_FILE_17xx26x,
                           B1 => n5372, B2 => fromRegsPortxREG_FILE_02xx26x, ZN
                           => n5270);
   U5912 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_31xx26x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_03xx26x, ZN
                           => n5269);
   U5913 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx26x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx26x, ZN
                           => n5268);
   U5914 : AOI22_X1 port map( A1 => n5371, A2 => fromRegsPortxREG_FILE_05xx26x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_07xx26x, ZN
                           => n5267);
   U5915 : AND4_X1 port map( A1 => n5270, A2 => n5269, A3 => n5268, A4 => n5267
                           , ZN => n5271);
   U5916 : NAND4_X1 port map( A1 => n5274, A2 => n5273, A3 => n5272, A4 => 
                           n5271, ZN => ashr_25xAx26x);
   U5917 : NAND2_X1 port map( A1 => n7534, A2 => n7505, ZN => n5973);
   U5918 : INV_X1 port map( A => n5973, ZN => n5848);
   U5919 : INV_X1 port map( A => n5848, ZN => n5957);
   U5920 : NAND2_X1 port map( A1 => n5760, A2 => n7531, ZN => n5761);
   U5921 : NOR4_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(2), A2 => n5957, 
                           A3 => n6388, A4 => n5761, ZN => n5440);
   U5922 : AND2_X1 port map( A1 => n5440, A2 => n5762, ZN => n5658);
   U5923 : INV_X1 port map( A => n5658, ZN => n5624);
   U5924 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_25xx31x, A2 => n5276,
                           B1 => fromRegsPortxREG_FILE_30xx31x, B2 => n5275, ZN
                           => n5286);
   U5925 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_29xx31x, A2 => n5278,
                           B1 => fromRegsPortxREG_FILE_26xx31x, B2 => n5277, ZN
                           => n5285);
   U5926 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_24xx31x, A2 => n5280,
                           B1 => fromRegsPortxREG_FILE_27xx31x, B2 => n5279, ZN
                           => n5284);
   U5927 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_31xx31x, A2 => n5282,
                           B1 => fromRegsPortxREG_FILE_28xx31x, B2 => n5281, ZN
                           => n5283);
   U5928 : NAND4_X1 port map( A1 => n5286, A2 => n5285, A3 => n5284, A4 => 
                           n5283, ZN => n5299);
   U5929 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_21xx31x, A2 => n5288,
                           B1 => fromRegsPortxREG_FILE_22xx31x, B2 => n5287, ZN
                           => n5297);
   U5930 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_20xx31x, A2 => n5290,
                           B1 => fromRegsPortxREG_FILE_23xx31x, B2 => n5289, ZN
                           => n5296);
   U5931 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_17xx31x, A2 => n5292,
                           B1 => fromRegsPortxREG_FILE_19xx31x, B2 => n5291, ZN
                           => n5295);
   U5932 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_18xx31x, A2 => n5293,
                           ZN => n5294);
   U5933 : NAND4_X1 port map( A1 => n5297, A2 => n5296, A3 => n5295, A4 => 
                           n5294, ZN => n5298);
   U5934 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5299
                           , A => n5298, ZN => n5312);
   U5935 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_12xx31x, A2 => n5301,
                           B1 => fromRegsPortxREG_FILE_10xx31x, B2 => n5300, ZN
                           => n5311);
   U5936 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_11xx31x, A2 => n5303,
                           B1 => fromRegsPortxREG_FILE_14xx31x, B2 => n5302, ZN
                           => n5307);
   U5937 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_15xx31x, A2 => n5305,
                           B1 => fromRegsPortxREG_FILE_13xx31x, B2 => n5304, ZN
                           => n5306);
   U5938 : NAND2_X1 port map( A1 => n5307, A2 => n5306, ZN => n5308);
   U5939 : AOI21_X1 port map( B1 => n5309, B2 => fromRegsPortxREG_FILE_16xx31x,
                           A => n5308, ZN => n5310);
   U5940 : OAI211_X1 port map( C1 => n5312, C2 => n5758, A => n5311, B => n5310
                           , ZN => n5314);
   U5941 : NAND2_X1 port map( A1 => n5314, A2 => n5313, ZN => n5334);
   U5942 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_06xx31x, A2 => n5316,
                           B1 => fromRegsPortxREG_FILE_03xx31x, B2 => n5315, ZN
                           => n5325);
   U5943 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_09xx31x, A2 => n5318,
                           B1 => fromRegsPortxREG_FILE_04xx31x, B2 => n5317, ZN
                           => n5324);
   U5944 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_05xx31x, A2 => n5320,
                           B1 => fromRegsPortxREG_FILE_07xx31x, B2 => n5319, ZN
                           => n5323);
   U5945 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_08xx31x, A2 => n5321,
                           ZN => n5322);
   U5946 : NAND4_X1 port map( A1 => n5325, A2 => n5324, A3 => n5323, A4 => 
                           n5322, ZN => n5332);
   U5947 : NAND2_X1 port map( A1 => n5326, A2 => fromRegsPortxREG_FILE_02xx31x,
                           ZN => n5329);
   U5948 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx31x, A2 => n5327,
                           ZN => n5328);
   U5949 : NAND2_X1 port map( A1 => n5329, A2 => n5328, ZN => n5330);
   U5950 : AOI21_X1 port map( B1 => n5332, B2 => n5331, A => n5330, ZN => n5333
                           );
   U5951 : NAND2_X1 port map( A1 => n5334, A2 => n5333, ZN => n7384);
   U5952 : XOR2_X1 port map( A => n7547, B => n7384, Z => n5386);
   U5953 : AOI22_X1 port map( A1 => n5336, A2 => fromRegsPortxREG_FILE_30xx31x,
                           B1 => n5335, B2 => fromRegsPortxREG_FILE_23xx31x, ZN
                           => n5346);
   U5954 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_11xx31x,
                           B1 => n5337, B2 => fromRegsPortxREG_FILE_09xx31x, ZN
                           => n5345);
   U5955 : AOI22_X1 port map( A1 => n5340, A2 => fromRegsPortxREG_FILE_07xx31x,
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_21xx31x, ZN
                           => n5344);
   U5956 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_16xx31x,
                           B1 => n5341, B2 => fromRegsPortxREG_FILE_15xx31x, ZN
                           => n5343);
   U5957 : AND4_X1 port map( A1 => n5346, A2 => n5345, A3 => n5344, A4 => n5343
                           , ZN => n5385);
   U5958 : AOI22_X1 port map( A1 => n5348, A2 => fromRegsPortxREG_FILE_29xx31x,
                           B1 => n5347, B2 => fromRegsPortxREG_FILE_17xx31x, ZN
                           => n5358);
   U5959 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_27xx31x,
                           B1 => n5349, B2 => fromRegsPortxREG_FILE_22xx31x, ZN
                           => n5357);
   U5960 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_03xx31x,
                           B1 => n5351, B2 => fromRegsPortxREG_FILE_20xx31x, ZN
                           => n5356);
   U5961 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_04xx31x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_12xx31x, ZN
                           => n5355);
   U5962 : AND4_X1 port map( A1 => n5358, A2 => n5357, A3 => n5356, A4 => n5355
                           , ZN => n5384);
   U5963 : AOI22_X1 port map( A1 => n5360, A2 => fromRegsPortxREG_FILE_25xx31x,
                           B1 => n5359, B2 => fromRegsPortxREG_FILE_06xx31x, ZN
                           => n5370);
   U5964 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_26xx31x,
                           B1 => n5361, B2 => fromRegsPortxREG_FILE_18xx31x, ZN
                           => n5369);
   U5965 : AOI22_X1 port map( A1 => n5364, A2 => fromRegsPortxREG_FILE_19xx31x,
                           B1 => n5363, B2 => fromRegsPortxREG_FILE_13xx31x, ZN
                           => n5368);
   U5966 : AOI22_X1 port map( A1 => n5366, A2 => fromRegsPortxREG_FILE_10xx31x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_14xx31x, ZN
                           => n5367);
   U5967 : AND4_X1 port map( A1 => n5370, A2 => n5369, A3 => n5368, A4 => n5367
                           , ZN => n5383);
   U5968 : AOI22_X1 port map( A1 => n5372, A2 => fromRegsPortxREG_FILE_02xx31x,
                           B1 => n5371, B2 => fromRegsPortxREG_FILE_05xx31x, ZN
                           => n5381);
   U5969 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_28xx31x,
                           B1 => n5373, B2 => fromRegsPortxREG_FILE_24xx31x, ZN
                           => n5380);
   U5970 : NAND2_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_08xx31x,
                           ZN => n5379);
   U5971 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_01xx31x,
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_31xx31x, ZN
                           => n5378);
   U5972 : AND4_X1 port map( A1 => n5381, A2 => n5380, A3 => n5379, A4 => n5378
                           , ZN => n5382);
   U5973 : NAND4_X1 port map( A1 => n5385, A2 => n5384, A3 => n5383, A4 => 
                           n5382, ZN => n7409);
   U5974 : XOR2_X1 port map( A => n5386, B => n7409, Z => n5387);
   U5975 : XOR2_X1 port map( A => DP_OP_679J1_122_3096xn2, B => n5387, Z => 
                           n5392);
   U5976 : OR4_X1 port map( A1 => DP_OP_679J1_122_3096xn88, A2 => 
                           DP_OP_679J1_122_3096xn87, A3 => 
                           DP_OP_679J1_122_3096xn71, A4 => 
                           DP_OP_679J1_122_3096xn69, ZN => n5388);
   U5977 : OR4_X1 port map( A1 => DP_OP_679J1_122_3096xn91, A2 => 
                           DP_OP_679J1_122_3096xn90, A3 => 
                           DP_OP_679J1_122_3096xn89, A4 => n5388, ZN => n5389);
   U5978 : OR4_X1 port map( A1 => DP_OP_679J1_122_3096xn94, A2 => 
                           DP_OP_679J1_122_3096xn93, A3 => 
                           DP_OP_679J1_122_3096xn92, A4 => n5389, ZN => n5390);
   U5979 : OR4_X1 port map( A1 => DP_OP_679J1_122_3096xn97, A2 => 
                           DP_OP_679J1_122_3096xn96, A3 => 
                           DP_OP_679J1_122_3096xn95, A4 => n5390, ZN => n5391);
   U5980 : OR4_X1 port map( A1 => n5392, A2 => DP_OP_679J1_122_3096xn99, A3 => 
                           DP_OP_679J1_122_3096xn98, A4 => n5391, ZN => n5398);
   U5981 : OR4_X1 port map( A1 => DP_OP_679J1_122_3096xn74, A2 => 
                           DP_OP_679J1_122_3096xn73, A3 => 
                           DP_OP_679J1_122_3096xn72, A4 => 
                           DP_OP_679J1_122_3096xn70, ZN => n5393);
   U5982 : OR4_X1 port map( A1 => DP_OP_679J1_122_3096xn77, A2 => 
                           DP_OP_679J1_122_3096xn76, A3 => 
                           DP_OP_679J1_122_3096xn75, A4 => n5393, ZN => n5394);
   U5983 : OR4_X1 port map( A1 => DP_OP_679J1_122_3096xn80, A2 => 
                           DP_OP_679J1_122_3096xn79, A3 => 
                           DP_OP_679J1_122_3096xn78, A4 => n5394, ZN => n5395);
   U5984 : OR4_X1 port map( A1 => DP_OP_679J1_122_3096xn83, A2 => 
                           DP_OP_679J1_122_3096xn82, A3 => 
                           DP_OP_679J1_122_3096xn81, A4 => n5395, ZN => n5396);
   U5985 : OR4_X1 port map( A1 => DP_OP_679J1_122_3096xn86, A2 => 
                           DP_OP_679J1_122_3096xn85, A3 => 
                           DP_OP_679J1_122_3096xn84, A4 => n5396, ZN => n5397);
   U5986 : NOR2_X1 port map( A1 => n5398, A2 => n5397, ZN => n5628);
   U5987 : INV_X1 port map( A => n7409, ZN => n7431);
   U5988 : NOR2_X1 port map( A1 => n7483, A2 => ashr_25xAx30x, ZN => n7324);
   U5989 : NOR2_X1 port map( A1 => n7477, A2 => ashr_25xAx25x, ZN => n7068);
   U5990 : OAI22_X1 port map( A1 => n7473, A2 => ashr_25xAx21x, B1 => n7472, B2
                           => ashr_25xAx20x, ZN => n5422);
   U5991 : AOI22_X1 port map( A1 => n7472, A2 => ashr_25xAx20x, B1 => n7471, B2
                           => ashr_25xAx19x, ZN => n5421);
   U5992 : INV_X1 port map( A => ashr_25xAx15x, ZN => n6789);
   U5993 : AOI22_X1 port map( A1 => n6789, A2 => n6774, B1 => intadd_2xAx3x, B2
                           => n6726, ZN => n5414);
   U5994 : NAND2_X1 port map( A1 => n7462, A2 => ashr_25xAx10x, ZN => n6525);
   U5995 : INV_X1 port map( A => ashr_25xAx9x, ZN => n6505);
   U5996 : NOR2_X1 port map( A1 => n6505, A2 => n6504, ZN => n6502);
   U5997 : NOR2_X1 port map( A1 => n7460, A2 => ashr_25xAx8x, ZN => n6465);
   U5998 : INV_X1 port map( A => ashr_25xAx7x, ZN => n6425);
   U5999 : INV_X1 port map( A => ashr_25xAx6x, ZN => n6357);
   U6000 : AOI22_X1 port map( A1 => n6425, A2 => n6406, B1 => n6357, B2 => 
                           n6353, ZN => n5406);
   U6001 : INV_X1 port map( A => ashr_25xAx5x, ZN => n5993);
   U6002 : NAND2_X1 port map( A1 => n5993, A2 => n5399, ZN => n6327);
   U6003 : NAND2_X1 port map( A1 => n7081, A2 => ashr_25xAx4x, ZN => n6257);
   U6004 : NOR2_X1 port map( A1 => intadd_4xAx0x, A2 => n7263, ZN => n6090);
   U6005 : NOR2_X1 port map( A1 => n7396, A2 => ashr_25xAx0x, ZN => n5683);
   U6006 : NOR2_X1 port map( A1 => n6144, A2 => ashr_25xAx1x, ZN => n6089);
   U6007 : INV_X2 port map( A => n7305, ZN => n7303);
   U6008 : OAI22_X1 port map( A1 => n5683, A2 => n6089, B1 => intadd_4xAx1x, B2
                           => n7303, ZN => n5400);
   U6009 : NAND2_X1 port map( A1 => intadd_4xAx1x, A2 => n7036, ZN => n6129);
   U6010 : NAND2_X1 port map( A1 => intadd_4xAx2x, A2 => n7203, ZN => n6186);
   U6011 : OAI211_X1 port map( C1 => n6090, C2 => n5400, A => n6129, B => n6186
                           , ZN => n5401);
   U6012 : OAI211_X1 port map( C1 => intadd_4xAx2x, C2 => n7203, A => n6257, B 
                           => n5401, ZN => n5402);
   U6013 : OAI211_X1 port map( C1 => n7081, C2 => ashr_25xAx4x, A => n6327, B 
                           => n5402, ZN => n5403);
   U6014 : NAND2_X1 port map( A1 => n7457, A2 => ashr_25xAx5x, ZN => n6316);
   U6015 : OAI211_X1 port map( C1 => n6357, C2 => n6353, A => n5403, B => n6316
                           , ZN => n5405);
   U6016 : INV_X1 port map( A => ashr_25xAx8x, ZN => n6443);
   U6017 : NOR2_X1 port map( A1 => n6443, A2 => n6445, ZN => n6466);
   U6018 : NOR2_X1 port map( A1 => n6425, A2 => n6406, ZN => n5404);
   U6019 : AOI211_X1 port map( C1 => n5406, C2 => n5405, A => n6466, B => n5404
                           , ZN => n5407);
   U6020 : AOI211_X1 port map( C1 => n6505, C2 => n6504, A => n6465, B => n5407
                           , ZN => n5408);
   U6021 : OAI22_X1 port map( A1 => n6502, A2 => n5408, B1 => n7462, B2 => 
                           ashr_25xAx10x, ZN => n5409);
   U6022 : AOI22_X1 port map( A1 => intadd_2xAx0x, A2 => n6616, B1 => n6525, B2
                           => n5409, ZN => n5411);
   U6023 : OAI22_X1 port map( A1 => intadd_2xAx0x, A2 => n6616, B1 => 
                           intadd_2xAx1x, B2 => n6658, ZN => n5410);
   U6024 : NAND2_X1 port map( A1 => intadd_2xAx1x, A2 => n6658, ZN => n6645);
   U6025 : NAND2_X1 port map( A1 => intadd_2xAx2x, A2 => n6702, ZN => n6690);
   U6026 : OAI211_X1 port map( C1 => n5411, C2 => n5410, A => n6645, B => n6690
                           , ZN => n5412);
   U6027 : NAND2_X1 port map( A1 => n7465, A2 => ashr_25xAx13x, ZN => n6689);
   U6028 : OAI211_X1 port map( C1 => intadd_2xAx3x, C2 => n6726, A => n5412, B 
                           => n6689, ZN => n5413);
   U6029 : AOI22_X1 port map( A1 => n7467, A2 => ashr_25xAx15x, B1 => n5414, B2
                           => n5413, ZN => n5415);
   U6030 : NAND2_X1 port map( A1 => n7468, A2 => ashr_25xAx16x, ZN => n6806);
   U6031 : NOR2_X1 port map( A1 => n7469, A2 => ashr_25xAx17x, ZN => n6831);
   U6032 : NOR2_X1 port map( A1 => n7468, A2 => ashr_25xAx16x, ZN => n6807);
   U6033 : AOI211_X1 port map( C1 => n5415, C2 => n6806, A => n6831, B => n6807
                           , ZN => n5417);
   U6034 : OAI22_X1 port map( A1 => intadd_1xAx0x, A2 => n6835, B1 => 
                           intadd_1xAx1x, B2 => n6891, ZN => n5416);
   U6035 : NAND2_X1 port map( A1 => intadd_1xAx1x, A2 => n6891, ZN => n6885);
   U6036 : NAND2_X1 port map( A1 => intadd_1xAx2x, A2 => n6918, ZN => n6917);
   U6037 : OAI211_X1 port map( C1 => n5417, C2 => n5416, A => n6885, B => n6917
                           , ZN => n5420);
   U6038 : OAI22_X1 port map( A1 => intadd_1xAx4x, A2 => n5717, B1 => 
                           intadd_1xAx5x, B2 => n6986, ZN => n5418);
   U6039 : AOI21_X1 port map( B1 => n7475, B2 => ashr_25xAx23x, A => n5418, ZN 
                           => n5419);
   U6040 : OAI221_X1 port map( B1 => n5422, B2 => n5421, C1 => n5422, C2 => 
                           n5420, A => n5419, ZN => n5424);
   U6041 : NOR2_X1 port map( A1 => n7475, A2 => ashr_25xAx23x, ZN => n7034);
   U6042 : NOR2_X1 port map( A1 => n7474, A2 => ashr_25xAx22x, ZN => n7004);
   U6043 : OAI22_X1 port map( A1 => intadd_1xAx6x, A2 => n7028, B1 => n7034, B2
                           => n7004, ZN => n5423);
   U6044 : AOI22_X1 port map( A1 => n7476, A2 => ashr_25xAx24x, B1 => n5424, B2
                           => n5423, ZN => n5425);
   U6045 : AOI211_X1 port map( C1 => intadd_1xAx7x, C2 => n5744, A => n7068, B 
                           => n5425, ZN => n5430);
   U6046 : INV_X1 port map( A => ashr_25xAx27x, ZN => n7180);
   U6047 : INV_X1 port map( A => ashr_25xAx26x, ZN => n7162);
   U6048 : AOI22_X1 port map( A1 => n7180, A2 => n7179, B1 => n7162, B2 => 
                           n7114, ZN => n5429);
   U6049 : INV_X1 port map( A => ashr_25xAx25x, ZN => n7122);
   U6050 : OAI22_X1 port map( A1 => n7162, A2 => n7114, B1 => n7122, B2 => 
                           n7093, ZN => n5428);
   U6051 : NAND2_X1 port map( A1 => n7481, A2 => ashr_25xAx29x, ZN => n5426);
   U6052 : NAND2_X1 port map( A1 => n7479, A2 => ashr_25xAx27x, ZN => n7177);
   U6053 : OAI211_X1 port map( C1 => intadd_3xAx0x, C2 => n7237, A => n5426, B 
                           => n7177, ZN => n5427);
   U6054 : AOI221_X1 port map( B1 => n5430, B2 => n5429, C1 => n5428, C2 => 
                           n5429, A => n5427, ZN => n5431);
   U6055 : AOI211_X1 port map( C1 => intadd_3xAx1x, C2 => n7247, A => n7324, B 
                           => n5431, ZN => n5433);
   U6056 : OAI211_X1 port map( C1 => intadd_3xAx1x, C2 => n7247, A => 
                           intadd_3xAx0x, B => n7237, ZN => n5432);
   U6057 : AOI22_X1 port map( A1 => n7483, A2 => ashr_25xAx30x, B1 => n5433, B2
                           => n5432, ZN => n5436);
   U6058 : INV_X1 port map( A => n7384, ZN => n7485);
   U6059 : NAND2_X1 port map( A1 => n7485, A2 => n7409, ZN => n5434);
   U6060 : AOI22_X1 port map( A1 => n7431, A2 => n7384, B1 => n5436, B2 => 
                           n5434, ZN => n5633);
   U6061 : NAND2_X1 port map( A1 => n7431, A2 => n7384, ZN => n5435);
   U6062 : AOI22_X1 port map( A1 => n5436, A2 => n5435, B1 => n7485, B2 => 
                           n7409, ZN => n5632);
   U6063 : AOI221_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(13), B2 => 
                           n5633, C1 => n6703, C2 => n5632, A => n6751, ZN => 
                           n5437);
   U6064 : AOI21_X1 port map( B1 => n5976, B2 => n5628, A => n5437, ZN => n5438
                           );
   U6065 : CLKBUF_X1 port map( A => n5657, Z => n5619);
   U6066 : INV_X2 port map( A => n5619, ZN => n5767);
   U6067 : NAND2_X1 port map( A1 => IF_ISAxpcReg_signal_2_port, A2 => 
                           IF_ISAxpcReg_signal_3_port, ZN => n5615);
   U6068 : INV_X1 port map( A => n5615, ZN => n5611);
   U6069 : NAND2_X1 port map( A1 => n5611, A2 => IF_ISAxpcReg_signal_4_port, ZN
                           => n5610);
   U6070 : INV_X1 port map( A => n5610, ZN => n5604);
   U6071 : NAND2_X1 port map( A1 => n5604, A2 => IF_ISAxpcReg_signal_5_port, ZN
                           => n5603);
   U6072 : NOR2_X1 port map( A1 => n5603, A2 => n7539, ZN => n5598);
   U6073 : NAND2_X1 port map( A1 => n5598, A2 => IF_ISAxpcReg_signal_7_port, ZN
                           => n5591);
   U6074 : NOR2_X1 port map( A1 => n5591, A2 => n7540, ZN => n5584);
   U6075 : NAND2_X1 port map( A1 => n5584, A2 => IF_ISAxpcReg_signal_9_port, ZN
                           => n5577);
   U6076 : NOR2_X1 port map( A1 => n5577, A2 => n7541, ZN => n5570);
   U6077 : NAND2_X1 port map( A1 => n5570, A2 => IF_ISAxpcReg_signal_11_port, 
                           ZN => n5563);
   U6078 : INV_X1 port map( A => n5563, ZN => n5439);
   U6079 : AND2_X1 port map( A1 => n5439, A2 => IF_ISAxpcReg_signal_12_port, ZN
                           => n5558);
   U6080 : NAND2_X1 port map( A1 => n5558, A2 => IF_ISAxpcReg_signal_13_port, 
                           ZN => n5553);
   U6081 : INV_X1 port map( A => n5553, ZN => n5547);
   U6082 : NAND2_X1 port map( A1 => n5547, A2 => IF_ISAxpcReg_signal_14_port, 
                           ZN => n5546);
   U6083 : INV_X1 port map( A => n5546, ZN => n5541);
   U6084 : NAND2_X1 port map( A1 => n5541, A2 => IF_ISAxpcReg_signal_15_port, 
                           ZN => n5540);
   U6085 : INV_X1 port map( A => n5540, ZN => n5536);
   U6086 : NAND2_X1 port map( A1 => n5536, A2 => IF_ISAxpcReg_signal_16_port, 
                           ZN => n5535);
   U6087 : INV_X1 port map( A => n5535, ZN => n5529);
   U6088 : NAND2_X1 port map( A1 => n5529, A2 => IF_ISAxpcReg_signal_17_port, 
                           ZN => n5528);
   U6089 : INV_X1 port map( A => n5528, ZN => n5522);
   U6090 : NAND2_X1 port map( A1 => n5522, A2 => IF_ISAxpcReg_signal_18_port, 
                           ZN => n5521);
   U6091 : INV_X1 port map( A => n5521, ZN => n5515);
   U6092 : NAND2_X1 port map( A1 => n5515, A2 => IF_ISAxpcReg_signal_19_port, 
                           ZN => n5514);
   U6093 : INV_X1 port map( A => n5514, ZN => n5509);
   U6094 : NAND2_X1 port map( A1 => n5509, A2 => IF_ISAxpcReg_signal_20_port, 
                           ZN => n5508);
   U6095 : INV_X1 port map( A => n5508, ZN => n5502);
   U6096 : NAND2_X1 port map( A1 => n5502, A2 => IF_ISAxpcReg_signal_21_port, 
                           ZN => n5501);
   U6097 : INV_X1 port map( A => n5501, ZN => n5495);
   U6098 : NAND2_X1 port map( A1 => n5495, A2 => IF_ISAxpcReg_signal_22_port, 
                           ZN => n5494);
   U6099 : INV_X1 port map( A => n5494, ZN => n5489);
   U6100 : NAND2_X1 port map( A1 => n5489, A2 => IF_ISAxpcReg_signal_23_port, 
                           ZN => n5488);
   U6101 : INV_X1 port map( A => n5488, ZN => n5482);
   U6102 : NAND2_X1 port map( A1 => n5482, A2 => IF_ISAxpcReg_signal_24_port, 
                           ZN => n5481);
   U6103 : INV_X1 port map( A => n5481, ZN => n5474);
   U6104 : NAND2_X1 port map( A1 => n5474, A2 => IF_ISAxpcReg_signal_25_port, 
                           ZN => n5473);
   U6105 : INV_X1 port map( A => n5473, ZN => n5466);
   U6106 : NAND2_X1 port map( A1 => n5466, A2 => IF_ISAxpcReg_signal_26_port, 
                           ZN => n5465);
   U6107 : INV_X1 port map( A => n5465, ZN => n5459);
   U6108 : NAND2_X1 port map( A1 => n5459, A2 => IF_ISAxpcReg_signal_27_port, 
                           ZN => n5458);
   U6109 : INV_X1 port map( A => n5458, ZN => n5453);
   U6110 : NAND2_X1 port map( A1 => n5453, A2 => IF_ISAxpcReg_signal_28_port, 
                           ZN => n5452);
   U6111 : INV_X1 port map( A => n5452, ZN => n5447);
   U6112 : NAND2_X1 port map( A1 => n5447, A2 => IF_ISAxpcReg_signal_29_port, 
                           ZN => n5446);
   U6113 : INV_X1 port map( A => n5446, ZN => n5654);
   U6114 : XOR2_X1 port map( A => n5654, B => IF_ISAxpcReg_signal_30_port, Z =>
                           n7357);
   U6115 : AOI22_X1 port map( A1 => n5767, A2 => n7357, B1 => intadd_0xSUMx28x,
                           B2 => n5619, ZN => n5949);
   U6116 : NOR2_X1 port map( A1 => IF_ISAxsection_2_port, A2 => n7534, ZN => 
                           n7454);
   U6117 : NAND2_X1 port map( A1 => IF_ISAxsection_2_port, A2 => n7534, ZN => 
                           n5982);
   U6118 : INV_X1 port map( A => n5982, ZN => n5645);
   U6119 : NOR2_X1 port map( A1 => n7454, A2 => n5645, ZN => n7449);
   U6120 : OR2_X1 port map( A1 => n5761, A2 => fromMemoryPortxLOADEDDATAx(6), 
                           ZN => n5768);
   U6121 : AOI21_X1 port map( B1 => n7449, B2 => n5768, A => rst, ZN => n5607);
   U6122 : CLKBUF_X1 port map( A => n5607, Z => n5659);
   U6123 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(12), A2 => n5440
                           , ZN => n5665);
   U6124 : INV_X1 port map( A => n5665, ZN => n5626);
   U6125 : NAND2_X1 port map( A1 => n5767, A2 => n5441, ZN => n5764);
   U6126 : CLKBUF_X1 port map( A => n5764, Z => n5585);
   U6127 : INV_X1 port map( A => n5585, ZN => n5656);
   U6128 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx28x, B1 => n7357,
                           B2 => n5585, ZN => n5952);
   U6129 : INV_X1 port map( A => n5952, ZN => n5442);
   U6130 : AOI22_X1 port map( A1 => n7357, A2 => n5659, B1 => n5626, B2 => 
                           n5442, ZN => n5445);
   U6131 : NAND2_X1 port map( A1 => n5848, A2 => n7531, ZN => n5979);
   U6132 : NOR3_X1 port map( A1 => n5769, A2 => n5760, A3 => n5979, ZN => n5567
                           );
   U6133 : CLKBUF_X1 port map( A => n5567, Z => n5662);
   U6134 : NOR3_X1 port map( A1 => n5957, A2 => n5769, A3 => n5761, ZN => n5661
                           );
   U6135 : INV_X1 port map( A => intadd_3xSUMx2x, ZN => n5443);
   U6136 : AOI22_X1 port map( A1 => intadd_0xSUMx28x, A2 => n5662, B1 => n5661,
                           B2 => n5443, ZN => n5444);
   U6137 : OAI211_X1 port map( C1 => n5624, C2 => n5949, A => n5445, B => n5444
                           , ZN => n7554);
   U6138 : OAI21_X1 port map( B1 => n5447, B2 => IF_ISAxpcReg_signal_29_port, A
                           => n5446, ZN => n5948);
   U6139 : INV_X1 port map( A => n5948, ZN => n7290);
   U6140 : AOI22_X1 port map( A1 => n5767, A2 => n7290, B1 => intadd_0xSUMx27x,
                           B2 => n5657, ZN => n5944);
   U6141 : INV_X1 port map( A => n5585, ZN => n5765);
   U6142 : AOI22_X1 port map( A1 => n5765, A2 => intadd_0xSUMx27x, B1 => n7290,
                           B2 => n5585, ZN => n5947);
   U6143 : INV_X1 port map( A => n5947, ZN => n5448);
   U6144 : AOI22_X1 port map( A1 => n7290, A2 => n5659, B1 => n5626, B2 => 
                           n5448, ZN => n5451);
   U6145 : INV_X1 port map( A => n5661, ZN => n5579);
   U6146 : INV_X1 port map( A => n5579, ZN => n5621);
   U6147 : INV_X1 port map( A => intadd_3xSUMx1x, ZN => n5449);
   U6148 : AOI22_X1 port map( A1 => intadd_0xSUMx27x, A2 => n5662, B1 => n5621,
                           B2 => n5449, ZN => n5450);
   U6149 : OAI211_X1 port map( C1 => n5624, C2 => n5944, A => n5451, B => n5450
                           , ZN => n7555);
   U6150 : OAI21_X1 port map( B1 => n5453, B2 => IF_ISAxpcReg_signal_28_port, A
                           => n5452, ZN => n5943);
   U6151 : INV_X1 port map( A => n5943, ZN => n7243);
   U6152 : AOI22_X1 port map( A1 => n5767, A2 => n7243, B1 => intadd_0xSUMx26x,
                           B2 => n5657, ZN => n5938);
   U6153 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx26x, B1 => n7243,
                           B2 => n5764, ZN => n5939);
   U6154 : INV_X1 port map( A => n5939, ZN => n5454);
   U6155 : AOI22_X1 port map( A1 => n7243, A2 => n5659, B1 => n5626, B2 => 
                           n5454, ZN => n5457);
   U6156 : INV_X1 port map( A => intadd_3xSUMx0x, ZN => n5455);
   U6157 : AOI22_X1 port map( A1 => intadd_0xSUMx26x, A2 => n5662, B1 => n5661,
                           B2 => n5455, ZN => n5456);
   U6158 : OAI211_X1 port map( C1 => n5624, C2 => n5938, A => n5457, B => n5456
                           , ZN => n7556);
   U6159 : OAI21_X1 port map( B1 => n5459, B2 => IF_ISAxpcReg_signal_27_port, A
                           => n5458, ZN => n5936);
   U6160 : INV_X1 port map( A => n5936, ZN => n7199);
   U6161 : AOI22_X1 port map( A1 => n5765, A2 => intadd_0xSUMx25x, B1 => n7199,
                           B2 => n5585, ZN => n5935);
   U6162 : INV_X1 port map( A => intadd_0xSUMx25x, ZN => n7181);
   U6163 : AOI22_X1 port map( A1 => n5767, A2 => n5936, B1 => n7181, B2 => 
                           n5657, ZN => n5931);
   U6164 : AOI22_X1 port map( A1 => n7199, A2 => n5659, B1 => n5931, B2 => 
                           n5658, ZN => n5464);
   U6165 : NOR2_X1 port map( A1 => n7122, A2 => add_x_26xBx25x, ZN => n6025);
   U6166 : AOI21_X1 port map( B1 => n7122, B2 => add_x_26xBx25x, A => n6025, ZN
                           => n5477);
   U6167 : NOR2_X1 port map( A1 => n5477, A2 => intadd_1xn1, ZN => n5460);
   U6168 : AOI21_X1 port map( B1 => ashr_25xAx25x, B2 => add_x_26xBx25x, A => 
                           n5460, ZN => n5469);
   U6169 : INV_X1 port map( A => n5461, ZN => n5937);
   U6170 : OAI22_X1 port map( A1 => ashr_25xAx27x, A2 => add_x_26xBx27x, B1 => 
                           n5462, B2 => n7180, ZN => n7178);
   U6171 : XNOR2_X1 port map( A => n5937, B => n7178, ZN => n5933);
   U6172 : AOI22_X1 port map( A1 => intadd_0xSUMx25x, A2 => n5662, B1 => n5621,
                           B2 => n5933, ZN => n5463);
   U6173 : OAI211_X1 port map( C1 => n5935, C2 => n5665, A => n5464, B => n5463
                           , ZN => n7557);
   U6174 : OAI21_X1 port map( B1 => n5466, B2 => IF_ISAxpcReg_signal_26_port, A
                           => n5465, ZN => n7111);
   U6175 : INV_X1 port map( A => n7111, ZN => n5468);
   U6176 : AOI22_X1 port map( A1 => n5767, A2 => n5468, B1 => intadd_0xSUMx24x,
                           B2 => n5657, ZN => n5925);
   U6177 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx24x, B1 => n5468,
                           B2 => n5585, ZN => n5926);
   U6178 : INV_X1 port map( A => n5926, ZN => n5467);
   U6179 : AOI22_X1 port map( A1 => n5468, A2 => n5659, B1 => n5626, B2 => 
                           n5467, ZN => n5472);
   U6180 : FA_X1 port map( A => n7162, B => n7120, CI => n5469, CO => n5461, S 
                           => n5927);
   U6181 : INV_X1 port map( A => n5927, ZN => n5470);
   U6182 : AOI22_X1 port map( A1 => intadd_0xSUMx24x, A2 => n5662, B1 => n5661,
                           B2 => n5470, ZN => n5471);
   U6183 : OAI211_X1 port map( C1 => n5624, C2 => n5925, A => n5472, B => n5471
                           , ZN => n7558);
   U6184 : OAI21_X1 port map( B1 => n5474, B2 => IF_ISAxpcReg_signal_25_port, A
                           => n5473, ZN => n7073);
   U6185 : INV_X1 port map( A => n7073, ZN => n5476);
   U6186 : AOI22_X1 port map( A1 => n5767, A2 => n5476, B1 => intadd_0xSUMx23x,
                           B2 => n5619, ZN => n5919);
   U6187 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx23x, B1 => n5476,
                           B2 => n5764, ZN => n5920);
   U6188 : INV_X1 port map( A => n5920, ZN => n5475);
   U6189 : AOI22_X1 port map( A1 => n5476, A2 => n5659, B1 => n5626, B2 => 
                           n5475, ZN => n5480);
   U6190 : XNOR2_X1 port map( A => n5477, B => intadd_1xn1, ZN => n5921);
   U6191 : INV_X1 port map( A => n5921, ZN => n5478);
   U6192 : AOI22_X1 port map( A1 => intadd_0xSUMx23x, A2 => n5662, B1 => n5478,
                           B2 => n5661, ZN => n5479);
   U6193 : OAI211_X1 port map( C1 => n5624, C2 => n5919, A => n5480, B => n5479
                           , ZN => n7559);
   U6194 : OAI21_X1 port map( B1 => n5482, B2 => IF_ISAxpcReg_signal_24_port, A
                           => n5481, ZN => n5918);
   U6195 : INV_X1 port map( A => n5918, ZN => n5484);
   U6196 : AOI22_X1 port map( A1 => n5767, A2 => n5484, B1 => intadd_0xSUMx22x,
                           B2 => n5657, ZN => n5913);
   U6197 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx22x, B1 => n5484,
                           B2 => n5764, ZN => n5914);
   U6198 : INV_X1 port map( A => n5914, ZN => n5483);
   U6199 : AOI22_X1 port map( A1 => n5484, A2 => n5659, B1 => n5626, B2 => 
                           n5483, ZN => n5487);
   U6200 : INV_X1 port map( A => intadd_1xSUMx7x, ZN => n5485);
   U6201 : AOI22_X1 port map( A1 => intadd_0xSUMx22x, A2 => n5662, B1 => n5621,
                           B2 => n5485, ZN => n5486);
   U6202 : OAI211_X1 port map( C1 => n5624, C2 => n5913, A => n5487, B => n5486
                           , ZN => n7560);
   U6203 : OAI21_X1 port map( B1 => n5489, B2 => IF_ISAxpcReg_signal_23_port, A
                           => n5488, ZN => n5912);
   U6204 : INV_X1 port map( A => n5912, ZN => n7033);
   U6205 : AOI22_X1 port map( A1 => n5767, A2 => n7033, B1 => intadd_0xSUMx21x,
                           B2 => n5657, ZN => n5908);
   U6206 : AOI22_X1 port map( A1 => n5765, A2 => intadd_0xSUMx21x, B1 => n7033,
                           B2 => n5764, ZN => n5911);
   U6207 : INV_X1 port map( A => n5911, ZN => n5490);
   U6208 : AOI22_X1 port map( A1 => n7033, A2 => n5659, B1 => n5626, B2 => 
                           n5490, ZN => n5493);
   U6209 : INV_X1 port map( A => intadd_1xSUMx6x, ZN => n5491);
   U6210 : AOI22_X1 port map( A1 => intadd_0xSUMx21x, A2 => n5662, B1 => n5621,
                           B2 => n5491, ZN => n5492);
   U6211 : OAI211_X1 port map( C1 => n5624, C2 => n5908, A => n5493, B => n5492
                           , ZN => n7561);
   U6212 : OAI21_X1 port map( B1 => n5495, B2 => IF_ISAxpcReg_signal_22_port, A
                           => n5494, ZN => n7014);
   U6213 : INV_X1 port map( A => n7014, ZN => n5497);
   U6214 : AOI22_X1 port map( A1 => n5767, A2 => n5497, B1 => intadd_0xSUMx20x,
                           B2 => n5657, ZN => n5903);
   U6215 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx20x, B1 => n5497,
                           B2 => n5764, ZN => n5904);
   U6216 : INV_X1 port map( A => n5904, ZN => n5496);
   U6217 : AOI22_X1 port map( A1 => n5497, A2 => n5659, B1 => n5626, B2 => 
                           n5496, ZN => n5500);
   U6218 : INV_X1 port map( A => intadd_1xSUMx5x, ZN => n5498);
   U6219 : AOI22_X1 port map( A1 => intadd_0xSUMx20x, A2 => n5662, B1 => n5621,
                           B2 => n5498, ZN => n5499);
   U6220 : OAI211_X1 port map( C1 => n5624, C2 => n5903, A => n5500, B => n5499
                           , ZN => n7562);
   U6221 : OAI21_X1 port map( B1 => n5502, B2 => IF_ISAxpcReg_signal_21_port, A
                           => n5501, ZN => n5902);
   U6222 : INV_X1 port map( A => n5902, ZN => n5504);
   U6223 : AOI22_X1 port map( A1 => n5767, A2 => n5504, B1 => intadd_0xSUMx19x,
                           B2 => n5657, ZN => n5897);
   U6224 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx19x, B1 => n5504,
                           B2 => n5764, ZN => n5898);
   U6225 : INV_X1 port map( A => n5898, ZN => n5503);
   U6226 : AOI22_X1 port map( A1 => n5504, A2 => n5659, B1 => n5626, B2 => 
                           n5503, ZN => n5507);
   U6227 : INV_X1 port map( A => intadd_1xSUMx4x, ZN => n5505);
   U6228 : AOI22_X1 port map( A1 => intadd_0xSUMx19x, A2 => n5662, B1 => n5621,
                           B2 => n5505, ZN => n5506);
   U6229 : OAI211_X1 port map( C1 => n5624, C2 => n5897, A => n5507, B => n5506
                           , ZN => n7563);
   U6230 : OAI21_X1 port map( B1 => n5509, B2 => IF_ISAxpcReg_signal_20_port, A
                           => n5508, ZN => n5896);
   U6231 : INV_X1 port map( A => n5896, ZN => n6955);
   U6232 : AOI22_X1 port map( A1 => n5767, A2 => n6955, B1 => intadd_0xSUMx18x,
                           B2 => n5657, ZN => n5891);
   U6233 : AOI22_X1 port map( A1 => n5765, A2 => intadd_0xSUMx18x, B1 => n6955,
                           B2 => n5764, ZN => n5892);
   U6234 : INV_X1 port map( A => n5892, ZN => n5510);
   U6235 : AOI22_X1 port map( A1 => n6955, A2 => n5659, B1 => n5626, B2 => 
                           n5510, ZN => n5513);
   U6236 : INV_X1 port map( A => intadd_1xSUMx3x, ZN => n5511);
   U6237 : AOI22_X1 port map( A1 => intadd_0xSUMx18x, A2 => n5662, B1 => n5621,
                           B2 => n5511, ZN => n5512);
   U6238 : OAI211_X1 port map( C1 => n5624, C2 => n5891, A => n5513, B => n5512
                           , ZN => n7564);
   U6239 : OAI21_X1 port map( B1 => n5515, B2 => IF_ISAxpcReg_signal_19_port, A
                           => n5514, ZN => n6923);
   U6240 : INV_X1 port map( A => n6923, ZN => n5517);
   U6241 : AOI22_X1 port map( A1 => n5767, A2 => n5517, B1 => intadd_0xSUMx17x,
                           B2 => n5657, ZN => n5885);
   U6242 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx17x, B1 => n5517,
                           B2 => n5764, ZN => n5887);
   U6243 : INV_X1 port map( A => n5887, ZN => n5516);
   U6244 : AOI22_X1 port map( A1 => n5517, A2 => n5659, B1 => n5626, B2 => 
                           n5516, ZN => n5520);
   U6245 : INV_X1 port map( A => intadd_1xSUMx2x, ZN => n5518);
   U6246 : AOI22_X1 port map( A1 => intadd_0xSUMx17x, A2 => n5567, B1 => n5621,
                           B2 => n5518, ZN => n5519);
   U6247 : OAI211_X1 port map( C1 => n5624, C2 => n5885, A => n5520, B => n5519
                           , ZN => n7565);
   U6248 : OAI21_X1 port map( B1 => n5522, B2 => IF_ISAxpcReg_signal_18_port, A
                           => n5521, ZN => n6889);
   U6249 : INV_X1 port map( A => n6889, ZN => n5524);
   U6250 : AOI22_X1 port map( A1 => n5767, A2 => n5524, B1 => intadd_0xSUMx16x,
                           B2 => n5657, ZN => n5881);
   U6251 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx16x, B1 => n5524,
                           B2 => n5764, ZN => n5884);
   U6252 : INV_X1 port map( A => n5884, ZN => n5523);
   U6253 : AOI22_X1 port map( A1 => n5524, A2 => n5659, B1 => n5626, B2 => 
                           n5523, ZN => n5527);
   U6254 : INV_X1 port map( A => intadd_1xSUMx1x, ZN => n5525);
   U6255 : AOI22_X1 port map( A1 => intadd_0xSUMx16x, A2 => n5567, B1 => n5621,
                           B2 => n5525, ZN => n5526);
   U6256 : OAI211_X1 port map( C1 => n5624, C2 => n5881, A => n5527, B => n5526
                           , ZN => n7566);
   U6257 : OAI21_X1 port map( B1 => n5529, B2 => IF_ISAxpcReg_signal_17_port, A
                           => n5528, ZN => n6834);
   U6258 : INV_X1 port map( A => n6834, ZN => n5531);
   U6259 : AOI22_X1 port map( A1 => n5767, A2 => n5531, B1 => intadd_0xSUMx15x,
                           B2 => n5657, ZN => n5877);
   U6260 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx15x, B1 => n5531,
                           B2 => n5764, ZN => n5880);
   U6261 : INV_X1 port map( A => n5880, ZN => n5530);
   U6262 : AOI22_X1 port map( A1 => n5531, A2 => n5659, B1 => n5626, B2 => 
                           n5530, ZN => n5534);
   U6263 : INV_X1 port map( A => intadd_1xSUMx0x, ZN => n5532);
   U6264 : AOI22_X1 port map( A1 => intadd_0xSUMx15x, A2 => n5662, B1 => n5621,
                           B2 => n5532, ZN => n5533);
   U6265 : OAI211_X1 port map( C1 => n5624, C2 => n5877, A => n5534, B => n5533
                           , ZN => n7567);
   U6266 : OAI21_X1 port map( B1 => n5536, B2 => IF_ISAxpcReg_signal_16_port, A
                           => n5535, ZN => n5875);
   U6267 : INV_X1 port map( A => n5875, ZN => n6804);
   U6268 : AOI22_X1 port map( A1 => n5767, A2 => n6804, B1 => intadd_0xSUMx14x,
                           B2 => n5657, ZN => n5870);
   U6269 : INV_X1 port map( A => ashr_25xAx16x, ZN => n6802);
   U6270 : AOI22_X1 port map( A1 => n6802, A2 => n6811, B1 => add_x_26xBx16x, 
                           B2 => ashr_25xAx16x, ZN => n6803);
   U6271 : AOI22_X1 port map( A1 => n6789, A2 => add_x_26xBx15x, B1 => n6778, 
                           B2 => ashr_25xAx15x, ZN => n6779);
   U6272 : OAI22_X1 port map( A1 => n6789, A2 => n6778, B1 => n6779, B2 => 
                           intadd_2xn1, ZN => n5876);
   U6273 : XOR2_X1 port map( A => n6803, B => n5876, Z => n5869);
   U6274 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx14x, B1 => n6804,
                           B2 => n5764, ZN => n5871);
   U6275 : INV_X1 port map( A => n5871, ZN => n5537);
   U6276 : AOI22_X1 port map( A1 => n5869, A2 => n5621, B1 => n5626, B2 => 
                           n5537, ZN => n5539);
   U6277 : AOI22_X1 port map( A1 => n6804, A2 => n5659, B1 => intadd_0xSUMx14x,
                           B2 => n5662, ZN => n5538);
   U6278 : OAI211_X1 port map( C1 => n5624, C2 => n5870, A => n5539, B => n5538
                           , ZN => n7568);
   U6279 : OAI21_X1 port map( B1 => n5541, B2 => IF_ISAxpcReg_signal_15_port, A
                           => n5540, ZN => n6777);
   U6280 : INV_X1 port map( A => n6777, ZN => n5543);
   U6281 : AOI22_X1 port map( A1 => n5767, A2 => n5543, B1 => intadd_0xSUMx13x,
                           B2 => n5657, ZN => n5864);
   U6282 : XOR2_X1 port map( A => n6779, B => intadd_2xn1, Z => n5863);
   U6283 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx13x, B1 => n5543,
                           B2 => n5764, ZN => n5865);
   U6284 : INV_X1 port map( A => n5865, ZN => n5542);
   U6285 : AOI22_X1 port map( A1 => n5863, A2 => n5621, B1 => n5626, B2 => 
                           n5542, ZN => n5545);
   U6286 : AOI22_X1 port map( A1 => n5543, A2 => n5607, B1 => intadd_0xSUMx13x,
                           B2 => n5662, ZN => n5544);
   U6287 : OAI211_X1 port map( C1 => n5624, C2 => n5864, A => n5545, B => n5544
                           , ZN => n7569);
   U6288 : OAI21_X1 port map( B1 => n5547, B2 => IF_ISAxpcReg_signal_14_port, A
                           => n5546, ZN => n6720);
   U6289 : INV_X1 port map( A => n6720, ZN => n5549);
   U6290 : AOI22_X1 port map( A1 => n5767, A2 => n5549, B1 => intadd_0xSUMx12x,
                           B2 => n5657, ZN => n5859);
   U6291 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx12x, B1 => n5549,
                           B2 => n5585, ZN => n5862);
   U6292 : INV_X1 port map( A => n5862, ZN => n5548);
   U6293 : AOI22_X1 port map( A1 => n5549, A2 => n5607, B1 => n5626, B2 => 
                           n5548, ZN => n5552);
   U6294 : INV_X1 port map( A => intadd_2xSUMx3x, ZN => n5550);
   U6295 : AOI22_X1 port map( A1 => intadd_0xSUMx12x, A2 => n5567, B1 => n5621,
                           B2 => n5550, ZN => n5551);
   U6296 : OAI211_X1 port map( C1 => n5624, C2 => n5859, A => n5552, B => n5551
                           , ZN => n7570);
   U6297 : OAI21_X1 port map( B1 => n5558, B2 => IF_ISAxpcReg_signal_13_port, A
                           => n5553, ZN => n5858);
   U6298 : INV_X1 port map( A => n5858, ZN => n6667);
   U6299 : AOI22_X1 port map( A1 => n5767, A2 => n6667, B1 => intadd_0xSUMx11x,
                           B2 => n5619, ZN => n5853);
   U6300 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx11x, B1 => n6667,
                           B2 => n5585, ZN => n5854);
   U6301 : INV_X1 port map( A => n5854, ZN => n5554);
   U6302 : AOI22_X1 port map( A1 => n6667, A2 => n5607, B1 => n5626, B2 => 
                           n5554, ZN => n5557);
   U6303 : INV_X1 port map( A => intadd_2xSUMx2x, ZN => n5555);
   U6304 : AOI22_X1 port map( A1 => intadd_0xSUMx11x, A2 => n5567, B1 => n5621,
                           B2 => n5555, ZN => n5556);
   U6305 : OAI211_X1 port map( C1 => n5624, C2 => n5853, A => n5557, B => n5556
                           , ZN => n7571);
   U6306 : AOI21_X1 port map( B1 => n5563, B2 => n7543, A => n5558, ZN => n6644
                           );
   U6307 : AOI22_X1 port map( A1 => n5767, A2 => n6644, B1 => intadd_0xSUMx10x,
                           B2 => n5657, ZN => n5846);
   U6308 : INV_X1 port map( A => intadd_0xSUMx10x, ZN => n6643);
   U6309 : INV_X1 port map( A => n6644, ZN => n5559);
   U6310 : AOI22_X1 port map( A1 => n5656, A2 => n6643, B1 => n5559, B2 => 
                           n5764, ZN => n5844);
   U6311 : AOI22_X1 port map( A1 => n6644, A2 => n5607, B1 => n5626, B2 => 
                           n5844, ZN => n5562);
   U6312 : INV_X1 port map( A => intadd_2xSUMx1x, ZN => n5560);
   U6313 : AOI22_X1 port map( A1 => intadd_0xSUMx10x, A2 => n5567, B1 => n5621,
                           B2 => n5560, ZN => n5561);
   U6314 : OAI211_X1 port map( C1 => n5624, C2 => n5846, A => n5562, B => n5561
                           , ZN => n7572);
   U6315 : OAI21_X1 port map( B1 => n5570, B2 => IF_ISAxpcReg_signal_11_port, A
                           => n5563, ZN => n6592);
   U6316 : INV_X1 port map( A => n6592, ZN => n5565);
   U6317 : AOI22_X1 port map( A1 => n5767, A2 => n5565, B1 => intadd_0xSUMx9x, 
                           B2 => n5657, ZN => n5838);
   U6318 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx9x, B1 => n5565, 
                           B2 => n5764, ZN => n5839);
   U6319 : INV_X1 port map( A => n5839, ZN => n5564);
   U6320 : AOI22_X1 port map( A1 => n5565, A2 => n5607, B1 => n5626, B2 => 
                           n5564, ZN => n5569);
   U6321 : INV_X1 port map( A => intadd_2xSUMx0x, ZN => n5566);
   U6322 : AOI22_X1 port map( A1 => intadd_0xSUMx9x, A2 => n5567, B1 => n5621, 
                           B2 => n5566, ZN => n5568);
   U6323 : OAI211_X1 port map( C1 => n5624, C2 => n5838, A => n5569, B => n5568
                           , ZN => n7573);
   U6324 : AOI21_X1 port map( B1 => n5577, B2 => n7541, A => n5570, ZN => n6532
                           );
   U6325 : AOI22_X1 port map( A1 => n5767, A2 => n6532, B1 => intadd_0xSUMx8x, 
                           B2 => n5657, ZN => n5830);
   U6326 : OAI22_X1 port map( A1 => ashr_25xAx9x, A2 => n6500, B1 => 
                           add_x_26xBx9x, B2 => n6505, ZN => n6503);
   U6327 : NOR2_X1 port map( A1 => n6443, A2 => n5586, ZN => n6460);
   U6328 : NOR2_X1 port map( A1 => ashr_25xAx4x, A2 => ashr_25xSHx4x, ZN => 
                           n5571);
   U6329 : NAND2_X1 port map( A1 => ashr_25xAx4x, A2 => ashr_25xSHx4x, ZN => 
                           n6259);
   U6330 : OAI21_X1 port map( B1 => n5571, B2 => intadd_4xn1, A => n6259, ZN =>
                           n5605);
   U6331 : INV_X1 port map( A => n5605, ZN => n5572);
   U6332 : AOI22_X1 port map( A1 => n5993, A2 => add_x_26xBx5x, B1 => n6307, B2
                           => ashr_25xAx5x, ZN => n5606);
   U6333 : INV_X1 port map( A => n5606, ZN => n6296);
   U6334 : AOI22_X1 port map( A1 => n5993, A2 => n6307, B1 => n5572, B2 => 
                           n6296, ZN => n5600);
   U6335 : OAI22_X1 port map( A1 => add_x_26xBx8x, A2 => ashr_25xAx8x, B1 => 
                           n6460, B2 => n5587, ZN => n5578);
   U6336 : AOI22_X1 port map( A1 => n6505, A2 => n6500, B1 => n6503, B2 => 
                           n5578, ZN => n5837);
   U6337 : INV_X1 port map( A => ashr_25xAx10x, ZN => n6553);
   U6338 : NOR2_X1 port map( A1 => n5835, A2 => n6553, ZN => n6565);
   U6339 : AOI21_X1 port map( B1 => n5835, B2 => n6553, A => n6565, ZN => n5573
                           );
   U6340 : INV_X1 port map( A => n5573, ZN => n6537);
   U6341 : XOR2_X1 port map( A => n5837, B => n6537, Z => n5829);
   U6342 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx8x, B1 => n6532, 
                           B2 => n5764, ZN => n5834);
   U6343 : OAI22_X1 port map( A1 => n5829, A2 => n5579, B1 => n5665, B2 => 
                           n5834, ZN => n5574);
   U6344 : INV_X1 port map( A => n5574, ZN => n5576);
   U6345 : AOI22_X1 port map( A1 => intadd_0xSUMx8x, A2 => n5662, B1 => n6532, 
                           B2 => n5659, ZN => n5575);
   U6346 : OAI211_X1 port map( C1 => n5624, C2 => n5830, A => n5576, B => n5575
                           , ZN => n7574);
   U6347 : OAI21_X1 port map( B1 => n5584, B2 => IF_ISAxpcReg_signal_9_port, A 
                           => n5577, ZN => n6495);
   U6348 : INV_X1 port map( A => n6495, ZN => n5581);
   U6349 : AOI22_X1 port map( A1 => n5767, A2 => n5581, B1 => intadd_0xSUMx7x, 
                           B2 => n5657, ZN => n5823);
   U6350 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx7x, B1 => n5581, 
                           B2 => n5764, ZN => n5822);
   U6351 : XOR2_X1 port map( A => n6503, B => n5578, Z => n5824);
   U6352 : OAI22_X1 port map( A1 => n5665, A2 => n5822, B1 => n5579, B2 => 
                           n5824, ZN => n5580);
   U6353 : INV_X1 port map( A => n5580, ZN => n5583);
   U6354 : AOI22_X1 port map( A1 => n5581, A2 => n5607, B1 => intadd_0xSUMx7x, 
                           B2 => n5662, ZN => n5582);
   U6355 : OAI211_X1 port map( C1 => n5624, C2 => n5823, A => n5583, B => n5582
                           , ZN => n7575);
   U6356 : AOI21_X1 port map( B1 => n5591, B2 => n7540, A => n5584, ZN => n6459
                           );
   U6357 : AOI22_X1 port map( A1 => n5767, A2 => n6459, B1 => intadd_0xSUMx6x, 
                           B2 => n5657, ZN => n5816);
   U6358 : AOI22_X1 port map( A1 => n5656, A2 => intadd_0xSUMx6x, B1 => n6459, 
                           B2 => n5585, ZN => n5821);
   U6359 : INV_X1 port map( A => n5821, ZN => n5588);
   U6360 : AOI22_X1 port map( A1 => n6443, A2 => add_x_26xBx8x, B1 => n5586, B2
                           => ashr_25xAx8x, ZN => n6469);
   U6361 : XNOR2_X1 port map( A => n5587, B => n6469, ZN => n5815);
   U6362 : AOI22_X1 port map( A1 => n5626, A2 => n5588, B1 => n5621, B2 => 
                           n5815, ZN => n5590);
   U6363 : AOI22_X1 port map( A1 => intadd_0xSUMx6x, A2 => n5662, B1 => n6459, 
                           B2 => n5659, ZN => n5589);
   U6364 : OAI211_X1 port map( C1 => n5624, C2 => n5816, A => n5590, B => n5589
                           , ZN => n7576);
   U6365 : OR2_X1 port map( A1 => n5598, A2 => IF_ISAxpcReg_signal_7_port, ZN 
                           => n5592);
   U6366 : AND2_X1 port map( A1 => n5592, A2 => n5591, ZN => n5594);
   U6367 : AOI22_X1 port map( A1 => n5765, A2 => intadd_0xSUMx5x, B1 => n5594, 
                           B2 => n5764, ZN => n5811);
   U6368 : INV_X1 port map( A => n5594, ZN => n6419);
   U6369 : INV_X1 port map( A => intadd_0xSUMx5x, ZN => n5593);
   U6370 : AOI22_X1 port map( A1 => n5767, A2 => n6419, B1 => n5593, B2 => 
                           n5657, ZN => n5809);
   U6371 : AOI22_X1 port map( A1 => n5594, A2 => n5607, B1 => n5809, B2 => 
                           n5658, ZN => n5597);
   U6372 : FA_X1 port map( A => ashr_25xAx7x, B => add_x_26xBx7x, CI => n5595, 
                           CO => n5587, S => n5813);
   U6373 : AOI22_X1 port map( A1 => n5813, A2 => n5621, B1 => intadd_0xSUMx5x, 
                           B2 => n5662, ZN => n5596);
   U6374 : OAI211_X1 port map( C1 => n5811, C2 => n5665, A => n5597, B => n5596
                           , ZN => n7577);
   U6375 : AOI21_X1 port map( B1 => n5603, B2 => n7539, A => n5598, ZN => n6362
                           );
   U6376 : AOI22_X1 port map( A1 => n5767, A2 => n6362, B1 => intadd_0xSUMx4x, 
                           B2 => n5657, ZN => n5802);
   U6377 : AOI22_X1 port map( A1 => n5765, A2 => intadd_0xSUMx4x, B1 => n6362, 
                           B2 => n5764, ZN => n5807);
   U6378 : INV_X1 port map( A => n5807, ZN => n5599);
   U6379 : AOI22_X1 port map( A1 => n6362, A2 => n5607, B1 => n5626, B2 => 
                           n5599, ZN => n5602);
   U6380 : FA_X1 port map( A => ashr_25xAx6x, B => add_x_26xBx6x, CI => n5600, 
                           CO => n5595, S => n5803);
   U6381 : AOI22_X1 port map( A1 => intadd_0xSUMx4x, A2 => n5662, B1 => n5803, 
                           B2 => n5621, ZN => n5601);
   U6382 : OAI211_X1 port map( C1 => n5624, C2 => n5802, A => n5602, B => n5601
                           , ZN => n7578);
   U6383 : OAI21_X1 port map( B1 => n5604, B2 => IF_ISAxpcReg_signal_5_port, A 
                           => n5603, ZN => n5801);
   U6384 : INV_X1 port map( A => n5801, ZN => n6306);
   U6385 : AOI22_X1 port map( A1 => n5765, A2 => intadd_0xSUMx3x, B1 => n6306, 
                           B2 => n5764, ZN => n5800);
   U6386 : INV_X1 port map( A => intadd_0xSUMx3x, ZN => n6315);
   U6387 : AOI22_X1 port map( A1 => n5767, A2 => n5801, B1 => n6315, B2 => 
                           n5657, ZN => n5797);
   U6388 : XNOR2_X1 port map( A => n5606, B => n5605, ZN => n5798);
   U6389 : AOI22_X1 port map( A1 => n5797, A2 => n5658, B1 => n5621, B2 => 
                           n5798, ZN => n5609);
   U6390 : AOI22_X1 port map( A1 => n6306, A2 => n5607, B1 => intadd_0xSUMx3x, 
                           B2 => n5662, ZN => n5608);
   U6391 : OAI211_X1 port map( C1 => n5800, C2 => n5665, A => n5609, B => n5608
                           , ZN => n7579);
   U6392 : OAI21_X1 port map( B1 => n5611, B2 => IF_ISAxpcReg_signal_4_port, A 
                           => n5610, ZN => n6258);
   U6393 : INV_X1 port map( A => n6258, ZN => n5790);
   U6394 : AOI22_X1 port map( A1 => n5767, A2 => n5790, B1 => intadd_0xSUMx2x, 
                           B2 => n5657, ZN => n5792);
   U6395 : INV_X1 port map( A => intadd_0xSUMx2x, ZN => n6285);
   U6396 : AOI22_X1 port map( A1 => n5765, A2 => n6285, B1 => n6258, B2 => 
                           n5764, ZN => n5791);
   U6397 : OAI21_X1 port map( B1 => ashr_25xSHx4x, B2 => ashr_25xAx4x, A => 
                           n6259, ZN => n6284);
   U6398 : XNOR2_X1 port map( A => intadd_4xn1, B => n6284, ZN => n5796);
   U6399 : INV_X1 port map( A => n5796, ZN => n5612);
   U6400 : AOI22_X1 port map( A1 => n5626, A2 => n5791, B1 => n5621, B2 => 
                           n5612, ZN => n5614);
   U6401 : AOI22_X1 port map( A1 => intadd_0xSUMx2x, A2 => n5662, B1 => n5790, 
                           B2 => n5659, ZN => n5613);
   U6402 : OAI211_X1 port map( C1 => n5624, C2 => n5792, A => n5614, B => n5613
                           , ZN => n7580);
   U6403 : OAI21_X1 port map( B1 => IF_ISAxpcReg_signal_2_port, B2 => 
                           IF_ISAxpcReg_signal_3_port, A => n5615, ZN => n6213)
                           ;
   U6404 : INV_X1 port map( A => n6213, ZN => n5784);
   U6405 : AOI22_X1 port map( A1 => n5767, A2 => n5784, B1 => intadd_0xSUMx1x, 
                           B2 => n5619, ZN => n5786);
   U6406 : INV_X1 port map( A => intadd_0xSUMx1x, ZN => n6239);
   U6407 : AOI22_X1 port map( A1 => n5765, A2 => n6239, B1 => n6213, B2 => 
                           n5764, ZN => n5785);
   U6408 : AOI22_X1 port map( A1 => n5784, A2 => n5659, B1 => n5785, B2 => 
                           n5626, ZN => n5618);
   U6409 : INV_X1 port map( A => intadd_4xSUMx2x, ZN => n5616);
   U6410 : AOI22_X1 port map( A1 => intadd_0xSUMx1x, A2 => n5662, B1 => n5661, 
                           B2 => n5616, ZN => n5617);
   U6411 : OAI211_X1 port map( C1 => n5624, C2 => n5786, A => n5618, B => n5617
                           , ZN => n7581);
   U6412 : INV_X1 port map( A => intadd_0xSUMx0x, ZN => n6117);
   U6413 : AOI22_X1 port map( A1 => n5765, A2 => n6117, B1 => 
                           IF_ISAxpcReg_signal_2_port, B2 => n5764, ZN => n5779
                           );
   U6414 : AOI22_X1 port map( A1 => n5767, A2 => n7542, B1 => n5619, B2 => 
                           intadd_0xSUMx0x, ZN => n5780);
   U6415 : INV_X1 port map( A => intadd_4xSUMx1x, ZN => n5620);
   U6416 : AOI22_X1 port map( A1 => intadd_0xSUMx0x, A2 => n5662, B1 => n5621, 
                           B2 => n5620, ZN => n5623);
   U6417 : NAND2_X1 port map( A1 => n5659, A2 => n7542, ZN => n5622);
   U6418 : OAI211_X1 port map( C1 => n5780, C2 => n5624, A => n5623, B => n5622
                           , ZN => n5625);
   U6419 : AOI21_X1 port map( B1 => n5779, B2 => n5626, A => n5625, ZN => n5627
                           );
   U6420 : INV_X1 port map( A => n5627, ZN => n7582);
   U6421 : NOR2_X1 port map( A1 => intadd_4xBx0x, A2 => n7538, ZN => 
                           intadd_0xCI);
   U6422 : INV_X1 port map( A => n5628, ZN => n5634);
   U6423 : INV_X1 port map( A => n5629, ZN => n5630);
   U6424 : INV_X1 port map( A => n5690, ZN => n5724);
   U6425 : NAND3_X1 port map( A1 => n5631, A2 => n5630, A3 => n5724, ZN => 
                           n6040);
   U6426 : OR2_X1 port map( A1 => n5716, A2 => n5690, ZN => n6038);
   U6427 : OAI22_X1 port map( A1 => n5633, A2 => n6040, B1 => n5632, B2 => 
                           n6038, ZN => n6042);
   U6428 : AOI21_X1 port map( B1 => n5634, B2 => n5679, A => n6042, ZN => n5639
                           );
   U6429 : NAND3_X1 port map( A1 => n5639, A2 => n5636, A3 => n5635, ZN => 
                           n5637);
   U6430 : OAI21_X1 port map( B1 => n5639, B2 => n5638, A => n5637, ZN => n5647
                           );
   U6431 : INV_X1 port map( A => n5647, ZN => n5640);
   U6432 : AOI22_X1 port map( A1 => n7454, A2 => IF_ISAxsection_0_port, B1 => 
                           n5641, B2 => n5640, ZN => n5667);
   U6433 : INV_X1 port map( A => n5667, ZN => n5643);
   U6434 : INV_X2 port map( A => n7412, ZN => n7414);
   U6435 : AOI21_X1 port map( B1 => n7414, B2 => n7538, A => intadd_0xCI, ZN =>
                           n6091);
   U6436 : INV_X1 port map( A => n6091, ZN => n5642);
   U6437 : AOI21_X1 port map( B1 => n7454, B2 => IF_ISAxsection_0_port, A => 
                           n7112, ZN => n5646);
   U6438 : NAND3_X1 port map( A1 => n5641, A2 => n7453, A3 => n5646, ZN => 
                           n5668);
   U6439 : OAI22_X1 port map( A1 => n5643, A2 => n5642, B1 => n5668, B2 => 
                           intadd_4xSUMx0x, ZN => n5644);
   U6440 : AND2_X1 port map( A1 => IF_ISAxsection_0_port, A2 => 
                           fromMemoryPort_sync_port, ZN => n7451);
   U6441 : NAND2_X1 port map( A1 => n5645, A2 => n7451, ZN => n7522);
   U6442 : NAND2_X1 port map( A1 => n5644, A2 => n7522, ZN => n5649);
   U6443 : NAND2_X1 port map( A1 => IF_ISAxsection_0_port, A2 => n5645, ZN => 
                           n6070);
   U6444 : NOR2_X1 port map( A1 => rst, A2 => n6070, ZN => n6629);
   U6445 : NAND2_X1 port map( A1 => fromMemoryPort_sync_port, A2 => n6629, ZN 
                           => n7527);
   U6446 : OAI211_X1 port map( C1 => n5647, C2 => n7453, A => n5646, B => n7527
                           , ZN => n5666);
   U6447 : NAND2_X1 port map( A1 => n5666, A2 => IF_ISAxN2460, ZN => n5648);
   U6448 : AOI21_X1 port map( B1 => n5649, B2 => n5648, A => rst, ZN => 
                           IF_ISAxN10904);
   U6449 : NAND2_X1 port map( A1 => n5650, A2 => fromMemoryPortxLOADEDDATAx(31)
                           , ZN => n5651);
   U6450 : NAND2_X1 port map( A1 => n5652, A2 => n5651, ZN => n7375);
   U6451 : INV_X1 port map( A => n7375, ZN => n7388);
   U6452 : AOI22_X1 port map( A1 => n7375, A2 => n7544, B1 => 
                           IF_ISAxpcReg_signal_31_port, B2 => n7388, ZN => 
                           n5653);
   U6453 : XNOR2_X1 port map( A => intadd_0xn1, B => n5653, ZN => n5963);
   U6454 : NAND2_X1 port map( A1 => n5654, A2 => IF_ISAxpcReg_signal_30_port, 
                           ZN => n5655);
   U6455 : XOR2_X1 port map( A => IF_ISAxpcReg_signal_31_port, B => n5655, Z =>
                           n5967);
   U6456 : INV_X1 port map( A => n5967, ZN => n7434);
   U6457 : AOI22_X1 port map( A1 => n5656, A2 => n5963, B1 => n7434, B2 => 
                           n5764, ZN => n5966);
   U6458 : INV_X1 port map( A => n5963, ZN => n7379);
   U6459 : AOI22_X1 port map( A1 => n5767, A2 => n5967, B1 => n7379, B2 => 
                           n5657, ZN => n5961);
   U6460 : AOI22_X1 port map( A1 => n7434, A2 => n5659, B1 => n5961, B2 => 
                           n5658, ZN => n5664);
   U6461 : NAND2_X1 port map( A1 => n7431, A2 => n7375, ZN => n6036);
   U6462 : OAI21_X1 port map( B1 => n7431, B2 => n7375, A => n6036, ZN => n5660
                           );
   U6463 : XNOR2_X1 port map( A => n5660, B => intadd_3xn1, ZN => n5970);
   U6464 : AOI22_X1 port map( A1 => n5963, A2 => n5662, B1 => n5970, B2 => 
                           n5661, ZN => n5663);
   U6465 : OAI211_X1 port map( C1 => n5966, C2 => n5665, A => n5664, B => n5663
                           , ZN => n7553);
   U6466 : OAI21_X1 port map( B1 => n5667, B2 => n5666, A => IF_ISAxN2459, ZN 
                           => n5672);
   U6467 : NAND2_X1 port map( A1 => n7410, A2 => ashr_25xAx0x, ZN => n6150);
   U6468 : INV_X2 port map( A => n7123, ZN => n7410);
   U6469 : NOR2_X1 port map( A1 => ashr_25xAx0x, A2 => n7410, ZN => n5994);
   U6470 : INV_X1 port map( A => n5994, ZN => n5987);
   U6471 : AOI21_X1 port map( B1 => n6150, B2 => n5987, A => n5668, ZN => n5669
                           );
   U6472 : INV_X1 port map( A => n5669, ZN => n5671);
   U6473 : NOR2_X1 port map( A1 => n7522, A2 => IF_ISAxN2459, ZN => n5670);
   U6474 : AOI211_X1 port map( C1 => n5672, C2 => n5671, A => rst, B => n5670, 
                           ZN => n7548);
   U6475 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => intadd_3xAx2x, ZN 
                           => DP_OP_719J1_125_1055xn164);
   U6476 : AOI21_X1 port map( B1 => n5673, B2 => n5674, A => intadd_3xAx1x, ZN 
                           => DP_OP_719J1_125_1055xn163);
   U6477 : AOI21_X1 port map( B1 => n5675, B2 => n7360, A => intadd_3xAx0x, ZN 
                           => DP_OP_719J1_125_1055xn162);
   U6478 : AOI21_X1 port map( B1 => n5675, B2 => n5674, A => n7180, ZN => 
                           DP_OP_719J1_125_1055xn161);
   U6479 : AOI21_X1 port map( B1 => n5675, B2 => n5674, A => n7162, ZN => 
                           DP_OP_719J1_125_1055xn160);
   U6480 : AOI21_X1 port map( B1 => n5675, B2 => n7360, A => n7122, ZN => 
                           DP_OP_719J1_125_1055xn159);
   U6481 : AOI21_X1 port map( B1 => n5675, B2 => n5674, A => intadd_1xAx7x, ZN 
                           => DP_OP_719J1_125_1055xn158);
   U6482 : AOI21_X1 port map( B1 => n5675, B2 => n7360, A => intadd_1xAx6x, ZN 
                           => DP_OP_719J1_125_1055xn157);
   U6483 : AOI21_X1 port map( B1 => n5675, B2 => n7360, A => intadd_1xAx5x, ZN 
                           => DP_OP_719J1_125_1055xn156);
   U6484 : AOI21_X1 port map( B1 => n5675, B2 => n7360, A => intadd_1xAx4x, ZN 
                           => DP_OP_719J1_125_1055xn155);
   U6485 : AOI21_X1 port map( B1 => n5675, B2 => n5676, A => intadd_1xAx3x, ZN 
                           => DP_OP_719J1_125_1055xn154);
   U6486 : AOI21_X1 port map( B1 => n5678, B2 => n5676, A => intadd_1xAx2x, ZN 
                           => DP_OP_719J1_125_1055xn153);
   U6487 : AOI21_X1 port map( B1 => n5675, B2 => n5676, A => intadd_1xAx1x, ZN 
                           => DP_OP_719J1_125_1055xn152);
   U6488 : AOI21_X1 port map( B1 => n5678, B2 => n5677, A => intadd_1xAx0x, ZN 
                           => DP_OP_719J1_125_1055xn151);
   U6489 : AOI21_X1 port map( B1 => n5675, B2 => n5677, A => n6802, ZN => 
                           DP_OP_719J1_125_1055xn150);
   U6490 : AOI21_X1 port map( B1 => n5675, B2 => n5676, A => n6789, ZN => 
                           DP_OP_719J1_125_1055xn149);
   U6491 : AOI21_X1 port map( B1 => n5678, B2 => n5677, A => intadd_2xAx3x, ZN 
                           => DP_OP_719J1_125_1055xn148);
   U6492 : AOI21_X1 port map( B1 => n5678, B2 => n5676, A => intadd_2xAx2x, ZN 
                           => DP_OP_719J1_125_1055xn147);
   U6493 : AOI21_X1 port map( B1 => n5678, B2 => n5677, A => intadd_2xAx1x, ZN 
                           => DP_OP_719J1_125_1055xn146);
   U6494 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => intadd_2xAx0x, ZN 
                           => DP_OP_719J1_125_1055xn145);
   U6495 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => n6553, ZN => 
                           DP_OP_719J1_125_1055xn144);
   U6496 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => n6505, ZN => 
                           DP_OP_719J1_125_1055xn143);
   U6497 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => n6443, ZN => 
                           DP_OP_719J1_125_1055xn142);
   U6498 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => n6425, ZN => 
                           DP_OP_719J1_125_1055xn141);
   U6499 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => n6357, ZN => 
                           DP_OP_719J1_125_1055xn140);
   U6500 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => n5993, ZN => 
                           DP_OP_719J1_125_1055xn139);
   U6501 : INV_X1 port map( A => ashr_25xAx4x, ZN => n6276);
   U6502 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => n6276, ZN => 
                           DP_OP_719J1_125_1055xn138);
   U6503 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => intadd_4xAx2x, ZN 
                           => DP_OP_719J1_125_1055xn137);
   U6504 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => intadd_4xAx1x, ZN 
                           => DP_OP_719J1_125_1055xn136);
   U6505 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => intadd_4xAx0x, ZN 
                           => DP_OP_719J1_125_1055xn135);
   U6506 : INV_X1 port map( A => ashr_25xAx0x, ZN => n6049);
   U6507 : AOI21_X1 port map( B1 => n5678, B2 => n7360, A => n6049, ZN => 
                           DP_OP_719J1_125_1055xn134);
   U6508 : NOR2_X1 port map( A1 => n5679, A2 => n5691, ZN => n5681);
   U6509 : NOR2_X1 port map( A1 => n5681, A2 => n5680, ZN => n7172);
   U6510 : NOR2_X1 port map( A1 => n7372, A2 => n7036, ZN => n6390);
   U6511 : INV_X1 port map( A => n7082, ZN => n7164);
   U6512 : INV_X2 port map( A => n7296, ZN => n7205);
   U6513 : NAND2_X1 port map( A1 => n7205, A2 => n7409, ZN => n6243);
   U6514 : OAI22_X1 port map( A1 => n7161, A2 => ashr_25xAx29x, B1 => 
                           ashr_25xAx30x, B2 => n7205, ZN => n6218);
   U6515 : OR2_X1 port map( A1 => n7399, A2 => n6218, ZN => n5709);
   U6516 : OAI21_X1 port map( B1 => n7164, B2 => n6243, A => n5709, ZN => n6678
                           );
   U6517 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx21x, B1 => 
                           ashr_25xAx22x, B2 => n7395, ZN => n6220);
   U6518 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx23x, B1 => 
                           ashr_25xAx24x, B2 => n7161, ZN => n6223);
   U6519 : AOI22_X1 port map( A1 => n6144, A2 => n6220, B1 => n6223, B2 => 
                           n7082, ZN => n6475);
   U6520 : INV_X1 port map( A => n7399, ZN => n6586);
   U6521 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx25x, B1 => 
                           ashr_25xAx26x, B2 => n7395, ZN => n6222);
   U6522 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx27x, B1 => 
                           ashr_25xAx28x, B2 => n7296, ZN => n6219);
   U6523 : AOI22_X1 port map( A1 => n6586, A2 => n6222, B1 => n6219, B2 => 
                           n7082, ZN => n6107);
   U6524 : AOI22_X1 port map( A1 => n7305, A2 => n6475, B1 => n6107, B2 => 
                           n7303, ZN => n6672);
   U6525 : NOR2_X1 port map( A1 => n6672, A2 => n7203, ZN => n5711);
   U6526 : AOI21_X1 port map( B1 => n6390, B2 => n6678, A => n5711, ZN => n6334
                           );
   U6527 : NAND2_X1 port map( A1 => n5688, A2 => n6043, ZN => n5682);
   U6528 : NOR2_X1 port map( A1 => n5687, A2 => n5682, ZN => n6373);
   U6529 : AND2_X1 port map( A1 => n6373, A2 => n7081, ZN => n7013);
   U6530 : INV_X1 port map( A => n7013, ZN => n7423);
   U6531 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx5x, B1 => 
                           ashr_25xAx4x, B2 => n7296, ZN => n6402);
   U6532 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx3x, B1 => 
                           ashr_25xAx2x, B2 => n7161, ZN => n6202);
   U6533 : AOI22_X1 port map( A1 => n6586, A2 => n6402, B1 => n6202, B2 => 
                           n7082, ZN => n6487);
   U6534 : INV_X1 port map( A => n5683, ZN => n5988);
   U6535 : OAI21_X1 port map( B1 => n7161, B2 => ashr_25xAx1x, A => n5988, ZN 
                           => n6201);
   U6536 : NOR2_X1 port map( A1 => n7263, A2 => n6201, ZN => n6489);
   U6537 : AOI22_X1 port map( A1 => n7038, A2 => n6487, B1 => n6489, B2 => 
                           n7303, ZN => n6676);
   U6538 : NOR2_X1 port map( A1 => n5687, A2 => n5690, ZN => n5722);
   U6539 : NOR2_X1 port map( A1 => n7081, A2 => n5708, ZN => n5684);
   U6540 : AND2_X1 port map( A1 => n5722, A2 => n5684, ZN => n7344);
   U6541 : NAND2_X1 port map( A1 => n7372, A2 => n7344, ZN => n7043);
   U6542 : OAI22_X1 port map( A1 => n6334, A2 => n7423, B1 => n6676, B2 => 
                           n7043, ZN => n5733);
   U6543 : INV_X1 port map( A => intadd_0xBx0x, ZN => n6991);
   U6544 : AOI22_X1 port map( A1 => n7410, A2 => intadd_1xAx4x, B1 => 
                           intadd_1xAx5x, B2 => n7408, ZN => n6227);
   U6545 : CLKBUF_X1 port map( A => n7408, Z => n7123);
   U6546 : OAI22_X1 port map( A1 => n7123, A2 => intadd_1xAx6x, B1 => 
                           intadd_1xAx7x, B2 => n7410, ZN => n6230);
   U6547 : CLKBUF_X1 port map( A => n7254, Z => n7125);
   U6548 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6227, B1 => n6230, B2
                           => n7125, ZN => n6506);
   U6549 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx27x, B1 => 
                           ashr_25xAx28x, B2 => n7408, ZN => n6226);
   U6550 : OAI22_X1 port map( A1 => n7123, A2 => n7122, B1 => n7162, B2 => 
                           n7410, ZN => n6229);
   U6551 : INV_X1 port map( A => n6229, ZN => n5685);
   U6552 : MUX2_X1 port map( A => n6226, B => n5685, S => intadd_4xBx0x, Z => 
                           n6096);
   U6553 : AOI22_X1 port map( A1 => n6991, A2 => n6506, B1 => n6096, B2 => 
                           n7046, ZN => n6669);
   U6554 : NOR2_X1 port map( A1 => intadd_4xBx2x, A2 => n7046, ZN => n6416);
   U6555 : NOR2_X1 port map( A1 => n7123, A2 => n7431, ZN => n6231);
   U6556 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx29x, B1 => 
                           ashr_25xAx30x, B2 => n7408, ZN => n6225);
   U6557 : NOR2_X1 port map( A1 => n7254, A2 => n6225, ZN => n5689);
   U6558 : AOI21_X1 port map( B1 => n6231, B2 => n7254, A => n5689, ZN => n7280
                           );
   U6559 : INV_X1 port map( A => n7280, ZN => n5686);
   U6560 : AOI22_X1 port map( A1 => n7231, A2 => n6669, B1 => n6416, B2 => 
                           n5686, ZN => n6303);
   U6561 : NOR2_X1 port map( A1 => n5712, A2 => n5687, ZN => n5725);
   U6562 : NAND2_X1 port map( A1 => n5688, A2 => n5725, ZN => n6095);
   U6563 : NOR2_X1 port map( A1 => ashr_25xSHx4x, A2 => n6095, ZN => n7159);
   U6564 : INV_X1 port map( A => n7159, ZN => n7216);
   U6565 : NOR2_X1 port map( A1 => intadd_4xBx0x, A2 => n7431, ZN => n6370);
   U6566 : NOR2_X1 port map( A1 => n6370, A2 => n5689, ZN => n6072);
   U6567 : NAND2_X1 port map( A1 => n7409, A2 => n6337, ZN => n6253);
   U6568 : OAI21_X1 port map( B1 => n6072, B2 => n7046, A => n6253, ZN => n6666
                           );
   U6569 : AOI22_X1 port map( A1 => n7231, A2 => n6669, B1 => n6666, B2 => 
                           ashr_25xSHx3x, ZN => n6302);
   U6570 : NOR3_X1 port map( A1 => n5697, A2 => n5690, A3 => n5696, ZN => n5707
                           );
   U6571 : NAND2_X1 port map( A1 => n6045, A2 => n5707, ZN => n6073);
   U6572 : INV_X1 port map( A => n6073, ZN => n6254);
   U6573 : OAI21_X1 port map( B1 => n7327, B2 => n7409, A => n6254, ZN => n7325
                           );
   U6574 : AOI21_X1 port map( B1 => n7327, B2 => n6302, A => n7325, ZN => n5705
                           );
   U6575 : INV_X1 port map( A => intadd_0xSUMx19x, ZN => n5694);
   U6576 : NAND2_X1 port map( A1 => n5692, A2 => n5691, ZN => n7380);
   U6577 : NAND2_X1 port map( A1 => intadd_1xAx4x, A2 => add_x_26xBx21x, ZN => 
                           n5693);
   U6578 : NOR3_X1 port map( A1 => n5695, A2 => n5697, A3 => n5712, ZN => n7316
                           );
   U6579 : CLKBUF_X1 port map( A => n7316, Z => n7406);
   U6580 : INV_X1 port map( A => n7406, ZN => n7310);
   U6581 : OAI22_X1 port map( A1 => n5694, A2 => n7380, B1 => n5693, B2 => 
                           n7310, ZN => n5704);
   U6582 : NOR3_X1 port map( A1 => n5696, A2 => n5713, A3 => n5708, ZN => n5989
                           );
   U6583 : INV_X1 port map( A => n5989, ZN => n7394);
   U6584 : NOR3_X1 port map( A1 => n5697, A2 => n5696, A3 => n5695, ZN => n5698
                           );
   U6585 : AND2_X1 port map( A1 => n6043, A2 => n5698, ZN => n7323);
   U6586 : CLKBUF_X1 port map( A => n7323, Z => n7067);
   U6587 : INV_X1 port map( A => n7067, ZN => n7393);
   U6588 : AOI211_X1 port map( C1 => n7394, C2 => n7393, A => ashr_25xAx21x, B 
                           => n7473, ZN => n5703);
   U6589 : NOR2_X1 port map( A1 => n5700, A2 => n5699, ZN => n5701);
   U6590 : OAI22_X1 port map( A1 => intadd_1xBx4x, A2 => n7223, B1 => n7112, B2
                           => n5902, ZN => n5702);
   U6591 : NOR4_X1 port map( A1 => n5705, A2 => n5704, A3 => n5703, A4 => n5702
                           , ZN => n5731);
   U6592 : NOR2_X1 port map( A1 => ashr_25xSHx4x, A2 => n5712, ZN => n5706);
   U6593 : AND2_X1 port map( A1 => n5722, A2 => n5706, ZN => n7416);
   U6594 : AND2_X1 port map( A1 => n7416, A2 => ashr_25xSHx3x, ZN => n7427);
   U6595 : AOI22_X1 port map( A1 => n7329, A2 => intadd_2xAx2x, B1 => 
                           intadd_2xAx1x, B2 => n7408, ZN => n6758);
   U6596 : AOI22_X1 port map( A1 => n7329, A2 => intadd_2xAx0x, B1 => n6553, B2
                           => n7408, ZN => n6577);
   U6597 : AOI22_X1 port map( A1 => n7414, A2 => n6758, B1 => n6577, B2 => 
                           n7254, ZN => n6840);
   U6598 : AOI22_X1 port map( A1 => n7410, A2 => n6505, B1 => n6443, B2 => 
                           n7408, ZN => n6576);
   U6599 : AOI22_X1 port map( A1 => n7410, A2 => n6425, B1 => n6357, B2 => 
                           n7408, ZN => n6392);
   U6600 : AOI22_X1 port map( A1 => n7414, A2 => n6576, B1 => n6392, B2 => 
                           n7125, ZN => n6480);
   U6601 : AOI22_X1 port map( A1 => n6991, A2 => n6840, B1 => n6480, B2 => 
                           intadd_0xBx0x, ZN => n6680);
   U6602 : INV_X1 port map( A => n5707, ZN => n7381);
   U6603 : NOR2_X1 port map( A1 => n7381, A2 => n5708, ZN => n6404);
   U6604 : INV_X1 port map( A => n6404, ZN => n6313);
   U6605 : INV_X1 port map( A => n7349, ZN => n7079);
   U6606 : NAND2_X1 port map( A1 => n7409, A2 => n7399, ZN => n6709);
   U6607 : NAND2_X1 port map( A1 => n6709, A2 => n5709, ZN => n6684);
   U6608 : NOR2_X1 port map( A1 => n7431, A2 => n7372, ZN => n6492);
   U6609 : NAND2_X1 port map( A1 => n6492, A2 => n7036, ZN => n6377);
   U6610 : INV_X1 port map( A => n6377, ZN => n5710);
   U6611 : AOI211_X1 port map( C1 => n6390, C2 => n6684, A => n5711, B => n5710
                           , ZN => n6314);
   U6612 : INV_X1 port map( A => n7416, ZN => n7339);
   U6613 : NOR2_X1 port map( A1 => ashr_25xSHx3x, A2 => n7339, ZN => n7049);
   U6614 : AOI22_X1 port map( A1 => n7329, A2 => intadd_1xAx4x, B1 => 
                           intadd_1xAx3x, B2 => n7408, ZN => n7045);
   U6615 : AOI22_X1 port map( A1 => n7329, A2 => intadd_1xAx2x, B1 => 
                           intadd_1xAx1x, B2 => n7408, ZN => n6925);
   U6616 : AOI22_X1 port map( A1 => n7414, A2 => n7045, B1 => n6925, B2 => 
                           n7254, ZN => n7089);
   U6617 : AOI22_X1 port map( A1 => n7329, A2 => intadd_1xAx0x, B1 => n6802, B2
                           => n7408, ZN => n6924);
   U6618 : AOI22_X1 port map( A1 => n7329, A2 => n6789, B1 => intadd_2xAx3x, B2
                           => n7408, ZN => n6759);
   U6619 : AOI22_X1 port map( A1 => n7414, A2 => n6924, B1 => n6759, B2 => 
                           n7412, ZN => n6841);
   U6620 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n7089, B1 => n6841, B2
                           => n7046, ZN => n7258);
   U6621 : INV_X1 port map( A => n7315, ZN => n7382);
   U6622 : INV_X1 port map( A => n7406, ZN => n7250);
   U6623 : INV_X1 port map( A => n5713, ZN => n5714);
   U6624 : NAND2_X1 port map( A1 => n6043, A2 => n5714, ZN => n5715);
   U6625 : AOI221_X1 port map( B1 => n7323, B2 => n7473, C1 => n7248, C2 => 
                           n5717, A => n7246, ZN => n5718);
   U6626 : OAI221_X1 port map( B1 => intadd_1xBx4x, B2 => n7382, C1 => 
                           add_x_26xBx21x, C2 => n7250, A => n5718, ZN => n5719
                           );
   U6627 : AOI22_X1 port map( A1 => n7049, A2 => n7258, B1 => ashr_25xAx21x, B2
                           => n5719, ZN => n5720);
   U6628 : OAI221_X1 port map( B1 => n7079, B2 => n7081, C1 => n7079, C2 => 
                           n6314, A => n5720, ZN => n5729);
   U6629 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx13x, B1 => 
                           ashr_25xAx12x, B2 => n7395, ZN => n6764);
   U6630 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx11x, B1 => 
                           ashr_25xAx10x, B2 => n7395, ZN => n6585);
   U6631 : AOI22_X1 port map( A1 => n7164, A2 => n6764, B1 => n6585, B2 => 
                           n7263, ZN => n6850);
   U6632 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx9x, B1 => 
                           ashr_25xAx8x, B2 => n7395, ZN => n6584);
   U6633 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx7x, B1 => 
                           ashr_25xAx6x, B2 => n7296, ZN => n6403);
   U6634 : AOI22_X1 port map( A1 => n6586, A2 => n6584, B1 => n6403, B2 => 
                           n7082, ZN => n6488);
   U6635 : AOI22_X1 port map( A1 => n7305, A2 => n6850, B1 => n6488, B2 => 
                           n7303, ZN => n6677);
   U6636 : AND2_X1 port map( A1 => n6043, A2 => n7081, ZN => n5721);
   U6637 : AND2_X1 port map( A1 => n5722, A2 => n5721, ZN => n7405);
   U6638 : INV_X1 port map( A => n7405, ZN => n7202);
   U6639 : NOR2_X1 port map( A1 => n7372, A2 => n7202, ZN => n7390);
   U6640 : INV_X1 port map( A => n7390, ZN => n7308);
   U6641 : AND2_X1 port map( A1 => n7405, A2 => n7372, ZN => n7301);
   U6642 : AOI22_X1 port map( A1 => n7205, A2 => intadd_1xAx4x, B1 => 
                           intadd_1xAx3x, B2 => n7296, ZN => n7035);
   U6643 : AOI22_X1 port map( A1 => n7205, A2 => intadd_1xAx2x, B1 => 
                           intadd_1xAx1x, B2 => n7161, ZN => n6929);
   U6644 : AOI22_X1 port map( A1 => n7164, A2 => n7035, B1 => n6929, B2 => 
                           n7399, ZN => n7084);
   U6645 : AOI22_X1 port map( A1 => n7205, A2 => intadd_1xAx0x, B1 => n6802, B2
                           => n7296, ZN => n6928);
   U6646 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx15x, B1 => 
                           ashr_25xAx14x, B2 => n7395, ZN => n6765);
   U6647 : INV_X1 port map( A => n6765, ZN => n5723);
   U6648 : AOI22_X1 port map( A1 => n7164, A2 => n6928, B1 => n5723, B2 => 
                           n7399, ZN => n6849);
   U6649 : AOI22_X1 port map( A1 => n7305, A2 => n7084, B1 => n6849, B2 => 
                           n7036, ZN => n7265);
   U6650 : AND2_X1 port map( A1 => n5725, A2 => n5724, ZN => n5726);
   U6651 : AND2_X1 port map( A1 => n5726, A2 => ashr_25xSHx4x, ZN => n7348);
   U6652 : NAND2_X1 port map( A1 => n7231, A2 => n7348, ZN => n6958);
   U6653 : INV_X1 port map( A => n6958, ZN => n7039);
   U6654 : AOI22_X1 port map( A1 => n7410, A2 => n5993, B1 => n6276, B2 => 
                           n7408, ZN => n6391);
   U6655 : AOI22_X1 port map( A1 => n7410, A2 => intadd_4xAx2x, B1 => 
                           intadd_4xAx1x, B2 => n7408, ZN => n6185);
   U6656 : AOI22_X1 port map( A1 => n7414, A2 => n6391, B1 => n6185, B2 => 
                           n7125, ZN => n6479);
   U6657 : AOI21_X1 port map( B1 => n7410, B2 => intadd_4xAx0x, A => n5994, ZN 
                           => n6184);
   U6658 : NAND2_X1 port map( A1 => n7414, A2 => n6184, ZN => n6481);
   U6659 : AOI22_X1 port map( A1 => n6991, A2 => n6479, B1 => n6481, B2 => 
                           intadd_0xBx0x, ZN => n6679);
   U6660 : AOI22_X1 port map( A1 => n7301, A2 => n7265, B1 => n7039, B2 => 
                           n6679, ZN => n5727);
   U6661 : OAI21_X1 port map( B1 => n6677, B2 => n7308, A => n5727, ZN => n5728
                           );
   U6662 : AOI211_X1 port map( C1 => n7427, C2 => n6680, A => n5729, B => n5728
                           , ZN => n5730);
   U6663 : OAI211_X1 port map( C1 => n6303, C2 => n7216, A => n5731, B => n5730
                           , ZN => n5732);
   U6664 : AOI211_X1 port map( C1 => DP_OP_719J1_125_1055xn90, C2 => n7172, A 
                           => n5733, B => n5732, ZN => n5735);
   U6665 : NAND2_X1 port map( A1 => n7516, A2 => n6070, ZN => n6829);
   U6666 : INV_X1 port map( A => n6829, ZN => n7023);
   U6667 : INV_X1 port map( A => n7023, ZN => n7529);
   U6668 : INV_X1 port map( A => n6629, ZN => n7435);
   U6669 : OAI22_X1 port map( A1 => n5735, A2 => n7529, B1 => n7435, B2 => 
                           n5734, ZN => IF_ISAxN10958);
   U6670 : NAND2_X1 port map( A1 => n7372, A2 => n7036, ZN => n7402);
   U6671 : INV_X1 port map( A => n7402, ZN => n7269);
   U6672 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx20x, B1 => 
                           ashr_25xAx19x, B2 => n7161, ZN => n6992);
   U6673 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx18x, B1 => 
                           ashr_25xAx17x, B2 => n7395, ZN => n6881);
   U6674 : AOI22_X1 port map( A1 => n7164, A2 => n6992, B1 => n6881, B2 => 
                           n7263, ZN => n6969);
   U6675 : NAND2_X1 port map( A1 => n7038, A2 => n7372, ZN => n7262);
   U6676 : INV_X1 port map( A => n7262, ZN => n7397);
   U6677 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx24x, B1 => 
                           ashr_25xAx23x, B2 => n7395, ZN => n7136);
   U6678 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx22x, B1 => 
                           ashr_25xAx21x, B2 => n7161, ZN => n6993);
   U6679 : AOI22_X1 port map( A1 => n7164, A2 => n7136, B1 => n6993, B2 => 
                           n7399, ZN => n7209);
   U6680 : AOI22_X1 port map( A1 => n7269, A2 => n6969, B1 => n7397, B2 => 
                           n7209, ZN => n5738);
   U6681 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx8x, B1 => 
                           ashr_25xAx7x, B2 => n7408, ZN => n6527);
   U6682 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx6x, B1 => 
                           ashr_25xAx5x, B2 => n7408, ZN => n6352);
   U6683 : AOI22_X1 port map( A1 => n7414, A2 => n6527, B1 => n6352, B2 => 
                           n7254, ZN => n6638);
   U6684 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx2x, B1 => 
                           ashr_25xAx1x, B2 => n7408, ZN => n6151);
   U6685 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx4x, B1 => 
                           ashr_25xAx3x, B2 => n7408, ZN => n6351);
   U6686 : MUX2_X1 port map( A => n6151, B => n6351, S => intadd_4xBx0x, Z => 
                           n6275);
   U6687 : INV_X1 port map( A => n6275, ZN => n5736);
   U6688 : AOI22_X1 port map( A1 => n6991, A2 => n6638, B1 => n5736, B2 => 
                           intadd_0xBx0x, ZN => n6796);
   U6689 : OR2_X1 port map( A1 => n7254, A2 => n6150, ZN => n6274);
   U6690 : INV_X1 port map( A => n6416, ZN => n6581);
   U6691 : OAI22_X1 port map( A1 => n6796, A2 => ashr_25xSHx3x, B1 => n6274, B2
                           => n6581, ZN => n6442);
   U6692 : AOI22_X1 port map( A1 => n7410, A2 => intadd_1xAx7x, B1 => n7122, B2
                           => n7123, ZN => n6154);
   U6693 : AOI22_X1 port map( A1 => n7410, A2 => n7162, B1 => n7180, B2 => 
                           n7123, ZN => n6365);
   U6694 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6154, B1 => n6365, B2
                           => n7254, ZN => n6277);
   U6695 : AOI22_X1 port map( A1 => n7410, A2 => intadd_3xAx0x, B1 => 
                           intadd_3xAx1x, B2 => n7123, ZN => n6364);
   U6696 : AOI22_X1 port map( A1 => n7410, A2 => intadd_3xAx2x, B1 => n7431, B2
                           => n7123, ZN => n6156);
   U6697 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6364, B1 => n6156, B2
                           => n7125, ZN => n7240);
   U6698 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6277, B1 => n7240, B2
                           => n7046, ZN => n6054);
   U6699 : NAND2_X1 port map( A1 => n7231, A2 => n6054, ZN => n5746);
   U6700 : INV_X1 port map( A => n5746, ZN => n6440);
   U6701 : AOI22_X1 port map( A1 => n7348, A2 => n6442, B1 => n7159, B2 => 
                           n6440, ZN => n5737);
   U6702 : OAI21_X1 port map( B1 => n5738, B2 => n7202, A => n5737, ZN => n5757
                           );
   U6703 : NOR2_X1 port map( A1 => n7476, A2 => ashr_25xAx24x, ZN => n5739);
   U6704 : NOR2_X1 port map( A1 => intadd_1xBx7x, A2 => ashr_25xAx24x, ZN => 
                           n6023);
   U6705 : AOI22_X1 port map( A1 => n5739, A2 => n7067, B1 => n6023, B2 => 
                           n7406, ZN => n5755);
   U6706 : INV_X1 port map( A => n7380, ZN => n7270);
   U6707 : OAI22_X1 port map( A1 => intadd_1xBx7x, A2 => n7223, B1 => n7476, B2
                           => n7394, ZN => n5740);
   U6708 : AOI21_X1 port map( B1 => intadd_0xSUMx22x, B2 => n7270, A => n5740, 
                           ZN => n5754);
   U6709 : NOR2_X1 port map( A1 => intadd_4xBx1x, A2 => ashr_25xSHx3x, ZN => 
                           n7418);
   U6710 : INV_X1 port map( A => n7418, ZN => n7126);
   U6711 : AOI22_X1 port map( A1 => n7329, A2 => intadd_1xAx3x, B1 => 
                           intadd_1xAx2x, B2 => n7408, ZN => n6988);
   U6712 : AOI22_X1 port map( A1 => n7329, A2 => intadd_1xAx1x, B1 => 
                           intadd_1xAx0x, B2 => n7408, ZN => n6875);
   U6713 : AOI22_X1 port map( A1 => n7414, A2 => n6988, B1 => n6875, B2 => 
                           n7412, ZN => n6965);
   U6714 : NAND2_X1 port map( A1 => intadd_4xBx2x, A2 => intadd_4xBx1x, ZN => 
                           n7411);
   U6715 : OAI22_X1 port map( A1 => n7123, A2 => intadd_1xAx7x, B1 => 
                           intadd_1xAx6x, B2 => n7410, ZN => n7124);
   U6716 : AOI22_X1 port map( A1 => n7329, A2 => intadd_1xAx5x, B1 => 
                           intadd_1xAx4x, B2 => n7408, ZN => n6989);
   U6717 : AOI22_X1 port map( A1 => n7414, A2 => n7124, B1 => n6989, B2 => 
                           n7125, ZN => n7225);
   U6718 : AOI22_X1 port map( A1 => n7329, A2 => n6802, B1 => n6789, B2 => 
                           n7408, ZN => n6874);
   U6719 : AOI22_X1 port map( A1 => n7329, A2 => ashr_25xAx14x, B1 => 
                           ashr_25xAx13x, B2 => n7408, ZN => n6729);
   U6720 : INV_X1 port map( A => n6729, ZN => n5741);
   U6721 : AOI22_X1 port map( A1 => n7414, A2 => n6874, B1 => n5741, B2 => 
                           n7254, ZN => n6964);
   U6722 : INV_X1 port map( A => n6964, ZN => n5742);
   U6723 : AOI22_X1 port map( A1 => n7329, A2 => ashr_25xAx12x, B1 => 
                           ashr_25xAx11x, B2 => n7408, ZN => n6728);
   U6724 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx10x, B1 => 
                           ashr_25xAx9x, B2 => n7408, ZN => n6528);
   U6725 : AOI22_X1 port map( A1 => n7414, A2 => n6728, B1 => n6528, B2 => 
                           n7125, ZN => n6637);
   U6726 : AOI22_X1 port map( A1 => n6991, A2 => n5742, B1 => n6637, B2 => 
                           intadd_0xBx0x, ZN => n6799);
   U6727 : OAI222_X1 port map( A1 => n7126, A2 => n6965, B1 => n7411, B2 => 
                           n7225, C1 => n6799, C2 => intadd_4xBx2x, ZN => n5743
                           );
   U6728 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx8x, B1 => 
                           ashr_25xAx7x, B2 => n7161, ZN => n6539);
   U6729 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx6x, B1 => 
                           ashr_25xAx5x, B2 => n7296, ZN => n6336);
   U6730 : AOI22_X1 port map( A1 => n6586, A2 => n6539, B1 => n6336, B2 => 
                           n7399, ZN => n6631);
   U6731 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx4x, B1 => 
                           ashr_25xAx3x, B2 => n7161, ZN => n6335);
   U6732 : NOR2_X1 port map( A1 => intadd_4xAx0x, A2 => n7205, ZN => n6050);
   U6733 : AOI21_X1 port map( B1 => n7205, B2 => ashr_25xAx2x, A => n6050, ZN 
                           => n6174);
   U6734 : AOI22_X1 port map( A1 => n6586, A2 => n6335, B1 => n6174, B2 => 
                           n7399, ZN => n6256);
   U6735 : AOI22_X1 port map( A1 => n7038, A2 => n6631, B1 => n6256, B2 => 
                           n7303, ZN => n6798);
   U6736 : NAND3_X1 port map( A1 => n7164, A2 => n7205, A3 => ashr_25xAx0x, ZN 
                           => n6053);
   U6737 : INV_X1 port map( A => n6390, ZN => n6588);
   U6738 : OAI22_X1 port map( A1 => n6798, A2 => n7203, B1 => n6053, B2 => 
                           n6588, ZN => n6453);
   U6739 : AOI22_X1 port map( A1 => n7416, A2 => n5743, B1 => n7344, B2 => 
                           n6453, ZN => n5753);
   U6740 : AOI221_X1 port map( B1 => n7323, B2 => n7476, C1 => n7248, C2 => 
                           n5744, A => n7246, ZN => n5745);
   U6741 : OAI221_X1 port map( B1 => intadd_1xBx7x, B2 => n7382, C1 => 
                           add_x_26xBx24x, C2 => n7250, A => n5745, ZN => n5751
                           );
   U6742 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx24x, B1 => 
                           ashr_25xAx25x, B2 => n7161, ZN => n6136);
   U6743 : AOI22_X1 port map( A1 => n7396, A2 => ashr_25xAx26x, B1 => 
                           ashr_25xAx27x, B2 => n7395, ZN => n6132);
   U6744 : AOI22_X1 port map( A1 => n6144, A2 => n6136, B1 => n6132, B2 => 
                           n7399, ZN => n6252);
   U6745 : AOI22_X1 port map( A1 => n7396, A2 => ashr_25xAx28x, B1 => 
                           ashr_25xAx29x, B2 => n7395, ZN => n6131);
   U6746 : AOI22_X1 port map( A1 => n7396, A2 => ashr_25xAx30x, B1 => n7409, B2
                           => n7395, ZN => n6133);
   U6747 : AOI22_X1 port map( A1 => n6144, A2 => n6131, B1 => n6133, B2 => 
                           n7082, ZN => n6624);
   U6748 : AOI22_X1 port map( A1 => n7038, A2 => n6252, B1 => n6624, B2 => 
                           n7303, ZN => n6436);
   U6749 : INV_X1 port map( A => n6492, ZN => n6546);
   U6750 : OAI21_X1 port map( B1 => n6436, B2 => n7203, A => n6546, ZN => n6457
                           );
   U6751 : OAI21_X1 port map( B1 => n7345, B2 => n6457, A => n7349, ZN => n5748
                           );
   U6752 : NOR2_X1 port map( A1 => n7431, A2 => intadd_4xBx2x, ZN => n6665);
   U6753 : INV_X1 port map( A => n6665, ZN => n6708);
   U6754 : NAND2_X1 port map( A1 => n6708, A2 => n5746, ZN => n6441);
   U6755 : INV_X1 port map( A => n7325, ZN => n7130);
   U6756 : OAI21_X1 port map( B1 => ashr_25xSHx4x, B2 => n6441, A => n7130, ZN 
                           => n5747);
   U6757 : OAI211_X1 port map( C1 => n7112, C2 => n5918, A => n5748, B => n5747
                           , ZN => n5750);
   U6758 : NAND2_X1 port map( A1 => n7372, A2 => n7013, ZN => n7188);
   U6759 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx16x, B1 => 
                           ashr_25xAx15x, B2 => n7296, ZN => n6880);
   U6760 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx14x, B1 => 
                           ashr_25xAx13x, B2 => n7395, ZN => n6734);
   U6761 : AOI22_X1 port map( A1 => n7164, A2 => n6880, B1 => n6734, B2 => 
                           n7263, ZN => n6968);
   U6762 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx12x, B1 => 
                           ashr_25xAx11x, B2 => n7161, ZN => n6733);
   U6763 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx10x, B1 => 
                           ashr_25xAx9x, B2 => n7161, ZN => n6540);
   U6764 : AOI22_X1 port map( A1 => n7164, A2 => n6733, B1 => n6540, B2 => 
                           n7082, ZN => n6632);
   U6765 : AOI22_X1 port map( A1 => n7038, A2 => n6968, B1 => n6632, B2 => 
                           n7303, ZN => n6797);
   U6766 : OAI22_X1 port map( A1 => n6436, A2 => n7188, B1 => n6797, B2 => 
                           n7308, ZN => n5749);
   U6767 : AOI211_X1 port map( C1 => ashr_25xAx24x, C2 => n5751, A => n5750, B 
                           => n5749, ZN => n5752);
   U6768 : NAND4_X1 port map( A1 => n5755, A2 => n5754, A3 => n5753, A4 => 
                           n5752, ZN => n5756);
   U6769 : AOI211_X1 port map( C1 => DP_OP_719J1_125_1055xn93, C2 => n7172, A 
                           => n5757, B => n5756, ZN => n5759);
   U6770 : OAI22_X1 port map( A1 => n5759, A2 => n7529, B1 => n5758, B2 => 
                           n7435, ZN => IF_ISAxN10961);
   U6771 : NAND2_X1 port map( A1 => ashr_25xAx0x, A2 => n7123, ZN => 
                           intadd_4xCI);
   U6772 : OR4_X1 port map( A1 => IF_ISAxsection_2_port, A2 => n5770, A3 => 
                           n5769, A4 => n5760, ZN => n5808);
   U6773 : INV_X1 port map( A => n5808, ZN => n5964);
   U6774 : NOR4_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(2), A2 => n6388, 
                           A3 => n5770, A4 => n5761, ZN => n5763);
   U6775 : AND2_X1 port map( A1 => n5763, A2 => n5762, ZN => n5962);
   U6776 : INV_X1 port map( A => n5962, ZN => n5886);
   U6777 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(12), A2 => n5763
                           , ZN => n5951);
   U6778 : OAI22_X1 port map( A1 => n5767, A2 => n5886, B1 => n5951, B2 => 
                           n5764, ZN => n5773);
   U6779 : OAI211_X1 port map( C1 => n5765, C2 => n5951, A => n5776, B => n7531
                           , ZN => n5766);
   U6780 : AOI21_X1 port map( B1 => n5767, B2 => n5962, A => n5766, ZN => n5771
                           );
   U6781 : NOR3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(2), A2 => 
                           fromMemoryPortxLOADEDDATAx(4), A3 => n5768, ZN => 
                           n5960);
   U6782 : NOR4_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(3), A2 => 
                           IF_ISAxsection_2_port, A3 => n5770, A4 => n5769, ZN 
                           => n5775);
   U6783 : NOR2_X2 port map( A1 => n5960, A2 => n5775, ZN => n5953);
   U6784 : OAI22_X1 port map( A1 => n5771, A2 => n7538, B1 => intadd_4xSUMx0x, 
                           B2 => n5953, ZN => n5772);
   U6785 : AOI221_X1 port map( B1 => n5964, B2 => n6091, C1 => n5773, C2 => 
                           n6091, A => n5772, ZN => n5774);
   U6786 : NAND2_X1 port map( A1 => n7454, A2 => n7519, ZN => n5777);
   U6787 : OAI22_X1 port map( A1 => n5774, A2 => n5973, B1 => n7538, B2 => 
                           n5777, ZN => n7622);
   U6788 : NAND2_X1 port map( A1 => n5848, A2 => n5775, ZN => n5852);
   U6789 : NOR2_X1 port map( A1 => n5957, A2 => n5951, ZN => n5845);
   U6790 : AND2_X1 port map( A1 => n5776, A2 => n7531, ZN => n5778);
   U6791 : OAI21_X1 port map( B1 => n5957, B2 => n5778, A => n5777, ZN => n5843
                           );
   U6792 : AOI22_X1 port map( A1 => n5845, A2 => n5779, B1 => n7542, B2 => 
                           n5843, ZN => n5783);
   U6793 : INV_X1 port map( A => n5960, ZN => n5847);
   U6794 : OAI22_X1 port map( A1 => intadd_4xSUMx1x, A2 => n5847, B1 => n5886, 
                           B2 => n5780, ZN => n5781);
   U6795 : OAI221_X1 port map( B1 => n5781, B2 => n5964, C1 => n5781, C2 => 
                           intadd_0xSUMx0x, A => n5848, ZN => n5782);
   U6796 : OAI211_X1 port map( C1 => intadd_4xSUMx1x, C2 => n5852, A => n5783, 
                           B => n5782, ZN => n7621);
   U6797 : AOI22_X1 port map( A1 => n5785, A2 => n5845, B1 => n5784, B2 => 
                           n5843, ZN => n5789);
   U6798 : INV_X1 port map( A => n5962, ZN => n5950);
   U6799 : OAI22_X1 port map( A1 => intadd_4xSUMx2x, A2 => n5847, B1 => n5950, 
                           B2 => n5786, ZN => n5787);
   U6800 : OAI221_X1 port map( B1 => n5787, B2 => n5964, C1 => n5787, C2 => 
                           intadd_0xSUMx1x, A => n5848, ZN => n5788);
   U6801 : OAI211_X1 port map( C1 => intadd_4xSUMx2x, C2 => n5852, A => n5789, 
                           B => n5788, ZN => n7620);
   U6802 : AOI22_X1 port map( A1 => n5791, A2 => n5845, B1 => n5790, B2 => 
                           n5843, ZN => n5795);
   U6803 : OAI22_X1 port map( A1 => n5796, A2 => n5847, B1 => n5886, B2 => 
                           n5792, ZN => n5793);
   U6804 : OAI221_X1 port map( B1 => n5793, B2 => n5964, C1 => n5793, C2 => 
                           intadd_0xSUMx2x, A => n5848, ZN => n5794);
   U6805 : OAI211_X1 port map( C1 => n5796, C2 => n5852, A => n5795, B => n5794
                           , ZN => n7619);
   U6806 : INV_X1 port map( A => n5843, ZN => n5968);
   U6807 : INV_X1 port map( A => n5845, ZN => n5965);
   U6808 : INV_X1 port map( A => n5953, ZN => n5932);
   U6809 : AOI222_X1 port map( A1 => n5798, A2 => n5932, B1 => n5962, B2 => 
                           n5797, C1 => n5964, C2 => intadd_0xSUMx3x, ZN => 
                           n5799);
   U6810 : OAI222_X1 port map( A1 => n5801, A2 => n5968, B1 => n5965, B2 => 
                           n5800, C1 => n5973, C2 => n5799, ZN => n7618);
   U6811 : INV_X1 port map( A => n5852, ZN => n5971);
   U6812 : AOI22_X1 port map( A1 => n5803, A2 => n5971, B1 => n6362, B2 => 
                           n5843, ZN => n5806);
   U6813 : INV_X1 port map( A => intadd_0xSUMx4x, ZN => n6345);
   U6814 : OAI22_X1 port map( A1 => n5808, A2 => n6345, B1 => n5886, B2 => 
                           n5802, ZN => n5804);
   U6815 : OAI221_X1 port map( B1 => n5804, B2 => n5960, C1 => n5804, C2 => 
                           n5803, A => n5848, ZN => n5805);
   U6816 : OAI211_X1 port map( C1 => n5807, C2 => n5965, A => n5806, B => n5805
                           , ZN => n7617);
   U6817 : INV_X1 port map( A => n5808, ZN => n5956);
   U6818 : AOI22_X1 port map( A1 => n5956, A2 => intadd_0xSUMx5x, B1 => n5962, 
                           B2 => n5809, ZN => n5810);
   U6819 : OAI21_X1 port map( B1 => n5811, B2 => n5951, A => n5810, ZN => n5812
                           );
   U6820 : AOI21_X1 port map( B1 => n5813, B2 => n5932, A => n5812, ZN => n5814
                           );
   U6821 : OAI22_X1 port map( A1 => n5968, A2 => n6419, B1 => n5814, B2 => 
                           n5973, ZN => n7616);
   U6822 : AOI22_X1 port map( A1 => n5971, A2 => n5815, B1 => n6459, B2 => 
                           n5843, ZN => n5820);
   U6823 : INV_X1 port map( A => n5815, ZN => n5817);
   U6824 : OAI22_X1 port map( A1 => n5817, A2 => n5847, B1 => n5886, B2 => 
                           n5816, ZN => n5818);
   U6825 : OAI221_X1 port map( B1 => n5818, B2 => n5964, C1 => n5818, C2 => 
                           intadd_0xSUMx6x, A => n5848, ZN => n5819);
   U6826 : OAI211_X1 port map( C1 => n5821, C2 => n5965, A => n5820, B => n5819
                           , ZN => n7615);
   U6827 : NOR2_X1 port map( A1 => n5822, A2 => n5951, ZN => n5826);
   U6828 : OAI22_X1 port map( A1 => n5953, A2 => n5824, B1 => n5886, B2 => 
                           n5823, ZN => n5825);
   U6829 : AOI211_X1 port map( C1 => intadd_0xSUMx7x, C2 => n5956, A => n5826, 
                           B => n5825, ZN => n5827);
   U6830 : OAI22_X1 port map( A1 => n5968, A2 => n6495, B1 => n5827, B2 => 
                           n5973, ZN => n7614);
   U6831 : INV_X1 port map( A => n5829, ZN => n5828);
   U6832 : AOI22_X1 port map( A1 => n5828, A2 => n5971, B1 => n6532, B2 => 
                           n5843, ZN => n5833);
   U6833 : OAI22_X1 port map( A1 => n5950, A2 => n5830, B1 => n5847, B2 => 
                           n5829, ZN => n5831);
   U6834 : OAI221_X1 port map( B1 => n5831, B2 => n5964, C1 => n5831, C2 => 
                           intadd_0xSUMx8x, A => n5848, ZN => n5832);
   U6835 : OAI211_X1 port map( C1 => n5834, C2 => n5965, A => n5833, B => n5832
                           , ZN => n7613);
   U6836 : NAND2_X1 port map( A1 => n6553, A2 => n5835, ZN => n5836);
   U6837 : AOI21_X1 port map( B1 => n5837, B2 => n5836, A => n6565, ZN => 
                           intadd_2xCI);
   U6838 : NOR2_X1 port map( A1 => n5953, A2 => intadd_2xSUMx0x, ZN => n5841);
   U6839 : OAI22_X1 port map( A1 => n5839, A2 => n5951, B1 => n5886, B2 => 
                           n5838, ZN => n5840);
   U6840 : AOI211_X1 port map( C1 => intadd_0xSUMx9x, C2 => n5964, A => n5841, 
                           B => n5840, ZN => n5842);
   U6841 : OAI22_X1 port map( A1 => n5968, A2 => n6592, B1 => n5842, B2 => 
                           n5973, ZN => n7612);
   U6842 : AOI22_X1 port map( A1 => n5845, A2 => n5844, B1 => n6644, B2 => 
                           n5843, ZN => n5851);
   U6843 : OAI22_X1 port map( A1 => intadd_2xSUMx1x, A2 => n5847, B1 => n5886, 
                           B2 => n5846, ZN => n5849);
   U6844 : OAI221_X1 port map( B1 => n5849, B2 => n5964, C1 => n5849, C2 => 
                           intadd_0xSUMx10x, A => n5848, ZN => n5850);
   U6845 : OAI211_X1 port map( C1 => intadd_2xSUMx1x, C2 => n5852, A => n5851, 
                           B => n5850, ZN => n7611);
   U6846 : NOR2_X1 port map( A1 => n5950, A2 => n5853, ZN => n5856);
   U6847 : OAI22_X1 port map( A1 => n5953, A2 => intadd_2xSUMx2x, B1 => n5854, 
                           B2 => n5951, ZN => n5855);
   U6848 : AOI211_X1 port map( C1 => intadd_0xSUMx11x, C2 => n5956, A => n5856,
                           B => n5855, ZN => n5857);
   U6849 : OAI22_X1 port map( A1 => n5968, A2 => n5858, B1 => n5857, B2 => 
                           n5973, ZN => n7610);
   U6850 : OAI22_X1 port map( A1 => n5953, A2 => intadd_2xSUMx3x, B1 => n5886, 
                           B2 => n5859, ZN => n5860);
   U6851 : AOI21_X1 port map( B1 => n5964, B2 => intadd_0xSUMx12x, A => n5860, 
                           ZN => n5861);
   U6852 : OAI222_X1 port map( A1 => n6720, A2 => n5968, B1 => n5965, B2 => 
                           n5862, C1 => n5973, C2 => n5861, ZN => n7609);
   U6853 : AND2_X1 port map( A1 => n5932, A2 => n5863, ZN => n5867);
   U6854 : OAI22_X1 port map( A1 => n5865, A2 => n5951, B1 => n5886, B2 => 
                           n5864, ZN => n5866);
   U6855 : AOI211_X1 port map( C1 => n5964, C2 => intadd_0xSUMx13x, A => n5867,
                           B => n5866, ZN => n5868);
   U6856 : OAI22_X1 port map( A1 => n5968, A2 => n6777, B1 => n5868, B2 => 
                           n5973, ZN => n7608);
   U6857 : AND2_X1 port map( A1 => n5932, A2 => n5869, ZN => n5873);
   U6858 : OAI22_X1 port map( A1 => n5871, A2 => n5951, B1 => n5886, B2 => 
                           n5870, ZN => n5872);
   U6859 : AOI211_X1 port map( C1 => n5964, C2 => intadd_0xSUMx14x, A => n5873,
                           B => n5872, ZN => n5874);
   U6860 : OAI22_X1 port map( A1 => n5968, A2 => n5875, B1 => n5874, B2 => 
                           n5973, ZN => n7607);
   U6861 : AOI22_X1 port map( A1 => ashr_25xAx16x, A2 => add_x_26xBx16x, B1 => 
                           n6803, B2 => n5876, ZN => intadd_1xCI);
   U6862 : OAI22_X1 port map( A1 => n5953, A2 => intadd_1xSUMx0x, B1 => n5886, 
                           B2 => n5877, ZN => n5878);
   U6863 : AOI21_X1 port map( B1 => n5964, B2 => intadd_0xSUMx15x, A => n5878, 
                           ZN => n5879);
   U6864 : OAI222_X1 port map( A1 => n6834, A2 => n5968, B1 => n5965, B2 => 
                           n5880, C1 => n5973, C2 => n5879, ZN => n7606);
   U6865 : OAI22_X1 port map( A1 => n5953, A2 => intadd_1xSUMx1x, B1 => n5886, 
                           B2 => n5881, ZN => n5882);
   U6866 : AOI21_X1 port map( B1 => n5964, B2 => intadd_0xSUMx16x, A => n5882, 
                           ZN => n5883);
   U6867 : OAI222_X1 port map( A1 => n6889, A2 => n5968, B1 => n5965, B2 => 
                           n5884, C1 => n5973, C2 => n5883, ZN => n7605);
   U6868 : NOR2_X1 port map( A1 => n5953, A2 => intadd_1xSUMx2x, ZN => n5889);
   U6869 : OAI22_X1 port map( A1 => n5887, A2 => n5951, B1 => n5886, B2 => 
                           n5885, ZN => n5888);
   U6870 : AOI211_X1 port map( C1 => intadd_0xSUMx17x, C2 => n5956, A => n5889,
                           B => n5888, ZN => n5890);
   U6871 : OAI22_X1 port map( A1 => n5968, A2 => n6923, B1 => n5890, B2 => 
                           n5973, ZN => n7604);
   U6872 : NOR2_X1 port map( A1 => n5953, A2 => intadd_1xSUMx3x, ZN => n5894);
   U6873 : OAI22_X1 port map( A1 => n5892, A2 => n5951, B1 => n5950, B2 => 
                           n5891, ZN => n5893);
   U6874 : AOI211_X1 port map( C1 => intadd_0xSUMx18x, C2 => n5956, A => n5894,
                           B => n5893, ZN => n5895);
   U6875 : OAI22_X1 port map( A1 => n5968, A2 => n5896, B1 => n5895, B2 => 
                           n5957, ZN => n7603);
   U6876 : NOR2_X1 port map( A1 => n5950, A2 => n5897, ZN => n5900);
   U6877 : OAI22_X1 port map( A1 => n5953, A2 => intadd_1xSUMx4x, B1 => n5898, 
                           B2 => n5951, ZN => n5899);
   U6878 : AOI211_X1 port map( C1 => intadd_0xSUMx19x, C2 => n5956, A => n5900,
                           B => n5899, ZN => n5901);
   U6879 : OAI22_X1 port map( A1 => n5968, A2 => n5902, B1 => n5901, B2 => 
                           n5957, ZN => n7602);
   U6880 : NOR2_X1 port map( A1 => n5950, A2 => n5903, ZN => n5906);
   U6881 : OAI22_X1 port map( A1 => n5953, A2 => intadd_1xSUMx5x, B1 => n5904, 
                           B2 => n5951, ZN => n5905);
   U6882 : AOI211_X1 port map( C1 => intadd_0xSUMx20x, C2 => n5956, A => n5906,
                           B => n5905, ZN => n5907);
   U6883 : OAI22_X1 port map( A1 => n5968, A2 => n7014, B1 => n5907, B2 => 
                           n5957, ZN => n7601);
   U6884 : OAI22_X1 port map( A1 => n5953, A2 => intadd_1xSUMx6x, B1 => n5950, 
                           B2 => n5908, ZN => n5909);
   U6885 : AOI21_X1 port map( B1 => n5964, B2 => intadd_0xSUMx21x, A => n5909, 
                           ZN => n5910);
   U6886 : OAI222_X1 port map( A1 => n5912, A2 => n5968, B1 => n5965, B2 => 
                           n5911, C1 => n5973, C2 => n5910, ZN => n7600);
   U6887 : NOR2_X1 port map( A1 => n5950, A2 => n5913, ZN => n5916);
   U6888 : OAI22_X1 port map( A1 => n5953, A2 => intadd_1xSUMx7x, B1 => n5914, 
                           B2 => n5951, ZN => n5915);
   U6889 : AOI211_X1 port map( C1 => intadd_0xSUMx22x, C2 => n5956, A => n5916,
                           B => n5915, ZN => n5917);
   U6890 : OAI22_X1 port map( A1 => n5968, A2 => n5918, B1 => n5917, B2 => 
                           n5957, ZN => n7599);
   U6891 : NOR2_X1 port map( A1 => n5950, A2 => n5919, ZN => n5923);
   U6892 : OAI22_X1 port map( A1 => n5953, A2 => n5921, B1 => n5920, B2 => 
                           n5951, ZN => n5922);
   U6893 : AOI211_X1 port map( C1 => intadd_0xSUMx23x, C2 => n5956, A => n5923,
                           B => n5922, ZN => n5924);
   U6894 : OAI22_X1 port map( A1 => n5968, A2 => n7073, B1 => n5924, B2 => 
                           n5957, ZN => n7598);
   U6895 : NOR2_X1 port map( A1 => n5950, A2 => n5925, ZN => n5929);
   U6896 : OAI22_X1 port map( A1 => n5953, A2 => n5927, B1 => n5926, B2 => 
                           n5951, ZN => n5928);
   U6897 : AOI211_X1 port map( C1 => intadd_0xSUMx24x, C2 => n5956, A => n5929,
                           B => n5928, ZN => n5930);
   U6898 : OAI22_X1 port map( A1 => n5968, A2 => n7111, B1 => n5930, B2 => 
                           n5957, ZN => n7597);
   U6899 : AOI222_X1 port map( A1 => n5933, A2 => n5932, B1 => n5962, B2 => 
                           n5931, C1 => n5964, C2 => intadd_0xSUMx25x, ZN => 
                           n5934);
   U6900 : OAI222_X1 port map( A1 => n5936, A2 => n5968, B1 => n5965, B2 => 
                           n5935, C1 => n5957, C2 => n5934, ZN => n7596);
   U6901 : OAI22_X1 port map( A1 => n7178, A2 => n5937, B1 => ashr_25xAx27x, B2
                           => add_x_26xBx27x, ZN => intadd_3xCI);
   U6902 : NOR2_X1 port map( A1 => n5950, A2 => n5938, ZN => n5941);
   U6903 : OAI22_X1 port map( A1 => n5953, A2 => intadd_3xSUMx0x, B1 => n5939, 
                           B2 => n5951, ZN => n5940);
   U6904 : AOI211_X1 port map( C1 => intadd_0xSUMx26x, C2 => n5956, A => n5941,
                           B => n5940, ZN => n5942);
   U6905 : OAI22_X1 port map( A1 => n5968, A2 => n5943, B1 => n5942, B2 => 
                           n5957, ZN => n7595);
   U6906 : OAI22_X1 port map( A1 => n5953, A2 => intadd_3xSUMx1x, B1 => n5950, 
                           B2 => n5944, ZN => n5945);
   U6907 : AOI21_X1 port map( B1 => n5964, B2 => intadd_0xSUMx27x, A => n5945, 
                           ZN => n5946);
   U6908 : OAI222_X1 port map( A1 => n5948, A2 => n5968, B1 => n5965, B2 => 
                           n5947, C1 => n5973, C2 => n5946, ZN => n7594);
   U6909 : INV_X1 port map( A => n7357, ZN => n5959);
   U6910 : NOR2_X1 port map( A1 => n5950, A2 => n5949, ZN => n5955);
   U6911 : OAI22_X1 port map( A1 => n5953, A2 => intadd_3xSUMx2x, B1 => n5952, 
                           B2 => n5951, ZN => n5954);
   U6912 : AOI211_X1 port map( C1 => intadd_0xSUMx28x, C2 => n5956, A => n5955,
                           B => n5954, ZN => n5958);
   U6913 : OAI22_X1 port map( A1 => n5968, A2 => n5959, B1 => n5958, B2 => 
                           n5957, ZN => n7593);
   U6914 : AOI222_X1 port map( A1 => n5964, A2 => n5963, B1 => n5962, B2 => 
                           n5961, C1 => n5960, C2 => n5970, ZN => n5974);
   U6915 : OAI22_X1 port map( A1 => n5968, A2 => n5967, B1 => n5966, B2 => 
                           n5965, ZN => n5969);
   U6916 : AOI21_X1 port map( B1 => n5971, B2 => n5970, A => n5969, ZN => n5972
                           );
   U6917 : OAI21_X1 port map( B1 => n5974, B2 => n5973, A => n5972, ZN => n7592
                           );
   U6918 : NOR3_X1 port map( A1 => n5976, A2 => n5975, A3 => n5979, ZN => n7590
                           );
   U6919 : AOI211_X1 port map( C1 => fromMemoryPortxLOADEDDATAx(5), C2 => 
                           fromMemoryPortxLOADEDDATAx(14), A => n5979, B => 
                           fromMemoryPortxLOADEDDATAx(13), ZN => n5977);
   U6920 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(12), A2 => n5977,
                           ZN => n7589);
   U6921 : NOR2_X1 port map( A1 => n7534, A2 => n7531, ZN => n5978);
   U6922 : AOI21_X1 port map( B1 => n5978, B2 => n7516, A => n5977, ZN => n7588
                           );
   U6923 : INV_X1 port map( A => n5979, ZN => n5981);
   U6924 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(5), A2 => n5981,
                           ZN => n5980);
   U6925 : INV_X1 port map( A => n5980, ZN => n7591);
   U6926 : NOR2_X1 port map( A1 => n7396, A2 => n5980, ZN => n7587);
   U6927 : NOR2_X1 port map( A1 => n7081, A2 => n5980, ZN => n7586);
   U6928 : NOR2_X1 port map( A1 => n7038, A2 => n5980, ZN => n7585);
   U6929 : NOR2_X1 port map( A1 => n7372, A2 => n5980, ZN => n7584);
   U6930 : NOR2_X1 port map( A1 => n6144, A2 => n5980, ZN => n7583);
   U6931 : NOR2_X1 port map( A1 => rst, A2 => IF_ISAxsection_0_port, ZN => 
                           n7552);
   U6932 : INV_X1 port map( A => n7552, ZN => n7549);
   U6933 : NAND2_X1 port map( A1 => IF_ISAxsection_0_port, A2 => n5981, ZN => 
                           n5983);
   U6934 : OAI22_X1 port map( A1 => n7448, A2 => n5983, B1 => n5982, B2 => 
                           n7549, ZN => n7551);
   U6935 : INV_X1 port map( A => n7454, ZN => n5985);
   U6936 : OAI22_X1 port map( A1 => n5985, A2 => n7549, B1 => n5984, B2 => 
                           n5983, ZN => n7550);
   U6937 : INV_X1 port map( A => n7248, ZN => n7385);
   U6938 : INV_X1 port map( A => n7067, ZN => n7313);
   U6939 : OAI221_X1 port map( B1 => n7205, B2 => n7385, C1 => n7296, C2 => 
                           n7313, A => n7383, ZN => n5986);
   U6940 : AOI221_X1 port map( B1 => n7406, B2 => n7410, C1 => n7315, C2 => 
                           n7123, A => n5986, ZN => n6048);
   U6941 : OAI22_X1 port map( A1 => n5988, A2 => n7313, B1 => n5987, B2 => 
                           n7310, ZN => n5992);
   U6942 : CLKBUF_X1 port map( A => n5989, Z => n7318);
   U6943 : AOI22_X1 port map( A1 => n7246, A2 => n7123, B1 => n7318, B2 => 
                           n7296, ZN => n5990);
   U6944 : OAI211_X1 port map( C1 => n7112, C2 => n7545, A => n5990, B => n6070
                           , ZN => n5991);
   U6945 : AOI211_X1 port map( C1 => IF_ISAxN2459, C2 => n7270, A => n5992, B 
                           => n5991, ZN => n6047);
   U6946 : NOR2_X1 port map( A1 => intadd_3xBx1x, A2 => ashr_25xAx29x, ZN => 
                           n7252);
   U6947 : AOI22_X1 port map( A1 => n7180, A2 => add_x_26xBx27x, B1 => n7162, 
                           B2 => add_x_26xBx26x, ZN => n6031);
   U6948 : NOR2_X1 port map( A1 => n7076, A2 => ashr_25xAx25x, ZN => n7070);
   U6949 : OAI22_X1 port map( A1 => intadd_1xAx6x, A2 => add_x_26xBx23x, B1 => 
                           intadd_1xAx2x, B2 => add_x_26xBx19x, ZN => n6020);
   U6950 : NOR2_X1 port map( A1 => intadd_1xBx0x, A2 => ashr_25xAx17x, ZN => 
                           n6837);
   U6951 : NOR2_X1 port map( A1 => n6802, A2 => add_x_26xBx16x, ZN => n6015);
   U6952 : NAND2_X1 port map( A1 => n5993, A2 => add_x_26xBx5x, ZN => n6000);
   U6953 : NOR2_X1 port map( A1 => intadd_4xBx2x, A2 => ashr_25xAx3x, ZN => 
                           n6200);
   U6954 : NOR2_X1 port map( A1 => intadd_4xAx2x, A2 => ashr_25xSHx3x, ZN => 
                           n6199);
   U6955 : NOR2_X1 port map( A1 => intadd_4xBx1x, A2 => ashr_25xAx2x, ZN => 
                           n6161);
   U6956 : NAND2_X1 port map( A1 => ashr_25xAx1x, A2 => n7414, ZN => n6093);
   U6957 : AOI22_X1 port map( A1 => n7125, A2 => intadd_4xAx0x, B1 => n6093, B2
                           => n5994, ZN => n5995);
   U6958 : INV_X1 port map( A => n5995, ZN => n5996);
   U6959 : OAI22_X1 port map( A1 => n6161, A2 => n5996, B1 => intadd_4xAx1x, B2
                           => intadd_0xBx0x, ZN => n5997);
   U6960 : OAI22_X1 port map( A1 => n7327, A2 => ashr_25xAx4x, B1 => n6199, B2 
                           => n5997, ZN => n5998);
   U6961 : OAI22_X1 port map( A1 => n6200, A2 => n5998, B1 => n6276, B2 => 
                           ashr_25xSHx4x, ZN => n5999);
   U6962 : AOI22_X1 port map( A1 => ashr_25xAx5x, A2 => n6307, B1 => n6000, B2 
                           => n5999, ZN => n6001);
   U6963 : NAND2_X1 port map( A1 => ashr_25xAx6x, A2 => n6359, ZN => n6356);
   U6964 : AOI22_X1 port map( A1 => n6357, A2 => add_x_26xBx6x, B1 => n6001, B2
                           => n6356, ZN => n6003);
   U6965 : NAND2_X1 port map( A1 => n6425, A2 => add_x_26xBx7x, ZN => n6432);
   U6966 : OAI22_X1 port map( A1 => n6553, A2 => add_x_26xBx10x, B1 => n6505, 
                           B2 => add_x_26xBx9x, ZN => n6007);
   U6967 : OAI22_X1 port map( A1 => n6425, A2 => add_x_26xBx7x, B1 => n6443, B2
                           => add_x_26xBx8x, ZN => n6002);
   U6968 : AOI211_X1 port map( C1 => n6003, C2 => n6432, A => n6007, B => n6002
                           , ZN => n6013);
   U6969 : OAI22_X1 port map( A1 => n6789, A2 => add_x_26xBx15x, B1 => 
                           intadd_2xAx0x, B2 => add_x_26xBx11x, ZN => n6005);
   U6970 : OAI22_X1 port map( A1 => intadd_2xAx3x, A2 => add_x_26xBx14x, B1 => 
                           intadd_2xAx1x, B2 => add_x_26xBx12x, ZN => n6004);
   U6971 : AOI211_X1 port map( C1 => intadd_2xBx2x, C2 => ashr_25xAx13x, A => 
                           n6005, B => n6004, ZN => n6012);
   U6972 : AOI22_X1 port map( A1 => n6505, A2 => add_x_26xBx9x, B1 => n6443, B2
                           => add_x_26xBx8x, ZN => n6008);
   U6973 : AOI22_X1 port map( A1 => intadd_2xAx0x, A2 => add_x_26xBx11x, B1 => 
                           n6553, B2 => add_x_26xBx10x, ZN => n6006);
   U6974 : OAI21_X1 port map( B1 => n6008, B2 => n6007, A => n6006, ZN => n6011
                           );
   U6975 : NAND2_X1 port map( A1 => n6789, A2 => add_x_26xBx15x, ZN => n6009);
   U6976 : NAND2_X1 port map( A1 => intadd_2xAx3x, A2 => add_x_26xBx14x, ZN => 
                           n6722);
   U6977 : NAND2_X1 port map( A1 => intadd_2xAx2x, A2 => add_x_26xBx13x, ZN => 
                           n6682);
   U6978 : NAND2_X1 port map( A1 => intadd_2xAx1x, A2 => add_x_26xBx12x, ZN => 
                           n6642);
   U6979 : NAND4_X1 port map( A1 => n6009, A2 => n6722, A3 => n6682, A4 => 
                           n6642, ZN => n6010);
   U6980 : AOI221_X1 port map( B1 => n6013, B2 => n6012, C1 => n6011, C2 => 
                           n6012, A => n6010, ZN => n6014);
   U6981 : OAI22_X1 port map( A1 => n6811, A2 => ashr_25xAx16x, B1 => n6015, B2
                           => n6014, ZN => n6018);
   U6982 : AOI22_X1 port map( A1 => intadd_1xBx3x, A2 => ashr_25xAx20x, B1 => 
                           intadd_1xBx1x, B2 => ashr_25xAx18x, ZN => n6017);
   U6983 : AOI22_X1 port map( A1 => intadd_1xBx5x, A2 => ashr_25xAx22x, B1 => 
                           intadd_1xBx4x, B2 => ashr_25xAx21x, ZN => n6016);
   U6984 : OAI211_X1 port map( C1 => n6837, C2 => n6018, A => n6017, B => n6016
                           , ZN => n6019);
   U6985 : AOI211_X1 port map( C1 => intadd_1xBx0x, C2 => ashr_25xAx17x, A => 
                           n6020, B => n6019, ZN => n6024);
   U6986 : NOR2_X1 port map( A1 => intadd_1xBx6x, A2 => ashr_25xAx23x, ZN => 
                           n7030);
   U6987 : NOR2_X1 port map( A1 => intadd_1xBx3x, A2 => ashr_25xAx20x, ZN => 
                           n6947);
   U6988 : NOR2_X1 port map( A1 => intadd_1xBx2x, A2 => ashr_25xAx19x, ZN => 
                           n6915);
   U6989 : AOI211_X1 port map( C1 => intadd_1xAx1x, C2 => add_x_26xBx18x, A => 
                           n6947, B => n6915, ZN => n6021);
   U6990 : NAND2_X1 port map( A1 => intadd_1xAx5x, A2 => add_x_26xBx22x, ZN => 
                           n7005);
   U6991 : OAI211_X1 port map( C1 => intadd_1xBx4x, C2 => ashr_25xAx21x, A => 
                           n6021, B => n7005, ZN => n6022);
   U6992 : NOR4_X1 port map( A1 => n6024, A2 => n6023, A3 => n7030, A4 => n6022
                           , ZN => n6026);
   U6993 : AOI211_X1 port map( C1 => intadd_1xBx7x, C2 => ashr_25xAx24x, A => 
                           n6026, B => n6025, ZN => n6027);
   U6994 : OAI22_X1 port map( A1 => n7070, A2 => n6027, B1 => n7162, B2 => 
                           add_x_26xBx26x, ZN => n6030);
   U6995 : NOR2_X1 port map( A1 => n7180, A2 => add_x_26xBx27x, ZN => n6029);
   U6996 : OAI22_X1 port map( A1 => intadd_3xAx1x, A2 => add_x_26xBx29x, B1 => 
                           intadd_3xAx0x, B2 => add_x_26xBx28x, ZN => n6028);
   U6997 : AOI211_X1 port map( C1 => n6031, C2 => n6030, A => n6029, B => n6028
                           , ZN => n6032);
   U6998 : AOI211_X1 port map( C1 => intadd_3xAx0x, C2 => add_x_26xBx28x, A => 
                           n7252, B => n6032, ZN => n6033);
   U6999 : NAND2_X1 port map( A1 => intadd_3xAx2x, A2 => add_x_26xBx30x, ZN => 
                           n7311);
   U7000 : AOI22_X1 port map( A1 => n6033, A2 => n7311, B1 => intadd_3xBx2x, B2
                           => ashr_25xAx30x, ZN => n6037);
   U7001 : NAND2_X1 port map( A1 => n7409, A2 => n7388, ZN => n6034);
   U7002 : INV_X1 port map( A => n6036, ZN => n7407);
   U7003 : AOI21_X1 port map( B1 => n6037, B2 => n6034, A => n7407, ZN => n6041
                           );
   U7004 : INV_X1 port map( A => n6034, ZN => n6035);
   U7005 : AOI21_X1 port map( B1 => n6037, B2 => n6036, A => n6035, ZN => n6039
                           );
   U7006 : OAI22_X1 port map( A1 => n6041, A2 => n6040, B1 => n6039, B2 => 
                           n6038, ZN => n6044);
   U7007 : AOI22_X1 port map( A1 => n6045, A2 => n6044, B1 => n6043, B2 => 
                           n6042, ZN => n6046);
   U7008 : OAI211_X1 port map( C1 => n6049, C2 => n6048, A => n6047, B => n6046
                           , ZN => n6069);
   U7009 : CLKBUF_X1 port map( A => n7172, Z => n7364);
   U7010 : AOI22_X1 port map( A1 => n7396, A2 => ashr_25xAx4x, B1 => 
                           ashr_25xAx5x, B2 => n7296, ZN => n6145);
   U7011 : AOI22_X1 port map( A1 => n7396, A2 => ashr_25xAx6x, B1 => 
                           ashr_25xAx7x, B2 => n7296, ZN => n6139);
   U7012 : AOI22_X1 port map( A1 => n6144, A2 => n6145, B1 => n6139, B2 => 
                           n7082, ZN => n6264);
   U7013 : AOI22_X1 port map( A1 => n7396, A2 => intadd_4xAx1x, B1 => 
                           intadd_4xAx2x, B2 => n7395, ZN => n6147);
   U7014 : INV_X1 port map( A => n6053, ZN => n6255);
   U7015 : AOI221_X1 port map( B1 => n6050, B2 => n7164, C1 => n6147, C2 => 
                           n7399, A => n6255, ZN => n6051);
   U7016 : AOI22_X1 port map( A1 => n7396, A2 => ashr_25xAx8x, B1 => 
                           ashr_25xAx9x, B2 => n7296, ZN => n6138);
   U7017 : AOI22_X1 port map( A1 => n7396, A2 => ashr_25xAx10x, B1 => 
                           ashr_25xAx11x, B2 => n7395, ZN => n6141);
   U7018 : AOI22_X1 port map( A1 => n6144, A2 => n6138, B1 => n6141, B2 => 
                           n7082, ZN => n6265);
   U7019 : AOI22_X1 port map( A1 => n7396, A2 => ashr_25xAx12x, B1 => 
                           ashr_25xAx13x, B2 => n7161, ZN => n6140);
   U7020 : AOI22_X1 port map( A1 => n7396, A2 => ashr_25xAx14x, B1 => 
                           ashr_25xAx15x, B2 => n7161, ZN => n6143);
   U7021 : AOI22_X1 port map( A1 => n6144, A2 => n6140, B1 => n6143, B2 => 
                           n7082, ZN => n6263);
   U7022 : AOI22_X1 port map( A1 => n7038, A2 => n6265, B1 => n6263, B2 => 
                           n7303, ZN => n6438);
   U7023 : AOI22_X1 port map( A1 => n6051, A2 => n7397, B1 => n7203, B2 => 
                           n6438, ZN => n6052);
   U7024 : AND2_X1 port map( A1 => n6404, A2 => n7081, ZN => n6687);
   U7025 : INV_X1 port map( A => n6687, ZN => n6518);
   U7026 : NAND2_X1 port map( A1 => n7423, A2 => n6518, ZN => n6716);
   U7027 : OAI211_X1 port map( C1 => n7402, C2 => n6264, A => n6052, B => n6716
                           , ZN => n6065);
   U7028 : NOR3_X1 port map( A1 => n7254, A2 => n6150, A3 => n7411, ZN => n6816
                           );
   U7029 : NOR2_X1 port map( A1 => n7262, A2 => n6053, ZN => n6815);
   U7030 : AOI22_X1 port map( A1 => n7416, A2 => n6816, B1 => n7405, B2 => 
                           n6815, ZN => n6064);
   U7031 : INV_X1 port map( A => n6373, ZN => n6412);
   U7032 : NOR2_X1 port map( A1 => n7081, A2 => n6412, ZN => n6750);
   U7033 : AND2_X1 port map( A1 => n6404, A2 => n7345, ZN => n6711);
   U7034 : AOI22_X1 port map( A1 => n7396, A2 => ashr_25xAx16x, B1 => 
                           ashr_25xAx17x, B2 => n7395, ZN => n6142);
   U7035 : AOI22_X1 port map( A1 => n7396, A2 => ashr_25xAx18x, B1 => 
                           ashr_25xAx19x, B2 => n7161, ZN => n6135);
   U7036 : AOI22_X1 port map( A1 => n6144, A2 => n6142, B1 => n6135, B2 => 
                           n7263, ZN => n6262);
   U7037 : AOI22_X1 port map( A1 => n7396, A2 => ashr_25xAx20x, B1 => 
                           ashr_25xAx21x, B2 => n7161, ZN => n6134);
   U7038 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx22x, B1 => 
                           ashr_25xAx23x, B2 => n7395, ZN => n6137);
   U7039 : AOI22_X1 port map( A1 => n6144, A2 => n6134, B1 => n6137, B2 => 
                           n7263, ZN => n6251);
   U7040 : AOI22_X1 port map( A1 => n7305, A2 => n6262, B1 => n6251, B2 => 
                           n7303, ZN => n6437);
   U7041 : AOI22_X1 port map( A1 => n7372, A2 => n6437, B1 => n6436, B2 => 
                           n7203, ZN => n6814);
   U7042 : OAI21_X1 port map( B1 => n6750, B2 => n6711, A => n6814, ZN => n6063
                           );
   U7043 : NAND2_X1 port map( A1 => n6054, A2 => ashr_25xSHx3x, ZN => n6056);
   U7044 : AOI22_X1 port map( A1 => n7410, A2 => n6802, B1 => intadd_1xAx0x, B2
                           => n7123, ZN => n6123);
   U7045 : AOI22_X1 port map( A1 => n7410, A2 => intadd_1xAx1x, B1 => 
                           intadd_1xAx2x, B2 => n7123, ZN => n6153);
   U7046 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6123, B1 => n6153, B2
                           => n7125, ZN => n6267);
   U7047 : AOI22_X1 port map( A1 => n7410, A2 => intadd_1xAx3x, B1 => 
                           intadd_1xAx4x, B2 => n7123, ZN => n6152);
   U7048 : AOI22_X1 port map( A1 => n7410, A2 => intadd_1xAx5x, B1 => 
                           intadd_1xAx6x, B2 => n7123, ZN => n6155);
   U7049 : AOI22_X1 port map( A1 => n7414, A2 => n6152, B1 => n6155, B2 => 
                           n7125, ZN => n6278);
   U7050 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6267, B1 => n6278, B2
                           => n7046, ZN => n6446);
   U7051 : NAND2_X1 port map( A1 => n6446, A2 => intadd_4xBx2x, ZN => n6055);
   U7052 : AND2_X1 port map( A1 => n6056, A2 => n6055, ZN => n6817);
   U7053 : INV_X1 port map( A => n6817, ZN => n6061);
   U7054 : NAND2_X1 port map( A1 => n6095, A2 => n6073, ZN => n6083);
   U7055 : INV_X1 port map( A => n7411, ZN => n7337);
   U7056 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx2x, B1 => 
                           ashr_25xAx3x, B2 => n7123, ZN => n6125);
   U7057 : OAI22_X1 port map( A1 => n7410, A2 => n6093, B1 => n7414, B2 => 
                           n6125, ZN => n6057);
   U7058 : AOI22_X1 port map( A1 => n7410, A2 => n6443, B1 => n6505, B2 => 
                           n7408, ZN => n6119);
   U7059 : AOI22_X1 port map( A1 => n7410, A2 => n6553, B1 => intadd_2xAx0x, B2
                           => n7408, ZN => n6122);
   U7060 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6119, B1 => n6122, B2
                           => n7125, ZN => n6271);
   U7061 : AOI22_X1 port map( A1 => n7410, A2 => intadd_2xAx1x, B1 => 
                           intadd_2xAx2x, B2 => n7123, ZN => n6121);
   U7062 : AOI22_X1 port map( A1 => n7410, A2 => intadd_2xAx3x, B1 => n6789, B2
                           => n7123, ZN => n6124);
   U7063 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6121, B1 => n6124, B2
                           => n7254, ZN => n6268);
   U7064 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6271, B1 => n6268, B2
                           => n7046, ZN => n6448);
   U7065 : AOI22_X1 port map( A1 => n7337, A2 => n6057, B1 => n6448, B2 => 
                           ashr_25xSHx3x, ZN => n6059);
   U7066 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx4x, B1 => 
                           ashr_25xAx5x, B2 => n7123, ZN => n6126);
   U7067 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx6x, B1 => 
                           ashr_25xAx7x, B2 => n7123, ZN => n6118);
   U7068 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6126, B1 => n6118, B2
                           => n7254, ZN => n6269);
   U7069 : AOI211_X1 port map( C1 => n7418, C2 => n6269, A => n6816, B => 
                           ashr_25xSHx4x, ZN => n6058);
   U7070 : NAND2_X1 port map( A1 => n6059, A2 => n6058, ZN => n6060);
   U7071 : OAI211_X1 port map( C1 => n6061, C2 => n7327, A => n6083, B => n6060
                           , ZN => n6062);
   U7072 : NAND4_X1 port map( A1 => n6065, A2 => n6064, A3 => n6063, A4 => 
                           n6062, ZN => n6066);
   U7073 : AOI21_X1 port map( B1 => DP_OP_719J1_125_1055xn69, B2 => n7364, A =>
                           n6066, ZN => n6067);
   U7074 : INV_X1 port map( A => n6067, ZN => n6068);
   U7075 : OAI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(0), A2 => n6070,
                           B1 => n6069, B2 => n6068, ZN => n6071);
   U7076 : NOR2_X1 port map( A1 => rst, A2 => n6071, ZN => IF_ISAxN10936);
   U7077 : OAI22_X1 port map( A1 => n7164, A2 => n7385, B1 => n7414, B2 => 
                           n7382, ZN => n6106);
   U7078 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6096, B1 => n6072, B2
                           => n7046, ZN => n6483);
   U7079 : AOI22_X1 port map( A1 => n7410, A2 => intadd_1xAx0x, B1 => 
                           intadd_1xAx1x, B2 => n7408, ZN => n6192);
   U7080 : AOI22_X1 port map( A1 => n7410, A2 => intadd_1xAx2x, B1 => 
                           intadd_1xAx3x, B2 => n7408, ZN => n6228);
   U7081 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6192, B1 => n6228, B2
                           => n7254, ZN => n6507);
   U7082 : OAI221_X1 port map( B1 => intadd_4xBx1x, B2 => n6506, C1 => n7046, 
                           C2 => n6507, A => n7231, ZN => n6097);
   U7083 : OAI21_X1 port map( B1 => n6483, B2 => intadd_4xBx2x, A => n6097, ZN 
                           => n6855);
   U7084 : INV_X1 port map( A => n6855, ZN => n6080);
   U7085 : NOR2_X1 port map( A1 => n6073, A2 => n7327, ZN => n6769);
   U7086 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx9x, B1 => 
                           ashr_25xAx10x, B2 => n7161, ZN => n6207);
   U7087 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx11x, B1 => 
                           ashr_25xAx12x, B2 => n7296, ZN => n6204);
   U7088 : AOI22_X1 port map( A1 => n6144, A2 => n6207, B1 => n6204, B2 => 
                           n7263, ZN => n6312);
   U7089 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx13x, B1 => 
                           ashr_25xAx14x, B2 => n7161, ZN => n6203);
   U7090 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx15x, B1 => 
                           ashr_25xAx16x, B2 => n7395, ZN => n6206);
   U7091 : AOI22_X1 port map( A1 => n6144, A2 => n6203, B1 => n6206, B2 => 
                           n7082, ZN => n6309);
   U7092 : AOI22_X1 port map( A1 => n7305, A2 => n6312, B1 => n6309, B2 => 
                           n7303, ZN => n6477);
   U7093 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx5x, B1 => 
                           ashr_25xAx6x, B2 => n7161, ZN => n6210);
   U7094 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx7x, B1 => 
                           ashr_25xAx8x, B2 => n7395, ZN => n6208);
   U7095 : AOI22_X1 port map( A1 => n6144, A2 => n6210, B1 => n6208, B2 => 
                           n7082, ZN => n6308);
   U7096 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx3x, B1 => 
                           ashr_25xAx4x, B2 => n7296, ZN => n6209);
   U7097 : INV_X1 port map( A => n6209, ZN => n6077);
   U7098 : NOR2_X1 port map( A1 => ashr_25xAx1x, A2 => n7161, ZN => n6075);
   U7099 : NOR2_X1 port map( A1 => n7396, A2 => ashr_25xAx2x, ZN => n6074);
   U7100 : NOR2_X1 port map( A1 => n6075, A2 => n6074, ZN => n6076);
   U7101 : MUX2_X1 port map( A => n6077, B => n6076, S => n7164, Z => n6078);
   U7102 : OAI22_X1 port map( A1 => n7402, A2 => n6308, B1 => n7262, B2 => 
                           n6078, ZN => n6079);
   U7103 : AOI211_X1 port map( C1 => n6477, C2 => n7203, A => n7345, B => n6079
                           , ZN => n6109);
   U7104 : AOI222_X1 port map( A1 => DP_OP_719J1_125_1055xn70, A2 => n7364, B1 
                           => n6080, B2 => n6769, C1 => n6404, C2 => n6109, ZN 
                           => n6081);
   U7105 : INV_X1 port map( A => n6081, ZN => n6105);
   U7106 : AOI22_X1 port map( A1 => n7410, A2 => intadd_4xAx0x, B1 => 
                           intadd_4xAx1x, B2 => n7408, ZN => n6082);
   U7107 : AOI22_X1 port map( A1 => n7410, A2 => intadd_4xAx2x, B1 => n6276, B2
                           => n7408, ZN => n6189);
   U7108 : AOI221_X1 port map( B1 => n6082, B2 => n7414, C1 => n6189, C2 => 
                           n7412, A => n7411, ZN => n6086);
   U7109 : NAND2_X1 port map( A1 => n7327, A2 => n6083, ZN => n6754);
   U7110 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx9x, B1 => 
                           ashr_25xAx10x, B2 => n7408, ZN => n6194);
   U7111 : INV_X1 port map( A => n6194, ZN => n6084);
   U7112 : AOI22_X1 port map( A1 => n7410, A2 => intadd_2xAx0x, B1 => 
                           intadd_2xAx1x, B2 => n7408, ZN => n6191);
   U7113 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6084, B1 => n6191, B2
                           => n7125, ZN => n6301);
   U7114 : AOI22_X1 port map( A1 => n7410, A2 => intadd_2xAx2x, B1 => 
                           intadd_2xAx3x, B2 => n7408, ZN => n6190);
   U7115 : AOI22_X1 port map( A1 => n7410, A2 => n6789, B1 => n6802, B2 => 
                           n7408, ZN => n6193);
   U7116 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6190, B1 => n6193, B2
                           => n7125, ZN => n6298);
   U7117 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6301, B1 => n6298, B2
                           => n7046, ZN => n6508);
   U7118 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx5x, B1 => 
                           ashr_25xAx6x, B2 => n7408, ZN => n6187);
   U7119 : AOI22_X1 port map( A1 => n7410, A2 => ashr_25xAx7x, B1 => 
                           ashr_25xAx8x, B2 => n7408, ZN => n6195);
   U7120 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6187, B1 => n6195, B2
                           => n7254, ZN => n6299);
   U7121 : OAI22_X1 port map( A1 => n7231, A2 => n6508, B1 => n6299, B2 => 
                           n7126, ZN => n6085);
   U7122 : NOR3_X1 port map( A1 => n6086, A2 => n6754, A3 => n6085, ZN => n6088
                           );
   U7123 : OAI22_X1 port map( A1 => n7414, A2 => n7383, B1 => n7112, B2 => 
                           n7538, ZN => n6087);
   U7124 : AOI211_X1 port map( C1 => n7323, C2 => n6089, A => n6088, B => n6087
                           , ZN => n6103);
   U7125 : AOI22_X1 port map( A1 => n7305, A2 => n6107, B1 => n6684, B2 => 
                           n7303, ZN => n6491);
   U7126 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx17x, B1 => 
                           ashr_25xAx18x, B2 => n7395, ZN => n6205);
   U7127 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx19x, B1 => 
                           ashr_25xAx20x, B2 => n7395, ZN => n6221);
   U7128 : AOI22_X1 port map( A1 => n6144, A2 => n6205, B1 => n6221, B2 => 
                           n7399, ZN => n6476);
   U7129 : AOI221_X1 port map( B1 => n6600, B2 => n6476, C1 => n7036, C2 => 
                           n6475, A => n7203, ZN => n6108);
   U7130 : AOI21_X1 port map( B1 => n7203, B2 => n6491, A => n6108, ZN => n6843
                           );
   U7131 : NAND2_X1 port map( A1 => intadd_4xAx0x, A2 => n7125, ZN => n6094);
   U7132 : AOI22_X1 port map( A1 => n6091, A2 => n7270, B1 => n6090, B2 => 
                           n7323, ZN => n6092);
   U7133 : OAI221_X1 port map( B1 => n7310, B2 => n6094, C1 => n7250, C2 => 
                           n6093, A => n6092, ZN => n6101);
   U7134 : NOR2_X1 port map( A1 => n7327, A2 => n6095, ZN => n6630);
   U7135 : INV_X1 port map( A => n6630, ZN => n6485);
   U7136 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6096, B1 => n7280, B2
                           => n7046, ZN => n6484);
   U7137 : OAI21_X1 port map( B1 => n7231, B2 => n6484, A => n6097, ZN => n6847
                           );
   U7138 : NOR2_X1 port map( A1 => n7411, A2 => n6481, ZN => n6856);
   U7139 : NAND2_X1 port map( A1 => n7397, A2 => n6489, ZN => n6848);
   U7140 : INV_X1 port map( A => n6848, ZN => n6098);
   U7141 : AOI22_X1 port map( A1 => n7416, A2 => n6856, B1 => n7405, B2 => 
                           n6098, ZN => n6099);
   U7142 : OAI21_X1 port map( B1 => n6485, B2 => n6847, A => n6099, ZN => n6100
                           );
   U7143 : AOI211_X1 port map( C1 => n6711, C2 => n6843, A => n6101, B => n6100
                           , ZN => n6102);
   U7144 : OAI211_X1 port map( C1 => n6586, C2 => n7394, A => n6103, B => n6102
                           , ZN => n6104);
   U7145 : AOI211_X1 port map( C1 => ashr_25xAx1x, C2 => n6106, A => n6105, B 
                           => n6104, ZN => n6112);
   U7146 : NOR2_X1 port map( A1 => n7383, A2 => n7529, ZN => n6572);
   U7147 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(1), A2 => n6629,
                           B1 => n6572, B2 => ashr_25xAx1x, ZN => n6111);
   U7148 : NAND2_X1 port map( A1 => n6750, A2 => n7023, ZN => n6664);
   U7149 : INV_X1 port map( A => n6664, ZN => n6474);
   U7150 : AOI22_X1 port map( A1 => n6600, A2 => n6107, B1 => n6678, B2 => 
                           n7303, ZN => n7074);
   U7151 : AOI21_X1 port map( B1 => n7203, B2 => n7074, A => n6108, ZN => n6857
                           );
   U7152 : NOR2_X1 port map( A1 => n6412, A2 => n7529, ZN => n6330);
   U7153 : AOI22_X1 port map( A1 => n6474, A2 => n6857, B1 => n6330, B2 => 
                           n6109, ZN => n6110);
   U7154 : OAI211_X1 port map( C1 => n6112, C2 => n7529, A => n6111, B => n6110
                           , ZN => IF_ISAxN10938);
   U7155 : INV_X1 port map( A => n6113, ZN => n7443);
   U7156 : AOI22_X1 port map( A1 => n7246, A2 => n6337, B1 => n7443, B2 => 
                           n7542, ZN => n6116);
   U7157 : OAI22_X1 port map( A1 => intadd_4xBx1x, A2 => n7382, B1 => n7305, B2
                           => n7385, ZN => n6114);
   U7158 : OAI21_X1 port map( B1 => n7246, B2 => n6114, A => ashr_25xAx2x, ZN 
                           => n6115);
   U7159 : OAI211_X1 port map( C1 => n7380, C2 => n6117, A => n6116, B => n6115
                           , ZN => n6181);
   U7160 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn71, A2 => n7364, ZN 
                           => n6179);
   U7161 : INV_X1 port map( A => n6118, ZN => n6120);
   U7162 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6120, B1 => n6119, B2
                           => n7125, ZN => n6341);
   U7163 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6122, B1 => n6121, B2
                           => n7254, ZN => n6340);
   U7164 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6124, B1 => n6123, B2
                           => n7125, ZN => n6339);
   U7165 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6340, B1 => n6339, B2
                           => n7046, ZN => n6533);
   U7166 : OAI221_X1 port map( B1 => n7414, B2 => n6126, C1 => n7125, C2 => 
                           n6125, A => n7337, ZN => n6127);
   U7167 : OAI21_X1 port map( B1 => n7231, B2 => n6533, A => n6127, ZN => n6128
                           );
   U7168 : AOI211_X1 port map( C1 => n7418, C2 => n6341, A => n6754, B => n6128
                           , ZN => n6168);
   U7169 : NAND2_X1 port map( A1 => n7038, A2 => ashr_25xAx2x, ZN => n6130);
   U7170 : AOI21_X1 port map( B1 => n6130, B2 => n6129, A => n7393, ZN => n6167
                           );
   U7171 : AOI22_X1 port map( A1 => n6144, A2 => n6132, B1 => n6131, B2 => 
                           n7399, ZN => n6714);
   U7172 : NOR2_X1 port map( A1 => n7036, A2 => n6714, ZN => n6170);
   U7173 : NOR2_X1 port map( A1 => n7263, A2 => n6133, ZN => n6705);
   U7174 : NOR2_X1 port map( A1 => n7038, A2 => n6705, ZN => n6171);
   U7175 : NOR2_X1 port map( A1 => n6170, A2 => n6171, ZN => n6524);
   U7176 : AOI22_X1 port map( A1 => n6586, A2 => n6135, B1 => n6134, B2 => 
                           n7399, ZN => n6346);
   U7177 : AOI22_X1 port map( A1 => n6586, A2 => n6137, B1 => n6136, B2 => 
                           n7399, ZN => n6715);
   U7178 : AOI22_X1 port map( A1 => n6600, A2 => n6346, B1 => n6715, B2 => 
                           n7303, ZN => n6550);
   U7179 : NOR2_X1 port map( A1 => n6550, A2 => n7203, ZN => n6172);
   U7180 : AOI21_X1 port map( B1 => n6524, B2 => n7203, A => n6172, ZN => n6888
                           );
   U7181 : INV_X1 port map( A => n6750, ZN => n6763);
   U7182 : AOI22_X1 port map( A1 => n6144, A2 => n6139, B1 => n6138, B2 => 
                           n7082, ZN => n6348);
   U7183 : AOI22_X1 port map( A1 => n6144, A2 => n6141, B1 => n6140, B2 => 
                           n7399, ZN => n6349);
   U7184 : AOI22_X1 port map( A1 => n6144, A2 => n6143, B1 => n6142, B2 => 
                           n7399, ZN => n6347);
   U7185 : AOI22_X1 port map( A1 => n6600, A2 => n6349, B1 => n6347, B2 => 
                           n7303, ZN => n6548);
   U7186 : INV_X1 port map( A => n6145, ZN => n6146);
   U7187 : AOI221_X1 port map( B1 => n6147, B2 => n7164, C1 => n6146, C2 => 
                           n7082, A => n7262, ZN => n6148);
   U7188 : AOI211_X1 port map( C1 => n7203, C2 => n6548, A => n6148, B => n7345
                           , ZN => n6149);
   U7189 : OAI21_X1 port map( B1 => n7402, B2 => n6348, A => n6149, ZN => n6169
                           );
   U7190 : OAI22_X1 port map( A1 => n6888, A2 => n6763, B1 => n6313, B2 => 
                           n6169, ZN => n6166);
   U7191 : AOI22_X1 port map( A1 => intadd_4xBx0x, A2 => n6151, B1 => n6150, B2
                           => n7125, ZN => n6526);
   U7192 : NAND2_X1 port map( A1 => n7337, A2 => n6526, ZN => n6887);
   U7193 : AOI22_X1 port map( A1 => n7414, A2 => n6153, B1 => n6152, B2 => 
                           n7254, ZN => n6338);
   U7194 : AOI22_X1 port map( A1 => n7414, A2 => n6155, B1 => n6154, B2 => 
                           n7125, ZN => n6367);
   U7195 : AOI22_X1 port map( A1 => n6991, A2 => n6338, B1 => n6367, B2 => 
                           n7046, ZN => n6534);
   U7196 : NOR2_X1 port map( A1 => n6534, A2 => ashr_25xSHx3x, ZN => n6159);
   U7197 : NAND2_X1 port map( A1 => n7414, A2 => n6156, ZN => n6746);
   U7198 : AOI221_X1 port map( B1 => n6365, B2 => n7414, C1 => n6364, C2 => 
                           n7412, A => n6337, ZN => n6157);
   U7199 : AOI21_X1 port map( B1 => n7046, B2 => n6746, A => n6157, ZN => n6543
                           );
   U7200 : NOR2_X1 port map( A1 => intadd_4xBx2x, A2 => n6543, ZN => n6160);
   U7201 : NOR2_X1 port map( A1 => n6159, A2 => n6160, ZN => n6871);
   U7202 : INV_X1 port map( A => n6157, ZN => n6158);
   U7203 : NAND2_X1 port map( A1 => n6370, A2 => n6158, ZN => n6551);
   U7204 : AOI21_X1 port map( B1 => n6160, B2 => n6551, A => n6159, ZN => n6893
                           );
   U7205 : OAI221_X1 port map( B1 => n6769, B2 => n6871, C1 => n6769, C2 => 
                           n6630, A => n6893, ZN => n6164);
   U7206 : NOR2_X1 port map( A1 => intadd_4xAx1x, A2 => intadd_0xBx0x, ZN => 
                           n6162);
   U7207 : OAI21_X1 port map( B1 => n6162, B2 => n6161, A => n7316, ZN => n6163
                           );
   U7208 : OAI211_X1 port map( C1 => n7339, C2 => n6887, A => n6164, B => n6163
                           , ZN => n6165);
   U7209 : NOR4_X1 port map( A1 => n6168, A2 => n6167, A3 => n6166, A4 => n6165
                           , ZN => n6178);
   U7210 : INV_X1 port map( A => n6169, ZN => n6176);
   U7211 : AOI21_X1 port map( B1 => n6171, B2 => n6709, A => n6170, ZN => n6545
                           );
   U7212 : AOI21_X1 port map( B1 => n6545, B2 => n7203, A => n6172, ZN => n6869
                           );
   U7213 : INV_X1 port map( A => n6711, ZN => n6499);
   U7214 : NAND2_X1 port map( A1 => n7205, A2 => ashr_25xAx0x, ZN => n6173);
   U7215 : AOI22_X1 port map( A1 => n6586, A2 => n6174, B1 => n6173, B2 => 
                           n7082, ZN => n6538);
   U7216 : NAND2_X1 port map( A1 => n7397, A2 => n6538, ZN => n6873);
   U7217 : OAI22_X1 port map( A1 => n6869, A2 => n6499, B1 => n7202, B2 => 
                           n6873, ZN => n6175);
   U7218 : AOI21_X1 port map( B1 => n6373, B2 => n6176, A => n6175, ZN => n6177
                           );
   U7219 : NAND3_X1 port map( A1 => n6179, A2 => n6178, A3 => n6177, ZN => 
                           n6180);
   U7220 : AOI211_X1 port map( C1 => n7318, C2 => n7036, A => n6181, B => n6180
                           , ZN => n6183);
   U7221 : OAI22_X1 port map( A1 => n6183, A2 => n6829, B1 => n6182, B2 => 
                           n7435, ZN => IF_ISAxN10939);
   U7222 : NOR2_X1 port map( A1 => intadd_4xAx2x, A2 => n7203, ZN => n6242);
   U7223 : AOI22_X1 port map( A1 => n7414, A2 => n6185, B1 => n6184, B2 => 
                           n7125, ZN => n6582);
   U7224 : OR2_X1 port map( A1 => n7411, A2 => n6582, ZN => n6935);
   U7225 : OAI22_X1 port map( A1 => n6186, A2 => n7313, B1 => n7339, B2 => 
                           n6935, ZN => n6241);
   U7226 : INV_X1 port map( A => n6187, ZN => n6188);
   U7227 : AOI221_X1 port map( B1 => n6189, B2 => intadd_4xBx0x, C1 => n6188, 
                           C2 => n7412, A => n7411, ZN => n6197);
   U7228 : AOI22_X1 port map( A1 => n7414, A2 => n6191, B1 => n6190, B2 => 
                           n7254, ZN => n6397);
   U7229 : AOI22_X1 port map( A1 => n7414, A2 => n6193, B1 => n6192, B2 => 
                           n7125, ZN => n6394);
   U7230 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6397, B1 => n6394, B2
                           => intadd_0xBx0x, ZN => n6604);
   U7231 : AOI22_X1 port map( A1 => n7414, A2 => n6195, B1 => n6194, B2 => 
                           n7254, ZN => n6395);
   U7232 : OAI22_X1 port map( A1 => n7231, A2 => n6604, B1 => n6395, B2 => 
                           n7126, ZN => n6196);
   U7233 : NOR3_X1 port map( A1 => n6197, A2 => n6754, A3 => n6196, ZN => n6198
                           );
   U7234 : AOI221_X1 port map( B1 => n6200, B2 => n7406, C1 => n6199, C2 => 
                           n7406, A => n6198, ZN => n6238);
   U7235 : OAI22_X1 port map( A1 => intadd_4xBx2x, A2 => n7382, B1 => n7372, B2
                           => n7385, ZN => n6236);
   U7236 : AOI22_X1 port map( A1 => n6586, A2 => n6202, B1 => n6201, B2 => 
                           n7082, ZN => n6583);
   U7237 : NAND2_X1 port map( A1 => n7397, A2 => n6583, ZN => n6914);
   U7238 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn72, A2 => n7172, ZN 
                           => n6217);
   U7239 : AOI22_X1 port map( A1 => n6586, A2 => n6204, B1 => n6203, B2 => 
                           n7082, ZN => n6400);
   U7240 : AOI22_X1 port map( A1 => n6586, A2 => n6206, B1 => n6205, B2 => 
                           n7082, ZN => n6398);
   U7241 : AOI22_X1 port map( A1 => n7038, A2 => n6400, B1 => n6398, B2 => 
                           n7303, ZN => n6603);
   U7242 : AOI22_X1 port map( A1 => n6586, A2 => n6208, B1 => n6207, B2 => 
                           n7399, ZN => n6399);
   U7243 : OAI221_X1 port map( B1 => n7164, B2 => n6210, C1 => n7263, C2 => 
                           n6209, A => n7397, ZN => n6211);
   U7244 : OAI211_X1 port map( C1 => n7402, C2 => n6399, A => n7081, B => n6211
                           , ZN => n6212);
   U7245 : AOI21_X1 port map( B1 => n6603, B2 => n7203, A => n6212, ZN => n6247
                           );
   U7246 : OAI22_X1 port map( A1 => n7372, A2 => n7394, B1 => n7112, B2 => 
                           n6213, ZN => n6215);
   U7247 : NOR2_X1 port map( A1 => n7383, A2 => intadd_4xBx2x, ZN => n6214);
   U7248 : AOI211_X1 port map( C1 => n6404, C2 => n6247, A => n6215, B => n6214
                           , ZN => n6216);
   U7249 : OAI211_X1 port map( C1 => n6914, C2 => n7202, A => n6217, B => n6216
                           , ZN => n6235);
   U7250 : AOI22_X1 port map( A1 => n6586, A2 => n6219, B1 => n6218, B2 => 
                           n7399, ZN => n6593);
   U7251 : AOI21_X1 port map( B1 => n6600, B2 => n6593, A => n7372, ZN => n6246
                           );
   U7252 : AOI22_X1 port map( A1 => n6586, A2 => n6221, B1 => n6220, B2 => 
                           n7082, ZN => n6599);
   U7253 : AOI22_X1 port map( A1 => n6586, A2 => n6223, B1 => n6222, B2 => 
                           n7399, ZN => n6598);
   U7254 : AOI221_X1 port map( B1 => n6600, B2 => n6599, C1 => n7036, C2 => 
                           n6598, A => n7203, ZN => n6244);
   U7255 : AOI221_X1 port map( B1 => n6246, B2 => n7431, C1 => n6246, C2 => 
                           n7305, A => n6244, ZN => n6224);
   U7256 : INV_X1 port map( A => n6224, ZN => n6927);
   U7257 : AOI22_X1 port map( A1 => n7414, A2 => n6226, B1 => n6225, B2 => 
                           n7254, ZN => n6414);
   U7258 : INV_X1 port map( A => n6253, ZN => n6369);
   U7259 : AOI21_X1 port map( B1 => intadd_4xBx1x, B2 => n6414, A => n6369, ZN 
                           => n6573);
   U7260 : AOI22_X1 port map( A1 => n7414, A2 => n6228, B1 => n6227, B2 => 
                           n7125, ZN => n6393);
   U7261 : OAI22_X1 port map( A1 => n7125, A2 => n6230, B1 => n6229, B2 => 
                           n7414, ZN => n6413);
   U7262 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6393, B1 => n6413, B2
                           => n7046, ZN => n6606);
   U7263 : NOR2_X1 port map( A1 => n6606, A2 => ashr_25xSHx3x, ZN => n6232);
   U7264 : AOI21_X1 port map( B1 => n6573, B2 => ashr_25xSHx3x, A => n6232, ZN 
                           => n6911);
   U7265 : AND2_X1 port map( A1 => n7414, A2 => n6231, ZN => n7392);
   U7266 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6414, B1 => n7392, B2
                           => n7046, ZN => n6595);
   U7267 : AOI21_X1 port map( B1 => n6595, B2 => ashr_25xSHx3x, A => n6232, ZN 
                           => n6909);
   U7268 : AOI22_X1 port map( A1 => n6769, A2 => n6911, B1 => n6630, B2 => 
                           n6909, ZN => n6233);
   U7269 : OAI21_X1 port map( B1 => n6499, B2 => n6927, A => n6233, ZN => n6234
                           );
   U7270 : AOI211_X1 port map( C1 => ashr_25xAx3x, C2 => n6236, A => n6235, B 
                           => n6234, ZN => n6237);
   U7271 : OAI211_X1 port map( C1 => n6239, C2 => n7380, A => n6238, B => n6237
                           , ZN => n6240);
   U7272 : AOI211_X1 port map( C1 => n6242, C2 => n7323, A => n6241, B => n6240
                           , ZN => n6250);
   U7273 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(3), A2 => n6629,
                           B1 => n6572, B2 => ashr_25xAx3x, ZN => n6249);
   U7274 : NOR2_X1 port map( A1 => n7263, A2 => n6243, ZN => n6757);
   U7275 : NAND2_X1 port map( A1 => n6757, A2 => n7036, ZN => n6245);
   U7276 : AOI21_X1 port map( B1 => n6246, B2 => n6245, A => n6244, ZN => n6910
                           );
   U7277 : AOI22_X1 port map( A1 => n6474, A2 => n6910, B1 => n6330, B2 => 
                           n6247, ZN => n6248);
   U7278 : OAI211_X1 port map( C1 => n6250, C2 => n7529, A => n6249, B => n6248
                           , ZN => IF_ISAxN10940);
   U7279 : MUX2_X1 port map( A => n6252, B => n6251, S => n7038, Z => n6625);
   U7280 : AOI22_X1 port map( A1 => n6625, A2 => n7372, B1 => n6624, B2 => 
                           n6390, ZN => n6948);
   U7281 : NAND2_X1 port map( A1 => n6948, A2 => n6377, ZN => n6974);
   U7282 : OAI21_X1 port map( B1 => n7240, B2 => n7046, A => n6253, ZN => n6641
                           );
   U7283 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6278, B1 => n6277, B2
                           => n7046, ZN => n6655);
   U7284 : OAI221_X1 port map( B1 => n7231, B2 => n6641, C1 => ashr_25xSHx3x, 
                           C2 => n6655, A => n6254, ZN => n6966);
   U7285 : AOI21_X1 port map( B1 => n7383, B2 => n6966, A => n7327, ZN => n6293
                           );
   U7286 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn73, A2 => n7364, ZN 
                           => n6291);
   U7287 : AOI22_X1 port map( A1 => n6600, A2 => n6256, B1 => n6255, B2 => 
                           n7303, ZN => n6961);
   U7288 : INV_X1 port map( A => n6961, ZN => n6633);
   U7289 : OAI22_X1 port map( A1 => n7112, A2 => n6258, B1 => n7393, B2 => 
                           n6257, ZN => n6261);
   U7290 : OAI22_X1 port map( A1 => n6276, A2 => n7383, B1 => n7382, B2 => 
                           n6259, ZN => n6260);
   U7291 : AOI211_X1 port map( C1 => n7301, C2 => n6633, A => n6261, B => n6260
                           , ZN => n6290);
   U7292 : AOI22_X1 port map( A1 => n7305, A2 => n6263, B1 => n6262, B2 => 
                           n7303, ZN => n6627);
   U7293 : OAI22_X1 port map( A1 => n7402, A2 => n6265, B1 => n6264, B2 => 
                           n7262, ZN => n6266);
   U7294 : AOI21_X1 port map( B1 => n7203, B2 => n6627, A => n6266, ZN => n6273
                           );
   U7295 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6268, B1 => n6267, B2
                           => n7046, ZN => n6654);
   U7296 : OAI22_X1 port map( A1 => n7231, A2 => n6654, B1 => n6269, B2 => 
                           n7411, ZN => n6270);
   U7297 : AOI211_X1 port map( C1 => n6271, C2 => n7418, A => n6754, B => n6270
                           , ZN => n6272);
   U7298 : AOI21_X1 port map( B1 => n6273, B2 => n6716, A => n6272, ZN => n6289
                           );
   U7299 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6275, B1 => n6274, B2
                           => intadd_0xBx0x, ZN => n6639);
   U7300 : OAI221_X1 port map( B1 => n6276, B2 => n7385, C1 => ashr_25xAx4x, C2
                           => n7313, A => n7394, ZN => n6282);
   U7301 : NOR2_X1 port map( A1 => n7240, A2 => n6337, ZN => n6280);
   U7302 : AOI221_X1 port map( B1 => n6278, B2 => intadd_4xBx1x, C1 => n6277, 
                           C2 => intadd_0xBx0x, A => ashr_25xSHx3x, ZN => n6279
                           );
   U7303 : AOI21_X1 port map( B1 => n6280, B2 => ashr_25xSHx3x, A => n6279, ZN 
                           => n6949);
   U7304 : OAI22_X1 port map( A1 => n6948, A2 => n6763, B1 => n6949, B2 => 
                           n6485, ZN => n6281);
   U7305 : AOI21_X1 port map( B1 => n7345, B2 => n6282, A => n6281, ZN => n6283
                           );
   U7306 : INV_X1 port map( A => n6283, ZN => n6287);
   U7307 : OAI22_X1 port map( A1 => n6285, A2 => n7380, B1 => n6284, B2 => 
                           n7310, ZN => n6286);
   U7308 : AOI211_X1 port map( C1 => n6639, C2 => n7049, A => n6287, B => n6286
                           , ZN => n6288);
   U7309 : NAND4_X1 port map( A1 => n6291, A2 => n6290, A3 => n6289, A4 => 
                           n6288, ZN => n6292);
   U7310 : AOI211_X1 port map( C1 => n6711, C2 => n6974, A => n6293, B => n6292
                           , ZN => n6295);
   U7311 : OAI22_X1 port map( A1 => n6295, A2 => n6829, B1 => n6294, B2 => 
                           n7435, ZN => IF_ISAxN10941);
   U7312 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(5), A2 => n6629,
                           B1 => n6572, B2 => ashr_25xAx5x, ZN => n6333);
   U7313 : INV_X1 port map( A => n6676, ZN => n6297);
   U7314 : AOI22_X1 port map( A1 => n6297, A2 => n7301, B1 => n7406, B2 => 
                           n6296, ZN => n6326);
   U7315 : AOI22_X1 port map( A1 => n6991, A2 => n6298, B1 => n6507, B2 => 
                           intadd_0xBx0x, ZN => n6668);
   U7316 : OAI22_X1 port map( A1 => n7231, A2 => n6668, B1 => n6299, B2 => 
                           n7411, ZN => n6300);
   U7317 : AOI211_X1 port map( C1 => n7418, C2 => n6301, A => n6754, B => n6300
                           , ZN => n6324);
   U7318 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn74, A2 => n7172, ZN 
                           => n6322);
   U7319 : OAI22_X1 port map( A1 => n7457, A2 => n7394, B1 => n6307, B2 => 
                           n7383, ZN => n6305);
   U7320 : INV_X1 port map( A => n6769, ZN => n6967);
   U7321 : OAI22_X1 port map( A1 => n6303, A2 => n6485, B1 => n6302, B2 => 
                           n6967, ZN => n6304);
   U7322 : AOI211_X1 port map( C1 => n6306, C2 => n7443, A => n6305, B => n6304
                           , ZN => n6321);
   U7323 : OAI22_X1 port map( A1 => n7457, A2 => n7385, B1 => n7382, B2 => 
                           n6307, ZN => n6319);
   U7324 : INV_X1 port map( A => n6308, ZN => n6310);
   U7325 : AOI22_X1 port map( A1 => n6600, A2 => n6309, B1 => n6476, B2 => 
                           n7303, ZN => n6673);
   U7326 : AOI22_X1 port map( A1 => n6310, A2 => n7397, B1 => n7203, B2 => 
                           n6673, ZN => n6311);
   U7327 : OAI211_X1 port map( C1 => n6312, C2 => n7402, A => n7081, B => n6311
                           , ZN => n6328);
   U7328 : OAI22_X1 port map( A1 => n6314, A2 => n6499, B1 => n6313, B2 => 
                           n6328, ZN => n6318);
   U7329 : OAI22_X1 port map( A1 => n6316, A2 => n7313, B1 => n6315, B2 => 
                           n7380, ZN => n6317);
   U7330 : AOI211_X1 port map( C1 => ashr_25xAx5x, C2 => n6319, A => n6318, B 
                           => n6317, ZN => n6320);
   U7331 : NAND3_X1 port map( A1 => n6322, A2 => n6321, A3 => n6320, ZN => 
                           n6323);
   U7332 : AOI211_X1 port map( C1 => n7049, C2 => n6679, A => n6324, B => n6323
                           , ZN => n6325);
   U7333 : OAI211_X1 port map( C1 => n6327, C2 => n7313, A => n6326, B => n6325
                           , ZN => n6331);
   U7334 : INV_X1 port map( A => n6328, ZN => n6329);
   U7335 : AOI22_X1 port map( A1 => n7023, A2 => n6331, B1 => n6330, B2 => 
                           n6329, ZN => n6332);
   U7336 : OAI211_X1 port map( C1 => n6334, C2 => n6664, A => n6333, B => n6332
                           , ZN => IF_ISAxN10942);
   U7337 : AOI22_X1 port map( A1 => n6586, A2 => n6336, B1 => n6335, B2 => 
                           n7082, ZN => n6541);
   U7338 : AOI22_X1 port map( A1 => n7038, A2 => n6541, B1 => n6538, B2 => 
                           n7303, ZN => n7008);
   U7339 : INV_X1 port map( A => n7301, ZN => n6997);
   U7340 : AOI22_X1 port map( A1 => n6991, A2 => n6339, B1 => n6338, B2 => 
                           n6337, ZN => n6742);
   U7341 : AOI22_X1 port map( A1 => n7337, A2 => n6341, B1 => n7418, B2 => 
                           n6340, ZN => n6342);
   U7342 : OAI21_X1 port map( B1 => intadd_4xBx2x, B2 => n6742, A => n6342, ZN 
                           => n6343);
   U7343 : OAI22_X1 port map( A1 => n7008, A2 => n6997, B1 => n6754, B2 => 
                           n6343, ZN => n6387);
   U7344 : NAND2_X1 port map( A1 => n6357, A2 => add_x_26xBx6x, ZN => n6344);
   U7345 : OAI22_X1 port map( A1 => n6345, A2 => n7380, B1 => n6344, B2 => 
                           n7310, ZN => n6386);
   U7346 : AOI22_X1 port map( A1 => n7038, A2 => n6347, B1 => n6346, B2 => 
                           n7303, ZN => n6719);
   U7347 : OAI22_X1 port map( A1 => n7402, A2 => n6349, B1 => n7262, B2 => 
                           n6348, ZN => n6350);
   U7348 : AOI211_X1 port map( C1 => n6719, C2 => n7203, A => n7345, B => n6350
                           , ZN => n6372);
   U7349 : AOI22_X1 port map( A1 => n7414, A2 => n6352, B1 => n6351, B2 => 
                           n7254, ZN => n6529);
   U7350 : AOI22_X1 port map( A1 => n6991, A2 => n6529, B1 => n6526, B2 => 
                           n7046, ZN => n6731);
   U7351 : INV_X1 port map( A => n6731, ZN => n7011);
   U7352 : AOI22_X1 port map( A1 => n6404, A2 => n6372, B1 => n7049, B2 => 
                           n7011, ZN => n6355);
   U7353 : OAI221_X1 port map( B1 => n7458, B2 => n6357, C1 => n6353, C2 => 
                           ashr_25xAx6x, A => n7323, ZN => n6354);
   U7354 : OAI211_X1 port map( C1 => n7310, C2 => n6356, A => n6355, B => n6354
                           , ZN => n6385);
   U7355 : AOI221_X1 port map( B1 => n6357, B2 => n7394, C1 => n7385, C2 => 
                           n7394, A => n7458, ZN => n6361);
   U7356 : AOI21_X1 port map( B1 => n7315, B2 => ashr_25xAx6x, A => n7246, ZN 
                           => n6358);
   U7357 : OAI22_X1 port map( A1 => n6359, A2 => n6358, B1 => n6357, B2 => 
                           n7383, ZN => n6360);
   U7358 : AOI211_X1 port map( C1 => n6362, C2 => n7443, A => n6361, B => n6360
                           , ZN => n6381);
   U7359 : INV_X1 port map( A => n6705, ZN => n6363);
   U7360 : OAI221_X1 port map( B1 => n7305, B2 => n6714, C1 => n7303, C2 => 
                           n6715, A => n7372, ZN => n6376);
   U7361 : OAI21_X1 port map( B1 => n6588, B2 => n6363, A => n6376, ZN => n7012
                           );
   U7362 : INV_X1 port map( A => n6746, ZN => n7294);
   U7363 : NAND2_X1 port map( A1 => intadd_4xBx1x, A2 => n7294, ZN => n6368);
   U7364 : AOI22_X1 port map( A1 => n7414, A2 => n6365, B1 => n6364, B2 => 
                           n7125, ZN => n6366);
   U7365 : AOI22_X1 port map( A1 => n6991, A2 => n6367, B1 => n6366, B2 => 
                           intadd_0xBx0x, ZN => n6743);
   U7366 : NAND2_X1 port map( A1 => n7231, A2 => n6743, ZN => n6371);
   U7367 : OAI21_X1 port map( B1 => n7231, B2 => n6368, A => n6371, ZN => n6987
                           );
   U7368 : AOI22_X1 port map( A1 => n6750, A2 => n7012, B1 => n6630, B2 => 
                           n6987, ZN => n6380);
   U7369 : AOI211_X1 port map( C1 => n7294, C2 => intadd_4xBx1x, A => n6370, B 
                           => n6369, ZN => n6706);
   U7370 : OAI21_X1 port map( B1 => n7231, B2 => n6706, A => n6371, ZN => n7019
                           );
   U7371 : AOI22_X1 port map( A1 => n6373, A2 => n6372, B1 => n6769, B2 => 
                           n7019, ZN => n6379);
   U7372 : INV_X1 port map( A => n6709, ZN => n6374);
   U7373 : OAI21_X1 port map( B1 => n6705, B2 => n6374, A => n6390, ZN => n6375
                           );
   U7374 : NAND3_X1 port map( A1 => n6377, A2 => n6376, A3 => n6375, ZN => 
                           n6999);
   U7375 : NAND2_X1 port map( A1 => n6711, A2 => n6999, ZN => n6378);
   U7376 : NAND4_X1 port map( A1 => n6381, A2 => n6380, A3 => n6379, A4 => 
                           n6378, ZN => n6382);
   U7377 : AOI21_X1 port map( B1 => DP_OP_719J1_125_1055xn75, B2 => n7172, A =>
                           n6382, ZN => n6383);
   U7378 : INV_X1 port map( A => n6383, ZN => n6384);
   U7379 : NOR4_X1 port map( A1 => n6387, A2 => n6386, A3 => n6385, A4 => n6384
                           , ZN => n6389);
   U7380 : OAI22_X1 port map( A1 => n6389, A2 => n6829, B1 => n6388, B2 => 
                           n7435, ZN => IF_ISAxN10943);
   U7381 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(7), ZN => n7438);
   U7382 : AOI22_X1 port map( A1 => n7038, A2 => n6598, B1 => n6593, B2 => 
                           n7303, ZN => n6784);
   U7383 : NOR2_X1 port map( A1 => n6784, A2 => n7203, ZN => n6409);
   U7384 : AOI21_X1 port map( B1 => n6390, B2 => n6757, A => n6409, ZN => n7055
                           );
   U7385 : AOI22_X1 port map( A1 => n7414, A2 => n6392, B1 => n6391, B2 => 
                           n7125, ZN => n6579);
   U7386 : AOI22_X1 port map( A1 => n6991, A2 => n6579, B1 => n6582, B2 => 
                           intadd_0xBx0x, ZN => n7040);
   U7387 : AOI22_X1 port map( A1 => n6991, A2 => n6394, B1 => n6393, B2 => 
                           intadd_0xBx0x, ZN => n6753);
   U7388 : OAI22_X1 port map( A1 => n7231, A2 => n6753, B1 => n6395, B2 => 
                           n7411, ZN => n6396);
   U7389 : AOI211_X1 port map( C1 => n7418, C2 => n6397, A => n6754, B => n6396
                           , ZN => n6434);
   U7390 : AOI22_X1 port map( A1 => n7038, A2 => n6398, B1 => n6599, B2 => 
                           n7303, ZN => n6783);
   U7391 : OAI22_X1 port map( A1 => n7402, A2 => n6400, B1 => n7262, B2 => 
                           n6399, ZN => n6401);
   U7392 : AOI211_X1 port map( C1 => n7203, C2 => n6783, A => n7345, B => n6401
                           , ZN => n6410);
   U7393 : AOI22_X1 port map( A1 => n6586, A2 => n6403, B1 => n6402, B2 => 
                           n7263, ZN => n6587);
   U7394 : AOI22_X1 port map( A1 => n6600, A2 => n6587, B1 => n6583, B2 => 
                           n7303, ZN => n7044);
   U7395 : INV_X1 port map( A => n7044, ZN => n7368);
   U7396 : AOI22_X1 port map( A1 => n6404, A2 => n6410, B1 => n7368, B2 => 
                           n7301, ZN => n6431);
   U7397 : NOR2_X1 port map( A1 => n6425, A2 => n7313, ZN => n6408);
   U7398 : AOI221_X1 port map( B1 => n7323, B2 => n6425, C1 => n7248, C2 => 
                           ashr_25xAx7x, A => n7318, ZN => n6405);
   U7399 : INV_X1 port map( A => n6405, ZN => n6407);
   U7400 : MUX2_X1 port map( A => n6408, B => n6407, S => n6406, Z => n6429);
   U7401 : NOR2_X1 port map( A1 => n6492, A2 => n6409, ZN => n7051);
   U7402 : INV_X1 port map( A => n6410, ZN => n6411);
   U7403 : OAI22_X1 port map( A1 => n7051, A2 => n6499, B1 => n6412, B2 => 
                           n6411, ZN => n6428);
   U7404 : INV_X1 port map( A => n6413, ZN => n6415);
   U7405 : AOI22_X1 port map( A1 => n6991, A2 => n6415, B1 => n6414, B2 => 
                           intadd_0xBx0x, ZN => n6756);
   U7406 : NOR2_X1 port map( A1 => n6756, A2 => ashr_25xSHx3x, ZN => n6417);
   U7407 : AOI21_X1 port map( B1 => n7392, B2 => n6416, A => n6417, ZN => n7032
                           );
   U7408 : NOR2_X1 port map( A1 => n6665, A2 => n6417, ZN => n7056);
   U7409 : OAI22_X1 port map( A1 => n7032, A2 => n6485, B1 => n7056, B2 => 
                           n6967, ZN => n6427);
   U7410 : NOR2_X1 port map( A1 => n7310, A2 => add_x_26xBx7x, ZN => n6418);
   U7411 : AOI211_X1 port map( C1 => n7315, C2 => add_x_26xBx7x, A => n7246, B 
                           => n6418, ZN => n6424);
   U7412 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn76, A2 => n7364, ZN 
                           => n6423);
   U7413 : OAI22_X1 port map( A1 => n7383, A2 => n6420, B1 => n7112, B2 => 
                           n6419, ZN => n6421);
   U7414 : AOI21_X1 port map( B1 => intadd_0xSUMx5x, B2 => n7270, A => n6421, 
                           ZN => n6422);
   U7415 : OAI211_X1 port map( C1 => n6425, C2 => n6424, A => n6423, B => n6422
                           , ZN => n6426);
   U7416 : NOR4_X1 port map( A1 => n6429, A2 => n6428, A3 => n6427, A4 => n6426
                           , ZN => n6430);
   U7417 : OAI211_X1 port map( C1 => n6432, C2 => n7250, A => n6431, B => n6430
                           , ZN => n6433);
   U7418 : AOI211_X1 port map( C1 => n7049, C2 => n7040, A => n6434, B => n6433
                           , ZN => n6435);
   U7419 : OAI222_X1 port map( A1 => n7438, A2 => n7435, B1 => n6664, B2 => 
                           n7055, C1 => n7529, C2 => n6435, ZN => IF_ISAxN10944
                           );
   U7420 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(8), ZN => n7439);
   U7421 : NOR2_X1 port map( A1 => n6436, A2 => n7203, ZN => n6439);
   U7422 : NOR2_X1 port map( A1 => n7423, A2 => n7529, ZN => n6628);
   U7423 : AOI22_X1 port map( A1 => n7372, A2 => n6438, B1 => n6437, B2 => 
                           n7203, ZN => n6458);
   U7424 : AOI22_X1 port map( A1 => n6474, A2 => n6439, B1 => n6628, B2 => 
                           n6458, ZN => n6473);
   U7425 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn77, A2 => n7364, ZN 
                           => n6456);
   U7426 : AOI22_X1 port map( A1 => n6769, A2 => n6441, B1 => n6630, B2 => 
                           n6440, ZN => n6455);
   U7427 : INV_X1 port map( A => n6442, ZN => n6451);
   U7428 : OAI21_X1 port map( B1 => n6443, B2 => n7385, A => n7394, ZN => n6444
                           );
   U7429 : NAND2_X1 port map( A1 => n6445, A2 => n6444, ZN => n6450);
   U7430 : OR2_X1 port map( A1 => n6446, A2 => n7231, ZN => n6447);
   U7431 : INV_X1 port map( A => n6754, ZN => n6741);
   U7432 : OAI211_X1 port map( C1 => n6448, C2 => ashr_25xSHx3x, A => n6447, B 
                           => n6741, ZN => n6449);
   U7433 : OAI211_X1 port map( C1 => n7339, C2 => n6451, A => n6450, B => n6449
                           , ZN => n6452);
   U7434 : AOI21_X1 port map( B1 => n7405, B2 => n6453, A => n6452, ZN => n6454
                           );
   U7435 : NAND3_X1 port map( A1 => n6456, A2 => n6455, A3 => n6454, ZN => 
                           n6471);
   U7436 : AOI22_X1 port map( A1 => n6687, A2 => n6458, B1 => n6711, B2 => 
                           n6457, ZN => n6468);
   U7437 : INV_X1 port map( A => intadd_0xSUMx6x, ZN => n6463);
   U7438 : AOI22_X1 port map( A1 => n7315, A2 => n6460, B1 => n6459, B2 => 
                           n7443, ZN => n6462);
   U7439 : OAI21_X1 port map( B1 => add_x_26xBx8x, B2 => ashr_25xAx8x, A => 
                           n7246, ZN => n6461);
   U7440 : OAI211_X1 port map( C1 => n6463, C2 => n7380, A => n6462, B => n6461
                           , ZN => n6464);
   U7441 : AOI221_X1 port map( B1 => n6466, B2 => n7323, C1 => n6465, C2 => 
                           n7067, A => n6464, ZN => n6467);
   U7442 : OAI211_X1 port map( C1 => n6469, C2 => n7250, A => n6468, B => n6467
                           , ZN => n6470);
   U7443 : OAI21_X1 port map( B1 => n6471, B2 => n6470, A => n7023, ZN => n6472
                           );
   U7444 : OAI211_X1 port map( C1 => n7435, C2 => n7439, A => n6473, B => n6472
                           , ZN => IF_ISAxN10945);
   U7445 : NAND2_X1 port map( A1 => n7372, A2 => n6474, ZN => n6623);
   U7446 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(9), A2 => n6629,
                           B1 => n6572, B2 => ashr_25xAx9x, ZN => n6523);
   U7447 : AOI22_X1 port map( A1 => n7038, A2 => n6476, B1 => n6475, B2 => 
                           n7303, ZN => n6478);
   U7448 : MUX2_X1 port map( A => n6478, B => n6477, S => n7372, Z => n6519);
   U7449 : AOI22_X1 port map( A1 => n6991, A2 => n6480, B1 => n6479, B2 => 
                           n7046, ZN => n6842);
   U7450 : INV_X1 port map( A => n6842, ZN => n6482);
   U7451 : OAI22_X1 port map( A1 => n6482, A2 => ashr_25xSHx3x, B1 => n6481, B2
                           => n6581, ZN => n7085);
   U7452 : AOI21_X1 port map( B1 => n7231, B2 => n6483, A => n6665, ZN => n7092
                           );
   U7453 : NAND2_X1 port map( A1 => n7231, A2 => n6484, ZN => n7078);
   U7454 : OAI22_X1 port map( A1 => n7092, A2 => n6967, B1 => n6485, B2 => 
                           n7078, ZN => n6486);
   U7455 : AOI21_X1 port map( B1 => n7416, B2 => n7085, A => n6486, ZN => n6517
                           );
   U7456 : AOI22_X1 port map( A1 => n7038, A2 => n6488, B1 => n6487, B2 => 
                           n7303, ZN => n6846);
   U7457 : INV_X1 port map( A => n6489, ZN => n6490);
   U7458 : OAI22_X1 port map( A1 => n7203, A2 => n6846, B1 => n6490, B2 => 
                           n6588, ZN => n7090);
   U7459 : INV_X1 port map( A => n6491, ZN => n6493);
   U7460 : AOI21_X1 port map( B1 => n6493, B2 => n7372, A => n6492, ZN => n7080
                           );
   U7461 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn78, A2 => n7172, ZN 
                           => n6498);
   U7462 : NAND3_X1 port map( A1 => n6504, A2 => n7248, A3 => ashr_25xAx9x, ZN 
                           => n6494);
   U7463 : OAI21_X1 port map( B1 => n7112, B2 => n6495, A => n6494, ZN => n6496
                           );
   U7464 : AOI21_X1 port map( B1 => n7246, B2 => add_x_26xBx9x, A => n6496, ZN 
                           => n6497);
   U7465 : OAI211_X1 port map( C1 => n7080, C2 => n6499, A => n6498, B => n6497
                           , ZN => n6515);
   U7466 : NOR2_X1 port map( A1 => n6505, A2 => n6500, ZN => n6501);
   U7467 : AOI22_X1 port map( A1 => n6502, A2 => n7067, B1 => n6501, B2 => 
                           n7315, ZN => n6513);
   U7468 : AOI22_X1 port map( A1 => intadd_0xSUMx7x, A2 => n7270, B1 => n6503, 
                           B2 => n7316, ZN => n6512);
   U7469 : OAI211_X1 port map( C1 => n7318, C2 => n7323, A => n6505, B => n6504
                           , ZN => n6511);
   U7470 : AOI22_X1 port map( A1 => n6991, A2 => n6507, B1 => n6506, B2 => 
                           n7046, ZN => n6509);
   U7471 : OAI221_X1 port map( B1 => n7231, B2 => n6509, C1 => ashr_25xSHx3x, 
                           C2 => n6508, A => n6741, ZN => n6510);
   U7472 : NAND4_X1 port map( A1 => n6513, A2 => n6512, A3 => n6511, A4 => 
                           n6510, ZN => n6514);
   U7473 : AOI211_X1 port map( C1 => n7405, C2 => n7090, A => n6515, B => n6514
                           , ZN => n6516);
   U7474 : OAI211_X1 port map( C1 => n6519, C2 => n6518, A => n6517, B => n6516
                           , ZN => n6521);
   U7475 : INV_X1 port map( A => n6519, ZN => n6520);
   U7476 : AOI22_X1 port map( A1 => n7023, A2 => n6521, B1 => n6628, B2 => 
                           n6520, ZN => n6522);
   U7477 : OAI211_X1 port map( C1 => n7074, C2 => n6623, A => n6523, B => n6522
                           , ZN => IF_ISAxN10946);
   U7478 : INV_X1 port map( A => n6524, ZN => n7118);
   U7479 : INV_X1 port map( A => intadd_0xSUMx8x, ZN => n6568);
   U7480 : OAI21_X1 port map( B1 => n7462, B2 => ashr_25xAx10x, A => n6525, ZN 
                           => n6531);
   U7481 : INV_X1 port map( A => n6526, ZN => n6530);
   U7482 : AOI22_X1 port map( A1 => n7414, A2 => n6528, B1 => n6527, B2 => 
                           n7254, ZN => n6730);
   U7483 : AOI22_X1 port map( A1 => n6991, A2 => n6730, B1 => n6529, B2 => 
                           intadd_0xBx0x, ZN => n6883);
   U7484 : OAI22_X1 port map( A1 => n6530, A2 => n6581, B1 => n6883, B2 => 
                           ashr_25xSHx3x, ZN => n7134);
   U7485 : AOI22_X1 port map( A1 => n7067, A2 => n6531, B1 => n7416, B2 => 
                           n7134, ZN => n6567);
   U7486 : AOI22_X1 port map( A1 => add_x_26xBx10x, A2 => n7246, B1 => n6532, 
                           B2 => n7443, ZN => n6536);
   U7487 : OAI221_X1 port map( B1 => n7231, B2 => n6534, C1 => ashr_25xSHx3x, 
                           C2 => n6533, A => n6741, ZN => n6535);
   U7488 : OAI211_X1 port map( C1 => n7310, C2 => n6537, A => n6536, B => n6535
                           , ZN => n6564);
   U7489 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn79, A2 => n7172, ZN 
                           => n6562);
   U7490 : INV_X1 port map( A => n6538, ZN => n6542);
   U7491 : AOI22_X1 port map( A1 => n6586, A2 => n6540, B1 => n6539, B2 => 
                           n7263, ZN => n6735);
   U7492 : AOI22_X1 port map( A1 => n7038, A2 => n6735, B1 => n6541, B2 => 
                           n7303, ZN => n6878);
   U7493 : OAI22_X1 port map( A1 => n6542, A2 => n6588, B1 => n6878, B2 => 
                           n7203, ZN => n7133);
   U7494 : NAND2_X1 port map( A1 => n7231, A2 => n6543, ZN => n7138);
   U7495 : INV_X1 port map( A => n7138, ZN => n6544);
   U7496 : AOI22_X1 port map( A1 => n7405, A2 => n7133, B1 => n6630, B2 => 
                           n6544, ZN => n6561);
   U7497 : INV_X1 port map( A => n6545, ZN => n6547);
   U7498 : OAI21_X1 port map( B1 => n6547, B2 => n7203, A => n6546, ZN => n7115
                           );
   U7499 : AND2_X1 port map( A1 => n6548, A2 => n7372, ZN => n6549);
   U7500 : AOI21_X1 port map( B1 => n6550, B2 => n7203, A => n6549, ZN => n6552
                           );
   U7501 : INV_X1 port map( A => n6552, ZN => n6558);
   U7502 : NAND3_X1 port map( A1 => n6708, A2 => n6551, A3 => n7138, ZN => 
                           n7129);
   U7503 : AOI22_X1 port map( A1 => n6687, A2 => n6552, B1 => n6769, B2 => 
                           n7129, ZN => n6557);
   U7504 : OAI21_X1 port map( B1 => n6553, B2 => n7385, A => n7394, ZN => n6554
                           );
   U7505 : NAND2_X1 port map( A1 => n6555, A2 => n6554, ZN => n6556);
   U7506 : OAI211_X1 port map( C1 => n7423, C2 => n6558, A => n6557, B => n6556
                           , ZN => n6559);
   U7507 : AOI21_X1 port map( B1 => n6711, B2 => n7115, A => n6559, ZN => n6560
                           );
   U7508 : NAND3_X1 port map( A1 => n6562, A2 => n6561, A3 => n6560, ZN => 
                           n6563);
   U7509 : AOI211_X1 port map( C1 => n6565, C2 => n7315, A => n6564, B => n6563
                           , ZN => n6566);
   U7510 : OAI211_X1 port map( C1 => n6568, C2 => n7380, A => n6567, B => n6566
                           , ZN => n6569);
   U7511 : AOI22_X1 port map( A1 => n6629, A2 => fromMemoryPortxLOADEDDATAx(10)
                           , B1 => n7023, B2 => n6569, ZN => n6571);
   U7512 : NAND2_X1 port map( A1 => n6572, A2 => ashr_25xAx10x, ZN => n6570);
   U7513 : OAI211_X1 port map( C1 => n6623, C2 => n7118, A => n6571, B => n6570
                           , ZN => IF_ISAxN10947);
   U7514 : AOI22_X1 port map( A1 => n7038, A2 => n6593, B1 => n6757, B2 => 
                           n7303, ZN => n7189);
   U7515 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(11), A2 => n6629
                           , B1 => n6572, B2 => ashr_25xAx11x, ZN => n6622);
   U7516 : INV_X1 port map( A => n6573, ZN => n6574);
   U7517 : AOI21_X1 port map( B1 => intadd_4xBx2x, B2 => n6574, A => n6665, ZN 
                           => n7158);
   U7518 : NOR2_X1 port map( A1 => intadd_2xAx0x, A2 => add_x_26xBx11x, ZN => 
                           n6575);
   U7519 : AOI22_X1 port map( A1 => intadd_0xSUMx9x, A2 => n7270, B1 => n6575, 
                           B2 => n7406, ZN => n6618);
   U7520 : OAI21_X1 port map( B1 => intadd_2xAx0x, B2 => n7385, A => n7394, ZN 
                           => n6615);
   U7521 : OAI221_X1 port map( B1 => n7246, B2 => n7315, C1 => n7246, C2 => 
                           ashr_25xAx11x, A => add_x_26xBx11x, ZN => n6591);
   U7522 : AOI22_X1 port map( A1 => n7414, A2 => n6577, B1 => n6576, B2 => 
                           n7254, ZN => n6760);
   U7523 : AND2_X1 port map( A1 => n6760, A2 => intadd_4xBx1x, ZN => n6578);
   U7524 : AOI21_X1 port map( B1 => n6579, B2 => intadd_0xBx0x, A => n6578, ZN 
                           => n6937);
   U7525 : INV_X1 port map( A => n6937, ZN => n6580);
   U7526 : OAI22_X1 port map( A1 => n6582, A2 => n6581, B1 => n6580, B2 => 
                           ashr_25xSHx3x, ZN => n7166);
   U7527 : INV_X1 port map( A => n6583, ZN => n6589);
   U7528 : AOI22_X1 port map( A1 => n6586, A2 => n6585, B1 => n6584, B2 => 
                           n7263, ZN => n6766);
   U7529 : AOI22_X1 port map( A1 => n7038, A2 => n6766, B1 => n6587, B2 => 
                           n7303, ZN => n6932);
   U7530 : OAI22_X1 port map( A1 => n6589, A2 => n6588, B1 => n6932, B2 => 
                           n7203, ZN => n7185);
   U7531 : AOI22_X1 port map( A1 => n7416, A2 => n7166, B1 => n7405, B2 => 
                           n7185, ZN => n6590);
   U7532 : OAI211_X1 port map( C1 => n7112, C2 => n6592, A => n6591, B => n6590
                           , ZN => n6614);
   U7533 : INV_X1 port map( A => n6593, ZN => n6594);
   U7534 : NAND2_X1 port map( A1 => n7409, A2 => n7262, ZN => n6710);
   U7535 : OAI21_X1 port map( B1 => n7262, B2 => n6594, A => n6710, ZN => n7186
                           );
   U7536 : NOR2_X1 port map( A1 => n6595, A2 => ashr_25xSHx3x, ZN => n7160);
   U7537 : AOI22_X1 port map( A1 => n6711, A2 => n7186, B1 => n6630, B2 => 
                           n7160, ZN => n6610);
   U7538 : NOR2_X1 port map( A1 => intadd_2xBx0x, A2 => ashr_25xAx11x, ZN => 
                           n6597);
   U7539 : AOI221_X1 port map( B1 => intadd_2xAx0x, B2 => n7463, C1 => 
                           ashr_25xAx11x, C2 => n6616, A => n7393, ZN => n6596)
                           ;
   U7540 : AOI21_X1 port map( B1 => n7406, B2 => n6597, A => n6596, ZN => n6609
                           );
   U7541 : AOI22_X1 port map( A1 => n6600, A2 => n6599, B1 => n6598, B2 => 
                           n7303, ZN => n6601);
   U7542 : AND2_X1 port map( A1 => n6601, A2 => n7203, ZN => n6602);
   U7543 : AOI21_X1 port map( B1 => n7372, B2 => n6603, A => n6602, ZN => n6619
                           );
   U7544 : NAND2_X1 port map( A1 => n6687, A2 => n6619, ZN => n6608);
   U7545 : OR2_X1 port map( A1 => n6604, A2 => ashr_25xSHx3x, ZN => n6605);
   U7546 : OAI211_X1 port map( C1 => intadd_4xBx2x, C2 => n6606, A => n6605, B 
                           => n6741, ZN => n6607);
   U7547 : NAND4_X1 port map( A1 => n6610, A2 => n6609, A3 => n6608, A4 => 
                           n6607, ZN => n6611);
   U7548 : AOI21_X1 port map( B1 => DP_OP_719J1_125_1055xn80, B2 => n7364, A =>
                           n6611, ZN => n6612);
   U7549 : INV_X1 port map( A => n6612, ZN => n6613);
   U7550 : AOI211_X1 port map( C1 => n6616, C2 => n6615, A => n6614, B => n6613
                           , ZN => n6617);
   U7551 : OAI211_X1 port map( C1 => n7158, C2 => n6967, A => n6618, B => n6617
                           , ZN => n6620);
   U7552 : AOI22_X1 port map( A1 => n7023, A2 => n6620, B1 => n6628, B2 => 
                           n6619, ZN => n6621);
   U7553 : OAI211_X1 port map( C1 => n7189, C2 => n6623, A => n6622, B => n6621
                           , ZN => IF_ISAxN10948);
   U7554 : NAND2_X1 port map( A1 => n7397, A2 => n6624, ZN => n7234);
   U7555 : INV_X1 port map( A => n6625, ZN => n6626);
   U7556 : AOI22_X1 port map( A1 => n7372, A2 => n6627, B1 => n6626, B2 => 
                           n7203, ZN => n6635);
   U7557 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(12), A2 => n6629
                           , B1 => n6628, B2 => n6635, ZN => n6663);
   U7558 : NAND2_X1 port map( A1 => n7337, A2 => n6630, ZN => n6776);
   U7559 : AOI22_X1 port map( A1 => n7305, A2 => n6632, B1 => n6631, B2 => 
                           n7303, ZN => n6960);
   U7560 : NOR2_X1 port map( A1 => n6633, A2 => n7372, ZN => n6634);
   U7561 : AOI21_X1 port map( B1 => n7372, B2 => n6960, A => n6634, ZN => n7212
                           );
   U7562 : AOI22_X1 port map( A1 => n7212, A2 => n7405, B1 => n6635, B2 => 
                           n6687, ZN => n6636);
   U7563 : INV_X1 port map( A => n6636, ZN => n6653);
   U7564 : MUX2_X1 port map( A => n6638, B => n6637, S => intadd_4xBx1x, Z => 
                           n6970);
   U7565 : INV_X1 port map( A => n6639, ZN => n6959);
   U7566 : NOR2_X1 port map( A1 => n6959, A2 => intadd_4xBx2x, ZN => n6640);
   U7567 : AOI21_X1 port map( B1 => intadd_4xBx2x, B2 => n6970, A => n6640, ZN 
                           => n7210);
   U7568 : AOI21_X1 port map( B1 => n7231, B2 => n6641, A => n6665, ZN => n7217
                           );
   U7569 : OAI22_X1 port map( A1 => n7210, A2 => n7339, B1 => n7217, B2 => 
                           n6967, ZN => n6652);
   U7570 : OAI22_X1 port map( A1 => n6643, A2 => n7380, B1 => n6642, B2 => 
                           n7310, ZN => n6651);
   U7571 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn81, A2 => n7364, ZN 
                           => n6649);
   U7572 : NAND2_X1 port map( A1 => n6710, A2 => n7234, ZN => n7224);
   U7573 : AOI22_X1 port map( A1 => n6711, A2 => n7224, B1 => n6644, B2 => 
                           n7443, ZN => n6648);
   U7574 : OAI22_X1 port map( A1 => intadd_2xBx1x, A2 => n7223, B1 => n6645, B2
                           => n7393, ZN => n6646);
   U7575 : AOI21_X1 port map( B1 => n7318, B2 => n6658, A => n6646, ZN => n6647
                           );
   U7576 : NAND3_X1 port map( A1 => n6649, A2 => n6648, A3 => n6647, ZN => 
                           n6650);
   U7577 : NOR4_X1 port map( A1 => n6653, A2 => n6652, A3 => n6651, A4 => n6650
                           , ZN => n6657);
   U7578 : OAI221_X1 port map( B1 => intadd_4xBx2x, B2 => n6655, C1 => 
                           ashr_25xSHx3x, C2 => n6654, A => n6741, ZN => n6656)
                           ;
   U7579 : OAI211_X1 port map( C1 => n7240, C2 => n6776, A => n6657, B => n6656
                           , ZN => n6661);
   U7580 : AOI221_X1 port map( B1 => n7323, B2 => n7464, C1 => n7248, C2 => 
                           n6658, A => n7246, ZN => n6659);
   U7581 : OAI221_X1 port map( B1 => intadd_2xBx1x, B2 => n7382, C1 => 
                           add_x_26xBx12x, C2 => n7250, A => n6659, ZN => n6660
                           );
   U7582 : OAI221_X1 port map( B1 => n6661, B2 => ashr_25xAx12x, C1 => n6661, 
                           C2 => n6660, A => n7023, ZN => n6662);
   U7583 : OAI211_X1 port map( C1 => n6664, C2 => n7234, A => n6663, B => n6662
                           , ZN => IF_ISAxN10949);
   U7584 : AOI21_X1 port map( B1 => intadd_4xBx2x, B2 => n6666, A => n6665, ZN 
                           => n7281);
   U7585 : INV_X1 port map( A => n7223, ZN => n7376);
   U7586 : AOI22_X1 port map( A1 => n6667, A2 => n7443, B1 => add_x_26xBx13x, 
                           B2 => n7376, ZN => n6671);
   U7587 : OAI221_X1 port map( B1 => intadd_4xBx2x, B2 => n6669, C1 => 
                           ashr_25xSHx3x, C2 => n6668, A => n6741, ZN => n6670)
                           ;
   U7588 : OAI211_X1 port map( C1 => n7281, C2 => n6967, A => n6671, B => n6670
                           , ZN => n6701);
   U7589 : NAND2_X1 port map( A1 => n6672, A2 => n7203, ZN => n6675);
   U7590 : NAND2_X1 port map( A1 => n6673, A2 => n7372, ZN => n6674);
   U7591 : NAND2_X1 port map( A1 => n6675, A2 => n6674, ZN => n6699);
   U7592 : AOI22_X1 port map( A1 => n7372, A2 => n6677, B1 => n6676, B2 => 
                           n7203, ZN => n7276);
   U7593 : NAND2_X1 port map( A1 => n7397, A2 => n6678, ZN => n7278);
   U7594 : AOI22_X1 port map( A1 => n7231, A2 => n6680, B1 => n6679, B2 => 
                           ashr_25xSHx3x, ZN => n7277);
   U7595 : OAI22_X1 port map( A1 => n6763, A2 => n7278, B1 => n7339, B2 => 
                           n7277, ZN => n6681);
   U7596 : AOI21_X1 port map( B1 => n7405, B2 => n7276, A => n6681, ZN => n6698
                           );
   U7597 : INV_X1 port map( A => intadd_0xSUMx11x, ZN => n6683);
   U7598 : OAI22_X1 port map( A1 => n6683, A2 => n7380, B1 => n6682, B2 => 
                           n7310, ZN => n6696);
   U7599 : INV_X1 port map( A => n6684, ZN => n6685);
   U7600 : OAI21_X1 port map( B1 => n6685, B2 => n7262, A => n6710, ZN => n7271
                           );
   U7601 : INV_X1 port map( A => n6699, ZN => n6686);
   U7602 : AOI222_X1 port map( A1 => DP_OP_719J1_125_1055xn82, A2 => n7364, B1 
                           => n6711, B2 => n7271, C1 => n6687, C2 => n6686, ZN 
                           => n6688);
   U7603 : INV_X1 port map( A => n6688, ZN => n6695);
   U7604 : AOI21_X1 port map( B1 => n6690, B2 => n6689, A => n7393, ZN => n6694
                           );
   U7605 : OAI221_X1 port map( B1 => intadd_2xBx2x, B2 => n7382, C1 => 
                           add_x_26xBx13x, C2 => n7250, A => n7383, ZN => n6691
                           );
   U7606 : AOI21_X1 port map( B1 => n7248, B2 => n6702, A => n6691, ZN => n6692
                           );
   U7607 : OAI22_X1 port map( A1 => n7280, A2 => n6776, B1 => intadd_2xAx2x, B2
                           => n6692, ZN => n6693);
   U7608 : NOR4_X1 port map( A1 => n6696, A2 => n6695, A3 => n6694, A4 => n6693
                           , ZN => n6697);
   U7609 : OAI211_X1 port map( C1 => n7423, C2 => n6699, A => n6698, B => n6697
                           , ZN => n6700);
   U7610 : AOI211_X1 port map( C1 => n7318, C2 => n6702, A => n6701, B => n6700
                           , ZN => n6704);
   U7611 : OAI22_X1 port map( A1 => n6704, A2 => n6829, B1 => n6703, B2 => 
                           n7435, ZN => IF_ISAxN10950);
   U7612 : NAND2_X1 port map( A1 => n7397, A2 => n6705, ZN => n7338);
   U7613 : INV_X1 port map( A => n7338, ZN => n6749);
   U7614 : OR2_X1 port map( A1 => n6706, A2 => ashr_25xSHx3x, ZN => n6707);
   U7615 : AND2_X1 port map( A1 => n6708, A2 => n6707, ZN => n7326);
   U7616 : INV_X1 port map( A => n7326, ZN => n6712);
   U7617 : NAND3_X1 port map( A1 => n7338, A2 => n6710, A3 => n6709, ZN => 
                           n7346);
   U7618 : AOI222_X1 port map( A1 => n6712, A2 => n6769, B1 => n7346, B2 => 
                           n6711, C1 => n7364, C2 => DP_OP_719J1_125_1055xn83, 
                           ZN => n6713);
   U7619 : INV_X1 port map( A => n6713, ZN => n6748);
   U7620 : AOI22_X1 port map( A1 => n7038, A2 => n6715, B1 => n6714, B2 => 
                           n7303, ZN => n6718);
   U7621 : INV_X1 port map( A => n6716, ZN => n6717);
   U7622 : AOI221_X1 port map( B1 => n6719, B2 => n7372, C1 => n6718, C2 => 
                           n7203, A => n6717, ZN => n6740);
   U7623 : OAI22_X1 port map( A1 => intadd_2xBx3x, A2 => n7223, B1 => n7112, B2
                           => n6720, ZN => n6725);
   U7624 : OAI221_X1 port map( B1 => n7466, B2 => n7385, C1 => n6726, C2 => 
                           n7313, A => n7383, ZN => n6721);
   U7625 : AOI221_X1 port map( B1 => n7406, B2 => intadd_2xBx3x, C1 => n7315, 
                           C2 => add_x_26xBx14x, A => n6721, ZN => n6723);
   U7626 : OAI22_X1 port map( A1 => intadd_2xAx3x, A2 => n6723, B1 => n7310, B2
                           => n6722, ZN => n6724);
   U7627 : AOI211_X1 port map( C1 => n7318, C2 => n6726, A => n6725, B => n6724
                           , ZN => n6738);
   U7628 : NOR2_X1 port map( A1 => n7466, A2 => ashr_25xAx14x, ZN => n6727);
   U7629 : AOI22_X1 port map( A1 => n6727, A2 => n7067, B1 => intadd_0xSUMx12x,
                           B2 => n7270, ZN => n6737);
   U7630 : AOI22_X1 port map( A1 => n7414, A2 => n6729, B1 => n6728, B2 => 
                           n7125, ZN => n6876);
   U7631 : AOI22_X1 port map( A1 => n6991, A2 => n6876, B1 => n6730, B2 => 
                           n7046, ZN => n6996);
   U7632 : AND2_X1 port map( A1 => n6731, A2 => ashr_25xSHx3x, ZN => n6732);
   U7633 : AOI21_X1 port map( B1 => intadd_4xBx2x, B2 => n6996, A => n6732, ZN 
                           => n7347);
   U7634 : AOI22_X1 port map( A1 => n7164, A2 => n6734, B1 => n6733, B2 => 
                           n7399, ZN => n6882);
   U7635 : AOI22_X1 port map( A1 => n7038, A2 => n6882, B1 => n6735, B2 => 
                           n7303, ZN => n7007);
   U7636 : AOI22_X1 port map( A1 => n7372, A2 => n7007, B1 => n7008, B2 => 
                           n7203, ZN => n7343);
   U7637 : AOI22_X1 port map( A1 => n7416, A2 => n7347, B1 => n7405, B2 => 
                           n7343, ZN => n6736);
   U7638 : NAND3_X1 port map( A1 => n6738, A2 => n6737, A3 => n6736, ZN => 
                           n6739);
   U7639 : NOR2_X1 port map( A1 => n6740, A2 => n6739, ZN => n6745);
   U7640 : OAI221_X1 port map( B1 => intadd_4xBx2x, B2 => n6743, C1 => 
                           ashr_25xSHx3x, C2 => n6742, A => n6741, ZN => n6744)
                           ;
   U7641 : OAI211_X1 port map( C1 => n6776, C2 => n6746, A => n6745, B => n6744
                           , ZN => n6747);
   U7642 : AOI211_X1 port map( C1 => n6750, C2 => n6749, A => n6748, B => n6747
                           , ZN => n6752);
   U7643 : OAI22_X1 port map( A1 => n6752, A2 => n6829, B1 => n6751, B2 => 
                           n7435, ZN => IF_ISAxN10951);
   U7644 : INV_X1 port map( A => n6753, ZN => n6755);
   U7645 : AOI221_X1 port map( B1 => n6756, B2 => ashr_25xSHx3x, C1 => n6755, 
                           C2 => intadd_4xBx2x, A => n6754, ZN => n6793);
   U7646 : NAND2_X1 port map( A1 => n7397, A2 => n6757, ZN => n7422);
   U7647 : AOI22_X1 port map( A1 => n7414, A2 => n6759, B1 => n6758, B2 => 
                           n7412, ZN => n6926);
   U7648 : AOI22_X1 port map( A1 => n6991, A2 => n6926, B1 => n6760, B2 => 
                           intadd_0xBx0x, ZN => n7054);
   U7649 : INV_X1 port map( A => n7040, ZN => n6761);
   U7650 : NOR2_X1 port map( A1 => n6761, A2 => intadd_4xBx2x, ZN => n6762);
   U7651 : AOI21_X1 port map( B1 => intadd_4xBx2x, B2 => n7054, A => n6762, ZN 
                           => n7367);
   U7652 : OAI22_X1 port map( A1 => n6763, A2 => n7422, B1 => n7339, B2 => 
                           n7367, ZN => n6792);
   U7653 : AOI22_X1 port map( A1 => n7164, A2 => n6765, B1 => n6764, B2 => 
                           n7082, ZN => n6930);
   U7654 : AOI22_X1 port map( A1 => n7305, A2 => n6930, B1 => n6766, B2 => 
                           n7036, ZN => n7371);
   U7655 : NOR2_X1 port map( A1 => n7467, A2 => ashr_25xAx15x, ZN => n6767);
   U7656 : AOI22_X1 port map( A1 => n6767, A2 => n7067, B1 => intadd_0xSUMx13x,
                           B2 => n7270, ZN => n6771);
   U7657 : NOR3_X1 port map( A1 => n7202, A2 => n7044, A3 => n7372, ZN => n6768
                           );
   U7658 : AOI21_X1 port map( B1 => n6769, B2 => n7409, A => n6768, ZN => n6770
                           );
   U7659 : OAI211_X1 port map( C1 => n7371, C2 => n6997, A => n6771, B => n6770
                           , ZN => n6772);
   U7660 : AOI21_X1 port map( B1 => DP_OP_719J1_125_1055xn84, B2 => n7172, A =>
                           n6772, ZN => n6773);
   U7661 : INV_X1 port map( A => n6773, ZN => n6791);
   U7662 : OAI221_X1 port map( B1 => n7467, B2 => n7385, C1 => n6774, C2 => 
                           n7313, A => n7383, ZN => n6775);
   U7663 : AOI21_X1 port map( B1 => n7315, B2 => add_x_26xBx15x, A => n6775, ZN
                           => n6788);
   U7664 : INV_X1 port map( A => n6776, ZN => n6782);
   U7665 : OAI22_X1 port map( A1 => n6778, A2 => n7223, B1 => n7112, B2 => 
                           n6777, ZN => n6781);
   U7666 : OAI22_X1 port map( A1 => n6779, A2 => n7310, B1 => n7467, B2 => 
                           n7394, ZN => n6780);
   U7667 : AOI211_X1 port map( C1 => n7392, C2 => n6782, A => n6781, B => n6780
                           , ZN => n6787);
   U7668 : OAI221_X1 port map( B1 => n7372, B2 => n6784, C1 => n7203, C2 => 
                           n6783, A => n7081, ZN => n6785);
   U7669 : OAI21_X1 port map( B1 => n7013, B2 => n7349, A => n6785, ZN => n6786
                           );
   U7670 : OAI211_X1 port map( C1 => n6789, C2 => n6788, A => n6787, B => n6786
                           , ZN => n6790);
   U7671 : NOR4_X1 port map( A1 => n6793, A2 => n6792, A3 => n6791, A4 => n6790
                           , ZN => n6795);
   U7672 : OAI22_X1 port map( A1 => n6795, A2 => n6829, B1 => n6794, B2 => 
                           n7435, ZN => IF_ISAxN10952);
   U7673 : INV_X1 port map( A => n7427, ZN => n6995);
   U7674 : OAI22_X1 port map( A1 => n6797, A2 => n6997, B1 => n6796, B2 => 
                           n6995, ZN => n6827);
   U7675 : INV_X1 port map( A => n7049, ZN => n6879);
   U7676 : OAI22_X1 port map( A1 => n6799, A2 => n6879, B1 => n6798, B2 => 
                           n7308, ZN => n6826);
   U7677 : AOI22_X1 port map( A1 => n7315, A2 => add_x_26xBx16x, B1 => n7248, 
                           B2 => n6805, ZN => n6801);
   U7678 : OAI21_X1 port map( B1 => n6814, B2 => n7345, A => n7349, ZN => n6800
                           );
   U7679 : OAI221_X1 port map( B1 => n6802, B2 => n6801, C1 => n6802, C2 => 
                           n7383, A => n6800, ZN => n6825);
   U7680 : AOI22_X1 port map( A1 => n7270, A2 => intadd_0xSUMx14x, B1 => n7406,
                           B2 => n6803, ZN => n6821);
   U7681 : AOI21_X1 port map( B1 => n7327, B2 => n6817, A => n7325, ZN => n6813
                           );
   U7682 : AOI22_X1 port map( A1 => n7318, A2 => n6805, B1 => n6804, B2 => 
                           n7443, ZN => n6810);
   U7683 : INV_X1 port map( A => n6806, ZN => n6808);
   U7684 : OAI21_X1 port map( B1 => n6808, B2 => n6807, A => n7323, ZN => n6809
                           );
   U7685 : OAI211_X1 port map( C1 => n6811, C2 => n7223, A => n6810, B => n6809
                           , ZN => n6812);
   U7686 : AOI211_X1 port map( C1 => n7013, C2 => n6814, A => n6813, B => n6812
                           , ZN => n6820);
   U7687 : AOI22_X1 port map( A1 => n6816, A2 => n7348, B1 => n6815, B2 => 
                           n7344, ZN => n6819);
   U7688 : OR2_X1 port map( A1 => n6817, A2 => n7216, ZN => n6818);
   U7689 : NAND4_X1 port map( A1 => n6821, A2 => n6820, A3 => n6819, A4 => 
                           n6818, ZN => n6822);
   U7690 : AOI21_X1 port map( B1 => n7364, B2 => DP_OP_719J1_125_1055xn85, A =>
                           n6822, ZN => n6823);
   U7691 : INV_X1 port map( A => n6823, ZN => n6824);
   U7692 : NOR4_X1 port map( A1 => n6827, A2 => n6826, A3 => n6825, A4 => n6824
                           , ZN => n6830);
   U7693 : OAI22_X1 port map( A1 => n6830, A2 => n6829, B1 => n6828, B2 => 
                           n7435, ZN => IF_ISAxN10953);
   U7694 : AOI22_X1 port map( A1 => n6831, A2 => n7067, B1 => intadd_0xSUMx15x,
                           B2 => n7270, ZN => n6833);
   U7695 : AOI22_X1 port map( A1 => n7318, A2 => n6835, B1 => add_x_26xBx17x, 
                           B2 => n7376, ZN => n6832);
   U7696 : OAI211_X1 port map( C1 => n7112, C2 => n6834, A => n6833, B => n6832
                           , ZN => n6866);
   U7697 : OAI221_X1 port map( B1 => n7469, B2 => n7385, C1 => n6835, C2 => 
                           n7313, A => n7383, ZN => n6836);
   U7698 : AOI221_X1 port map( B1 => n7406, B2 => intadd_1xBx0x, C1 => n7315, 
                           C2 => add_x_26xBx17x, A => n6836, ZN => n6839);
   U7699 : INV_X1 port map( A => n6837, ZN => n6838);
   U7700 : OAI22_X1 port map( A1 => intadd_1xAx0x, A2 => n6839, B1 => n7310, B2
                           => n6838, ZN => n6865);
   U7701 : AOI22_X1 port map( A1 => n6991, A2 => n6841, B1 => n6840, B2 => 
                           intadd_0xBx0x, ZN => n7107);
   U7702 : AOI22_X1 port map( A1 => n7427, A2 => n6842, B1 => n7049, B2 => 
                           n7107, ZN => n6845);
   U7703 : OAI21_X1 port map( B1 => n6843, B2 => n7345, A => n7349, ZN => n6844
                           );
   U7704 : OAI211_X1 port map( C1 => n7308, C2 => n6846, A => n6845, B => n6844
                           , ZN => n6864);
   U7705 : AND2_X1 port map( A1 => DP_OP_719J1_125_1055xn86, A2 => n7364, ZN =>
                           n6862);
   U7706 : INV_X1 port map( A => n7344, ZN => n7369);
   U7707 : OAI22_X1 port map( A1 => n7369, A2 => n6848, B1 => n7216, B2 => 
                           n6847, ZN => n6861);
   U7708 : OR2_X1 port map( A1 => n6849, A2 => n7036, ZN => n6852);
   U7709 : NAND2_X1 port map( A1 => n6850, A2 => n7036, ZN => n6851);
   U7710 : AND2_X1 port map( A1 => n6852, A2 => n6851, ZN => n7075);
   U7711 : INV_X1 port map( A => n7075, ZN => n6853);
   U7712 : NAND2_X1 port map( A1 => n7301, A2 => n6853, ZN => n6854);
   U7713 : NOR2_X1 port map( A1 => n7325, A2 => n7327, ZN => n7283);
   U7714 : INV_X1 port map( A => n7283, ZN => n7157);
   U7715 : OAI211_X1 port map( C1 => n7325, C2 => n6855, A => n6854, B => n7157
                           , ZN => n6860);
   U7716 : AOI22_X1 port map( A1 => n7013, A2 => n6857, B1 => n7348, B2 => 
                           n6856, ZN => n6858);
   U7717 : INV_X1 port map( A => n6858, ZN => n6859);
   U7718 : OR4_X1 port map( A1 => n6862, A2 => n6861, A3 => n6860, A4 => n6859,
                           ZN => n6863);
   U7719 : NOR4_X1 port map( A1 => n6866, A2 => n6865, A3 => n6864, A4 => n6863
                           , ZN => n6868);
   U7720 : OAI22_X1 port map( A1 => n6868, A2 => n7529, B1 => n6867, B2 => 
                           n7435, ZN => IF_ISAxN10954);
   U7721 : NAND2_X1 port map( A1 => n7081, A2 => n6869, ZN => n6870);
   U7722 : AOI22_X1 port map( A1 => n7159, A2 => n6871, B1 => n7349, B2 => 
                           n6870, ZN => n6872);
   U7723 : OAI21_X1 port map( B1 => n7369, B2 => n6873, A => n6872, ZN => n6906
                           );
   U7724 : AOI22_X1 port map( A1 => n7414, A2 => n6875, B1 => n6874, B2 => 
                           n7254, ZN => n6990);
   U7725 : INV_X1 port map( A => n6990, ZN => n6877);
   U7726 : AOI22_X1 port map( A1 => n6991, A2 => n6877, B1 => n6876, B2 => 
                           intadd_0xBx0x, ZN => n7131);
   U7727 : OAI22_X1 port map( A1 => n7131, A2 => n6879, B1 => n6878, B2 => 
                           n7308, ZN => n6905);
   U7728 : AOI22_X1 port map( A1 => n7164, A2 => n6881, B1 => n6880, B2 => 
                           n7082, ZN => n6994);
   U7729 : AOI22_X1 port map( A1 => n7038, A2 => n6994, B1 => n6882, B2 => 
                           n7036, ZN => n7119);
   U7730 : OAI22_X1 port map( A1 => n7119, A2 => n6997, B1 => n6883, B2 => 
                           n6995, ZN => n6904);
   U7731 : INV_X1 port map( A => intadd_0xSUMx16x, ZN => n6884);
   U7732 : OAI22_X1 port map( A1 => n6885, A2 => n7313, B1 => n6884, B2 => 
                           n7380, ZN => n6901);
   U7733 : AOI221_X1 port map( B1 => n7323, B2 => n7470, C1 => n7248, C2 => 
                           n6891, A => n7246, ZN => n6886);
   U7734 : OAI221_X1 port map( B1 => intadd_1xBx1x, B2 => n7382, C1 => 
                           add_x_26xBx18x, C2 => n7250, A => n6886, ZN => n6898
                           );
   U7735 : INV_X1 port map( A => n7348, ZN => n7366);
   U7736 : OAI22_X1 port map( A1 => n6888, A2 => n7423, B1 => n7366, B2 => 
                           n6887, ZN => n6897);
   U7737 : OAI22_X1 port map( A1 => intadd_1xBx1x, A2 => n7223, B1 => n7112, B2
                           => n6889, ZN => n6890);
   U7738 : AOI211_X1 port map( C1 => n7318, C2 => n6891, A => n6890, B => n7283
                           , ZN => n6895);
   U7739 : NOR2_X1 port map( A1 => intadd_1xBx1x, A2 => ashr_25xAx18x, ZN => 
                           n6892);
   U7740 : AOI22_X1 port map( A1 => n7130, A2 => n6893, B1 => n6892, B2 => 
                           n7406, ZN => n6894);
   U7741 : NAND2_X1 port map( A1 => n6895, A2 => n6894, ZN => n6896);
   U7742 : AOI211_X1 port map( C1 => n6898, C2 => ashr_25xAx18x, A => n6897, B 
                           => n6896, ZN => n6899);
   U7743 : INV_X1 port map( A => n6899, ZN => n6900);
   U7744 : AOI211_X1 port map( C1 => DP_OP_719J1_125_1055xn87, C2 => n7172, A 
                           => n6901, B => n6900, ZN => n6902);
   U7745 : INV_X1 port map( A => n6902, ZN => n6903);
   U7746 : NOR4_X1 port map( A1 => n6906, A2 => n6905, A3 => n6904, A4 => n6903
                           , ZN => n6908);
   U7747 : OAI22_X1 port map( A1 => n6908, A2 => n7529, B1 => n6907, B2 => 
                           n7435, ZN => IF_ISAxN10955);
   U7748 : AOI22_X1 port map( A1 => n7013, A2 => n6910, B1 => n7159, B2 => 
                           n6909, ZN => n6913);
   U7749 : OAI21_X1 port map( B1 => n6911, B2 => ashr_25xSHx4x, A => n7130, ZN 
                           => n6912);
   U7750 : OAI211_X1 port map( C1 => n6914, C2 => n7369, A => n6913, B => n6912
                           , ZN => n6944);
   U7751 : INV_X1 port map( A => n6915, ZN => n6916);
   U7752 : OAI22_X1 port map( A1 => n6917, A2 => n7313, B1 => n6916, B2 => 
                           n7310, ZN => n6943);
   U7753 : AOI22_X1 port map( A1 => n7318, A2 => n6918, B1 => add_x_26xBx19x, 
                           B2 => n7376, ZN => n6922);
   U7754 : AOI221_X1 port map( B1 => n7323, B2 => n7471, C1 => n7248, C2 => 
                           n6918, A => n7246, ZN => n6919);
   U7755 : OAI221_X1 port map( B1 => intadd_1xBx2x, B2 => n7382, C1 => 
                           add_x_26xBx19x, C2 => n7310, A => n6919, ZN => n6920
                           );
   U7756 : AOI22_X1 port map( A1 => n7270, A2 => intadd_0xSUMx17x, B1 => 
                           ashr_25xAx19x, B2 => n6920, ZN => n6921);
   U7757 : OAI211_X1 port map( C1 => n7112, C2 => n6923, A => n6922, B => n6921
                           , ZN => n6942);
   U7758 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn88, A2 => n7364, ZN 
                           => n6940);
   U7759 : AOI22_X1 port map( A1 => n7414, A2 => n6925, B1 => n6924, B2 => 
                           n7412, ZN => n7047);
   U7760 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n7047, B1 => n6926, B2
                           => intadd_0xBx0x, ZN => n7193);
   U7761 : AOI21_X1 port map( B1 => n7081, B2 => n6927, A => n7079, ZN => n6934
                           );
   U7762 : AOI22_X1 port map( A1 => n7164, A2 => n6929, B1 => n6928, B2 => 
                           n7263, ZN => n7037);
   U7763 : INV_X1 port map( A => n7037, ZN => n6931);
   U7764 : AOI22_X1 port map( A1 => n7305, A2 => n6931, B1 => n6930, B2 => 
                           n7036, ZN => n7190);
   U7765 : OAI22_X1 port map( A1 => n7190, A2 => n6997, B1 => n6932, B2 => 
                           n7308, ZN => n6933);
   U7766 : AOI211_X1 port map( C1 => n7049, C2 => n7193, A => n6934, B => n6933
                           , ZN => n6939);
   U7767 : INV_X1 port map( A => n6935, ZN => n6936);
   U7768 : AOI22_X1 port map( A1 => n7427, A2 => n6937, B1 => n7348, B2 => 
                           n6936, ZN => n6938);
   U7769 : NAND3_X1 port map( A1 => n6940, A2 => n6939, A3 => n6938, ZN => 
                           n6941);
   U7770 : NOR4_X1 port map( A1 => n6944, A2 => n6943, A3 => n6942, A4 => n6941
                           , ZN => n6946);
   U7771 : OAI22_X1 port map( A1 => n6946, A2 => n7529, B1 => n6945, B2 => 
                           n7435, ZN => IF_ISAxN10956);
   U7772 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn89, A2 => n7364, ZN 
                           => n6954);
   U7773 : AOI22_X1 port map( A1 => intadd_0xSUMx18x, A2 => n7270, B1 => n6947,
                           B2 => n7406, ZN => n6953);
   U7774 : INV_X1 port map( A => n6948, ZN => n6951);
   U7775 : INV_X1 port map( A => n6949, ZN => n6950);
   U7776 : AOI22_X1 port map( A1 => n7013, A2 => n6951, B1 => n7159, B2 => 
                           n6950, ZN => n6952);
   U7777 : NAND3_X1 port map( A1 => n6954, A2 => n6953, A3 => n6952, ZN => 
                           n6981);
   U7778 : OAI211_X1 port map( C1 => n7318, C2 => n7323, A => intadd_1xAx3x, B 
                           => n6962, ZN => n6957);
   U7779 : AOI22_X1 port map( A1 => n6955, A2 => n7443, B1 => add_x_26xBx20x, 
                           B2 => n7376, ZN => n6956);
   U7780 : OAI211_X1 port map( C1 => n6959, C2 => n6958, A => n6957, B => n6956
                           , ZN => n6980);
   U7781 : OAI22_X1 port map( A1 => n6961, A2 => n7043, B1 => n6960, B2 => 
                           n7308, ZN => n6979);
   U7782 : OAI221_X1 port map( B1 => n7472, B2 => n7385, C1 => n6962, C2 => 
                           n7313, A => n7383, ZN => n6963);
   U7783 : AOI221_X1 port map( B1 => n7406, B2 => intadd_1xBx3x, C1 => n7315, 
                           C2 => add_x_26xBx20x, A => n6963, ZN => n6977);
   U7784 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n6965, B1 => n6964, B2
                           => intadd_0xBx0x, ZN => n7230);
   U7785 : AOI22_X1 port map( A1 => n7431, A2 => ashr_25xSHx4x, B1 => n6967, B2
                           => n6966, ZN => n6973);
   U7786 : AOI22_X1 port map( A1 => n7305, A2 => n6969, B1 => n6968, B2 => 
                           n7036, ZN => n7204);
   U7787 : INV_X1 port map( A => n6970, ZN => n6971);
   U7788 : OAI22_X1 port map( A1 => n7204, A2 => n6997, B1 => n6971, B2 => 
                           n6995, ZN => n6972);
   U7789 : AOI211_X1 port map( C1 => n7049, C2 => n7230, A => n6973, B => n6972
                           , ZN => n6976);
   U7790 : OAI21_X1 port map( B1 => n7345, B2 => n6974, A => n7349, ZN => n6975
                           );
   U7791 : OAI211_X1 port map( C1 => intadd_1xAx3x, C2 => n6977, A => n6976, B 
                           => n6975, ZN => n6978);
   U7792 : NOR4_X1 port map( A1 => n6981, A2 => n6980, A3 => n6979, A4 => n6978
                           , ZN => n6983);
   U7793 : OAI22_X1 port map( A1 => n6983, A2 => n7529, B1 => n6982, B2 => 
                           n7435, ZN => IF_ISAxN10957);
   U7794 : AOI221_X1 port map( B1 => n7323, B2 => n7474, C1 => n7248, C2 => 
                           n6986, A => n7246, ZN => n6984);
   U7795 : OAI221_X1 port map( B1 => intadd_1xBx5x, B2 => n7382, C1 => 
                           add_x_26xBx22x, C2 => n7250, A => n6984, ZN => n6985
                           );
   U7796 : AOI22_X1 port map( A1 => n7270, A2 => intadd_0xSUMx20x, B1 => 
                           ashr_25xAx22x, B2 => n6985, ZN => n7003);
   U7797 : AOI22_X1 port map( A1 => n7159, A2 => n6987, B1 => n7318, B2 => 
                           n6986, ZN => n7002);
   U7798 : AOI22_X1 port map( A1 => n7414, A2 => n6989, B1 => n6988, B2 => 
                           n7412, ZN => n7127);
   U7799 : AOI22_X1 port map( A1 => n6991, A2 => n7127, B1 => n6990, B2 => 
                           intadd_0xBx0x, ZN => n7293);
   U7800 : AOI22_X1 port map( A1 => n7164, A2 => n6993, B1 => n6992, B2 => 
                           n7399, ZN => n7137);
   U7801 : AOI22_X1 port map( A1 => n7305, A2 => n7137, B1 => n6994, B2 => 
                           n7036, ZN => n7309);
   U7802 : OAI22_X1 port map( A1 => n7309, A2 => n6997, B1 => n6996, B2 => 
                           n6995, ZN => n6998);
   U7803 : AOI21_X1 port map( B1 => n7049, B2 => n7293, A => n6998, ZN => n7001
                           );
   U7804 : OAI21_X1 port map( B1 => n7345, B2 => n6999, A => n7349, ZN => n7000
                           );
   U7805 : NAND4_X1 port map( A1 => n7003, A2 => n7002, A3 => n7001, A4 => 
                           n7000, ZN => n7025);
   U7806 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn91, A2 => n7364, ZN 
                           => n7022);
   U7807 : INV_X1 port map( A => n7004, ZN => n7006);
   U7808 : OAI22_X1 port map( A1 => n7006, A2 => n7393, B1 => n7005, B2 => 
                           n7310, ZN => n7010);
   U7809 : OAI22_X1 port map( A1 => n7008, A2 => n7043, B1 => n7007, B2 => 
                           n7308, ZN => n7009);
   U7810 : AOI211_X1 port map( C1 => n7039, C2 => n7011, A => n7010, B => n7009
                           , ZN => n7021);
   U7811 : NAND2_X1 port map( A1 => n7013, A2 => n7012, ZN => n7017);
   U7812 : NOR2_X1 port map( A1 => n7112, A2 => n7014, ZN => n7015);
   U7813 : AOI21_X1 port map( B1 => add_x_26xBx22x, B2 => n7376, A => n7015, ZN
                           => n7016);
   U7814 : NAND2_X1 port map( A1 => n7017, A2 => n7016, ZN => n7018);
   U7815 : AOI211_X1 port map( C1 => n7019, C2 => n7130, A => n7283, B => n7018
                           , ZN => n7020);
   U7816 : NAND3_X1 port map( A1 => n7022, A2 => n7021, A3 => n7020, ZN => 
                           n7024);
   U7817 : OAI21_X1 port map( B1 => n7025, B2 => n7024, A => n7023, ZN => n7026
                           );
   U7818 : OAI21_X1 port map( B1 => n7435, B2 => n7027, A => n7026, ZN => 
                           IF_ISAxN10959);
   U7819 : AOI221_X1 port map( B1 => n7323, B2 => n7475, C1 => n7248, C2 => 
                           n7028, A => n7246, ZN => n7029);
   U7820 : OAI221_X1 port map( B1 => intadd_1xBx6x, B2 => n7382, C1 => 
                           add_x_26xBx23x, C2 => n7250, A => n7029, ZN => n7064
                           );
   U7821 : AOI22_X1 port map( A1 => intadd_0xSUMx21x, A2 => n7270, B1 => n7030,
                           B2 => n7406, ZN => n7031);
   U7822 : OAI21_X1 port map( B1 => n7032, B2 => n7216, A => n7031, ZN => n7063
                           );
   U7823 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn92, A2 => n7364, ZN 
                           => n7061);
   U7824 : AOI22_X1 port map( A1 => n7067, A2 => n7034, B1 => n7033, B2 => 
                           n7443, ZN => n7042);
   U7825 : AOI22_X1 port map( A1 => n7205, A2 => intadd_1xAx6x, B1 => 
                           intadd_1xAx5x, B2 => n7395, ZN => n7083);
   U7826 : AOI22_X1 port map( A1 => n7164, A2 => n7083, B1 => n7035, B2 => 
                           n7263, ZN => n7165);
   U7827 : AOI22_X1 port map( A1 => n7038, A2 => n7165, B1 => n7037, B2 => 
                           n7036, ZN => n7389);
   U7828 : AOI22_X1 port map( A1 => n7040, A2 => n7039, B1 => n7301, B2 => 
                           n7389, ZN => n7041);
   U7829 : OAI211_X1 port map( C1 => n7044, C2 => n7043, A => n7042, B => n7041
                           , ZN => n7053);
   U7830 : AOI22_X1 port map( A1 => n7329, A2 => intadd_1xAx6x, B1 => 
                           intadd_1xAx5x, B2 => n7408, ZN => n7087);
   U7831 : AOI22_X1 port map( A1 => n7414, A2 => n7087, B1 => n7045, B2 => 
                           n7412, ZN => n7175);
   U7832 : AOI22_X1 port map( A1 => intadd_4xBx1x, A2 => n7175, B1 => n7047, B2
                           => n7046, ZN => n7426);
   U7833 : INV_X1 port map( A => n7371, ZN => n7048);
   U7834 : AOI22_X1 port map( A1 => n7049, A2 => n7426, B1 => n7390, B2 => 
                           n7048, ZN => n7050);
   U7835 : OAI221_X1 port map( B1 => n7079, B2 => n7081, C1 => n7079, C2 => 
                           n7051, A => n7050, ZN => n7052);
   U7836 : AOI211_X1 port map( C1 => n7427, C2 => n7054, A => n7053, B => n7052
                           , ZN => n7060);
   U7837 : OAI22_X1 port map( A1 => n7423, A2 => n7055, B1 => n7223, B2 => 
                           intadd_1xBx6x, ZN => n7058);
   U7838 : OAI22_X1 port map( A1 => n7394, A2 => n7475, B1 => n7325, B2 => 
                           n7056, ZN => n7057);
   U7839 : NOR3_X1 port map( A1 => n7058, A2 => n7057, A3 => n7283, ZN => n7059
                           );
   U7840 : NAND3_X1 port map( A1 => n7061, A2 => n7060, A3 => n7059, ZN => 
                           n7062);
   U7841 : AOI211_X1 port map( C1 => ashr_25xAx23x, C2 => n7064, A => n7063, B 
                           => n7062, ZN => n7066);
   U7842 : OAI22_X1 port map( A1 => n7066, A2 => n7529, B1 => n7065, B2 => 
                           n7435, ZN => IF_ISAxN10960);
   U7843 : AOI22_X1 port map( A1 => n7068, A2 => n7067, B1 => intadd_0xSUMx23x,
                           B2 => n7270, ZN => n7072);
   U7844 : OAI22_X1 port map( A1 => n7076, A2 => n7223, B1 => n7477, B2 => 
                           n7394, ZN => n7069);
   U7845 : AOI21_X1 port map( B1 => n7070, B2 => n7406, A => n7069, ZN => n7071
                           );
   U7846 : OAI211_X1 port map( C1 => n7112, C2 => n7073, A => n7072, B => n7071
                           , ZN => n7106);
   U7847 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn94, A2 => n7364, ZN 
                           => n7104);
   U7848 : OAI22_X1 port map( A1 => n7075, A2 => n7308, B1 => n7074, B2 => 
                           n7188, ZN => n7102);
   U7849 : OAI221_X1 port map( B1 => n7076, B2 => n7315, C1 => add_x_26xBx25x, 
                           C2 => n7316, A => ashr_25xAx25x, ZN => n7077);
   U7850 : OAI21_X1 port map( B1 => n7216, B2 => n7078, A => n7077, ZN => n7101
                           );
   U7851 : AOI21_X1 port map( B1 => n7081, B2 => n7080, A => n7079, ZN => n7100
                           );
   U7852 : AOI22_X1 port map( A1 => n7205, A2 => n7122, B1 => intadd_1xAx7x, B2
                           => n7395, ZN => n7163);
   U7853 : AOI22_X1 port map( A1 => n7164, A2 => n7163, B1 => n7083, B2 => 
                           n7082, ZN => n7268);
   U7854 : OAI22_X1 port map( A1 => n7084, A2 => n7402, B1 => n7268, B2 => 
                           n7262, ZN => n7086);
   U7855 : AOI22_X1 port map( A1 => n7405, A2 => n7086, B1 => n7348, B2 => 
                           n7085, ZN => n7098);
   U7856 : AOI22_X1 port map( A1 => n7329, A2 => ashr_25xAx25x, B1 => 
                           ashr_25xAx24x, B2 => n7408, ZN => n7174);
   U7857 : INV_X1 port map( A => n7174, ZN => n7088);
   U7858 : AOI22_X1 port map( A1 => n7414, A2 => n7088, B1 => n7087, B2 => 
                           n7412, ZN => n7253);
   U7859 : OAI22_X1 port map( A1 => n7089, A2 => n7126, B1 => n7253, B2 => 
                           n7411, ZN => n7091);
   U7860 : AOI22_X1 port map( A1 => n7416, A2 => n7091, B1 => n7344, B2 => 
                           n7090, ZN => n7097);
   U7861 : INV_X1 port map( A => n7092, ZN => n7095);
   U7862 : OAI221_X1 port map( B1 => n7477, B2 => n7385, C1 => n7093, C2 => 
                           n7313, A => n7383, ZN => n7094);
   U7863 : AOI22_X1 port map( A1 => n7130, A2 => n7095, B1 => n7094, B2 => 
                           ashr_25xAx25x, ZN => n7096);
   U7864 : NAND4_X1 port map( A1 => n7098, A2 => n7097, A3 => n7157, A4 => 
                           n7096, ZN => n7099);
   U7865 : NOR4_X1 port map( A1 => n7102, A2 => n7101, A3 => n7100, A4 => n7099
                           , ZN => n7103);
   U7866 : NAND2_X1 port map( A1 => n7104, A2 => n7103, ZN => n7105);
   U7867 : AOI211_X1 port map( C1 => n7427, C2 => n7107, A => n7106, B => n7105
                           , ZN => n7109);
   U7868 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(25), ZN => n7108);
   U7869 : OAI22_X1 port map( A1 => n7109, A2 => n7529, B1 => n7108, B2 => 
                           n7435, ZN => IF_ISAxN10962);
   U7870 : OAI221_X1 port map( B1 => n7478, B2 => n7385, C1 => n7114, C2 => 
                           n7313, A => n7383, ZN => n7110);
   U7871 : AOI221_X1 port map( B1 => n7406, B2 => n7120, C1 => n7315, C2 => 
                           add_x_26xBx26x, A => n7110, ZN => n7113);
   U7872 : OAI22_X1 port map( A1 => n7162, A2 => n7113, B1 => n7112, B2 => 
                           n7111, ZN => n7151);
   U7873 : OAI211_X1 port map( C1 => n7318, C2 => n7323, A => n7162, B => n7114
                           , ZN => n7117);
   U7874 : OAI21_X1 port map( B1 => n7345, B2 => n7115, A => n7349, ZN => n7116
                           );
   U7875 : OAI211_X1 port map( C1 => n7120, C2 => n7223, A => n7117, B => n7116
                           , ZN => n7150);
   U7876 : OAI22_X1 port map( A1 => n7119, A2 => n7308, B1 => n7118, B2 => 
                           n7188, ZN => n7149);
   U7877 : NOR2_X1 port map( A1 => n7120, A2 => ashr_25xAx26x, ZN => n7121);
   U7878 : AOI22_X1 port map( A1 => intadd_0xSUMx24x, A2 => n7270, B1 => n7121,
                           B2 => n7406, ZN => n7145);
   U7879 : OAI22_X1 port map( A1 => n7123, A2 => n7162, B1 => n7122, B2 => 
                           n7410, ZN => n7226);
   U7880 : OAI22_X1 port map( A1 => n7125, A2 => n7226, B1 => n7124, B2 => 
                           n7414, ZN => n7334);
   U7881 : OAI22_X1 port map( A1 => n7334, A2 => n7411, B1 => n7127, B2 => 
                           n7126, ZN => n7128);
   U7882 : AOI22_X1 port map( A1 => n7130, A2 => n7129, B1 => n7416, B2 => 
                           n7128, ZN => n7144);
   U7883 : INV_X1 port map( A => n7131, ZN => n7132);
   U7884 : AOI21_X1 port map( B1 => n7427, B2 => n7132, A => n7283, ZN => n7143
                           );
   U7885 : AOI22_X1 port map( A1 => n7348, A2 => n7134, B1 => n7344, B2 => 
                           n7133, ZN => n7135);
   U7886 : INV_X1 port map( A => n7135, ZN => n7141);
   U7887 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx26x, B1 => 
                           ashr_25xAx25x, B2 => n7161, ZN => n7206);
   U7888 : AOI22_X1 port map( A1 => n7164, A2 => n7206, B1 => n7136, B2 => 
                           n7263, ZN => n7304);
   U7889 : AOI22_X1 port map( A1 => n7269, A2 => n7137, B1 => n7397, B2 => 
                           n7304, ZN => n7139);
   U7890 : OAI22_X1 port map( A1 => n7139, A2 => n7202, B1 => n7216, B2 => 
                           n7138, ZN => n7140);
   U7891 : NOR2_X1 port map( A1 => n7141, A2 => n7140, ZN => n7142);
   U7892 : NAND4_X1 port map( A1 => n7145, A2 => n7144, A3 => n7143, A4 => 
                           n7142, ZN => n7146);
   U7893 : AOI21_X1 port map( B1 => DP_OP_719J1_125_1055xn95, B2 => n7172, A =>
                           n7146, ZN => n7147);
   U7894 : INV_X1 port map( A => n7147, ZN => n7148);
   U7895 : NOR4_X1 port map( A1 => n7151, A2 => n7150, A3 => n7149, A4 => n7148
                           , ZN => n7153);
   U7896 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(26), ZN => n7152);
   U7897 : OAI22_X1 port map( A1 => n7153, A2 => n7529, B1 => n7152, B2 => 
                           n7435, ZN => IF_ISAxN10963);
   U7898 : AOI22_X1 port map( A1 => n7179, A2 => n7248, B1 => add_x_26xBx27x, 
                           B2 => n7315, ZN => n7154);
   U7899 : AOI21_X1 port map( B1 => n7383, B2 => n7154, A => n7180, ZN => n7155
                           );
   U7900 : AOI21_X1 port map( B1 => n7318, B2 => n7179, A => n7155, ZN => n7156
                           );
   U7901 : OAI211_X1 port map( C1 => n7325, C2 => n7158, A => n7157, B => n7156
                           , ZN => n7171);
   U7902 : AOI22_X1 port map( A1 => n7160, A2 => n7159, B1 => add_x_26xBx27x, 
                           B2 => n7376, ZN => n7169);
   U7903 : AOI22_X1 port map( A1 => n7205, A2 => n7180, B1 => n7162, B2 => 
                           n7161, ZN => n7264);
   U7904 : AOI22_X1 port map( A1 => n7164, A2 => n7264, B1 => n7163, B2 => 
                           n7263, ZN => n7403);
   U7905 : OAI22_X1 port map( A1 => n7165, A2 => n7402, B1 => n7403, B2 => 
                           n7262, ZN => n7167);
   U7906 : AOI22_X1 port map( A1 => n7405, A2 => n7167, B1 => n7348, B2 => 
                           n7166, ZN => n7168);
   U7907 : NAND2_X1 port map( A1 => n7169, A2 => n7168, ZN => n7170);
   U7908 : AOI211_X1 port map( C1 => DP_OP_719J1_125_1055xn96, C2 => n7172, A 
                           => n7171, B => n7170, ZN => n7173);
   U7909 : INV_X1 port map( A => n7173, ZN => n7198);
   U7910 : AOI22_X1 port map( A1 => n7329, A2 => ashr_25xAx27x, B1 => 
                           ashr_25xAx26x, B2 => n7408, ZN => n7255);
   U7911 : AOI22_X1 port map( A1 => n7414, A2 => n7255, B1 => n7174, B2 => 
                           n7254, ZN => n7417);
   U7912 : INV_X1 port map( A => n7175, ZN => n7176);
   U7913 : AOI22_X1 port map( A1 => n7337, A2 => n7417, B1 => n7418, B2 => 
                           n7176, ZN => n7196);
   U7914 : OAI22_X1 port map( A1 => n7178, A2 => n7310, B1 => n7177, B2 => 
                           n7393, ZN => n7184);
   U7915 : NAND2_X1 port map( A1 => n7180, A2 => n7179, ZN => n7182);
   U7916 : OAI22_X1 port map( A1 => n7182, A2 => n7393, B1 => n7181, B2 => 
                           n7380, ZN => n7183);
   U7917 : AOI211_X1 port map( C1 => n7344, C2 => n7185, A => n7184, B => n7183
                           , ZN => n7195);
   U7918 : OAI21_X1 port map( B1 => n7345, B2 => n7186, A => n7349, ZN => n7187
                           );
   U7919 : INV_X1 port map( A => n7187, ZN => n7192);
   U7920 : OAI22_X1 port map( A1 => n7190, A2 => n7308, B1 => n7189, B2 => 
                           n7188, ZN => n7191);
   U7921 : AOI211_X1 port map( C1 => n7427, C2 => n7193, A => n7192, B => n7191
                           , ZN => n7194);
   U7922 : OAI211_X1 port map( C1 => n7196, C2 => n7339, A => n7195, B => n7194
                           , ZN => n7197);
   U7923 : AOI211_X1 port map( C1 => n7199, C2 => n7443, A => n7198, B => n7197
                           , ZN => n7201);
   U7924 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(27), ZN => n7200);
   U7925 : OAI22_X1 port map( A1 => n7201, A2 => n7529, B1 => n7200, B2 => 
                           n7435, ZN => IF_ISAxN10964);
   U7926 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn97, A2 => n7364, ZN 
                           => n7215);
   U7927 : AOI21_X1 port map( B1 => n7204, B2 => n7203, A => n7202, ZN => n7208
                           );
   U7928 : AOI22_X1 port map( A1 => n7205, A2 => ashr_25xAx28x, B1 => 
                           ashr_25xAx27x, B2 => n7395, ZN => n7295);
   U7929 : OAI221_X1 port map( B1 => n6586, B2 => n7206, C1 => n7399, C2 => 
                           n7295, A => n7397, ZN => n7207);
   U7930 : OAI211_X1 port map( C1 => n7402, C2 => n7209, A => n7208, B => n7207
                           , ZN => n7214);
   U7931 : INV_X1 port map( A => n7210, ZN => n7211);
   U7932 : AOI22_X1 port map( A1 => n7344, A2 => n7212, B1 => n7348, B2 => 
                           n7211, ZN => n7213);
   U7933 : NAND3_X1 port map( A1 => n7215, A2 => n7214, A3 => n7213, ZN => 
                           n7242);
   U7934 : NOR2_X1 port map( A1 => n7411, A2 => n7216, ZN => n7391);
   U7935 : INV_X1 port map( A => n7391, ZN => n7279);
   U7936 : AOI21_X1 port map( B1 => n7327, B2 => n7217, A => n7325, ZN => n7222
                           );
   U7937 : OAI221_X1 port map( B1 => n7480, B2 => n7385, C1 => n7237, C2 => 
                           n7313, A => n7383, ZN => n7218);
   U7938 : AOI221_X1 port map( B1 => n7406, B2 => intadd_3xBx0x, C1 => n7315, 
                           C2 => add_x_26xBx28x, A => n7218, ZN => n7220);
   U7939 : NAND2_X1 port map( A1 => intadd_3xAx0x, A2 => n7237, ZN => n7219);
   U7940 : OAI22_X1 port map( A1 => intadd_3xAx0x, A2 => n7220, B1 => n7393, B2
                           => n7219, ZN => n7221);
   U7941 : AOI211_X1 port map( C1 => n7270, C2 => intadd_0xSUMx26x, A => n7222,
                           B => n7221, ZN => n7239);
   U7942 : AOI221_X1 port map( B1 => ashr_25xAx28x, B2 => n7223, C1 => n7310, 
                           C2 => n7223, A => intadd_3xBx0x, ZN => n7236);
   U7943 : OAI21_X1 port map( B1 => n7345, B2 => n7224, A => n7349, ZN => n7233
                           );
   U7944 : AOI21_X1 port map( B1 => n7418, B2 => n7225, A => n7339, ZN => n7229
                           );
   U7945 : INV_X1 port map( A => n7226, ZN => n7227);
   U7946 : AOI22_X1 port map( A1 => n7329, A2 => ashr_25xAx28x, B1 => 
                           ashr_25xAx27x, B2 => n7408, ZN => n7328);
   U7947 : OAI221_X1 port map( B1 => n7414, B2 => n7227, C1 => n7412, C2 => 
                           n7328, A => n7337, ZN => n7228);
   U7948 : OAI211_X1 port map( C1 => n7231, C2 => n7230, A => n7229, B => n7228
                           , ZN => n7232);
   U7949 : OAI211_X1 port map( C1 => n7234, C2 => n7423, A => n7233, B => n7232
                           , ZN => n7235);
   U7950 : AOI211_X1 port map( C1 => n7318, C2 => n7237, A => n7236, B => n7235
                           , ZN => n7238);
   U7951 : OAI211_X1 port map( C1 => n7240, C2 => n7279, A => n7239, B => n7238
                           , ZN => n7241);
   U7952 : AOI211_X1 port map( C1 => n7243, C2 => n7443, A => n7242, B => n7241
                           , ZN => n7245);
   U7953 : OAI22_X1 port map( A1 => n7245, A2 => n7529, B1 => n7244, B2 => 
                           n7435, ZN => IF_ISAxN10965);
   U7954 : NAND2_X1 port map( A1 => intadd_3xAx1x, A2 => n7247, ZN => n7261);
   U7955 : AOI221_X1 port map( B1 => n7323, B2 => n7481, C1 => n7248, C2 => 
                           n7247, A => n7246, ZN => n7249);
   U7956 : OAI221_X1 port map( B1 => intadd_3xBx1x, B2 => n7382, C1 => 
                           add_x_26xBx29x, C2 => n7250, A => n7249, ZN => n7251
                           );
   U7957 : AOI22_X1 port map( A1 => n7406, A2 => n7252, B1 => ashr_25xAx29x, B2
                           => n7251, ZN => n7260);
   U7958 : AOI21_X1 port map( B1 => n7418, B2 => n7253, A => n7339, ZN => n7257
                           );
   U7959 : AOI22_X1 port map( A1 => n7329, A2 => ashr_25xAx29x, B1 => 
                           ashr_25xAx28x, B2 => n7123, ZN => n7413);
   U7960 : OAI221_X1 port map( B1 => n7414, B2 => n7255, C1 => n7254, C2 => 
                           n7413, A => n7337, ZN => n7256);
   U7961 : OAI211_X1 port map( C1 => intadd_4xBx2x, C2 => n7258, A => n7257, B 
                           => n7256, ZN => n7259);
   U7962 : OAI211_X1 port map( C1 => n7393, C2 => n7261, A => n7260, B => n7259
                           , ZN => n7289);
   U7963 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn98, A2 => n7364, ZN 
                           => n7287);
   U7964 : AOI22_X1 port map( A1 => n7205, A2 => intadd_3xAx1x, B1 => 
                           intadd_3xAx0x, B2 => n7296, ZN => n7400);
   U7965 : AOI221_X1 port map( B1 => n7400, B2 => n7164, C1 => n7264, C2 => 
                           n7263, A => n7262, ZN => n7267);
   U7966 : OAI21_X1 port map( B1 => n7372, B2 => n7265, A => n7405, ZN => n7266
                           );
   U7967 : AOI211_X1 port map( C1 => n7269, C2 => n7268, A => n7267, B => n7266
                           , ZN => n7275);
   U7968 : AOI22_X1 port map( A1 => intadd_0xSUMx27x, A2 => n7270, B1 => 
                           add_x_26xBx29x, B2 => n7376, ZN => n7273);
   U7969 : OAI21_X1 port map( B1 => n7345, B2 => n7271, A => n7349, ZN => n7272
                           );
   U7970 : OAI211_X1 port map( C1 => n7481, C2 => n7394, A => n7273, B => n7272
                           , ZN => n7274);
   U7971 : AOI211_X1 port map( C1 => n7344, C2 => n7276, A => n7275, B => n7274
                           , ZN => n7286);
   U7972 : OAI22_X1 port map( A1 => n7423, A2 => n7278, B1 => n7366, B2 => 
                           n7277, ZN => n7284);
   U7973 : OAI22_X1 port map( A1 => n7325, A2 => n7281, B1 => n7280, B2 => 
                           n7279, ZN => n7282);
   U7974 : NOR3_X1 port map( A1 => n7284, A2 => n7283, A3 => n7282, ZN => n7285
                           );
   U7975 : NAND3_X1 port map( A1 => n7287, A2 => n7286, A3 => n7285, ZN => 
                           n7288);
   U7976 : AOI211_X1 port map( C1 => n7290, C2 => n7443, A => n7289, B => n7288
                           , ZN => n7292);
   U7977 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(29), ZN => n7291);
   U7978 : OAI22_X1 port map( A1 => n7292, A2 => n7529, B1 => n7291, B2 => 
                           n7435, ZN => IF_ISAxN10966);
   U7979 : AOI22_X1 port map( A1 => n7391, A2 => n7294, B1 => n7427, B2 => 
                           n7293, ZN => n7307);
   U7980 : INV_X1 port map( A => n7295, ZN => n7300);
   U7981 : NOR2_X1 port map( A1 => n7296, A2 => ashr_25xAx30x, ZN => n7298);
   U7982 : NOR2_X1 port map( A1 => n7396, A2 => ashr_25xAx29x, ZN => n7297);
   U7983 : NOR2_X1 port map( A1 => n7298, A2 => n7297, ZN => n7299);
   U7984 : MUX2_X1 port map( A => n7300, B => n7299, S => n6586, Z => n7302);
   U7985 : OAI221_X1 port map( B1 => n7305, B2 => n7304, C1 => n7303, C2 => 
                           n7302, A => n7301, ZN => n7306);
   U7986 : OAI211_X1 port map( C1 => n7309, C2 => n7308, A => n7307, B => n7306
                           , ZN => n7356);
   U7987 : NAND2_X1 port map( A1 => DP_OP_719J1_125_1055xn99, A2 => n7364, ZN 
                           => n7354);
   U7988 : INV_X1 port map( A => intadd_0xSUMx28x, ZN => n7312);
   U7989 : OAI22_X1 port map( A1 => n7312, A2 => n7380, B1 => n7311, B2 => 
                           n7310, ZN => n7322);
   U7990 : OAI221_X1 port map( B1 => n7483, B2 => n7385, C1 => n7317, C2 => 
                           n7313, A => n7383, ZN => n7314);
   U7991 : AOI221_X1 port map( B1 => n7316, B2 => intadd_3xBx2x, C1 => n7315, 
                           C2 => add_x_26xBx30x, A => n7314, ZN => n7320);
   U7992 : AOI22_X1 port map( A1 => n7318, A2 => n7317, B1 => add_x_26xBx30x, 
                           B2 => n7376, ZN => n7319);
   U7993 : OAI21_X1 port map( B1 => intadd_3xAx2x, B2 => n7320, A => n7319, ZN 
                           => n7321);
   U7994 : AOI211_X1 port map( C1 => n7324, C2 => n7323, A => n7322, B => n7321
                           , ZN => n7353);
   U7995 : AOI21_X1 port map( B1 => n7327, B2 => n7326, A => n7325, ZN => n7342
                           );
   U7996 : INV_X1 port map( A => n7328, ZN => n7333);
   U7997 : NOR2_X1 port map( A1 => ashr_25xAx30x, A2 => n7123, ZN => n7331);
   U7998 : NOR2_X1 port map( A1 => n7329, A2 => ashr_25xAx29x, ZN => n7330);
   U7999 : NOR2_X1 port map( A1 => n7331, A2 => n7330, ZN => n7332);
   U8000 : MUX2_X1 port map( A => n7333, B => n7332, S => n7414, Z => n7336);
   U8001 : INV_X1 port map( A => n7334, ZN => n7335);
   U8002 : AOI22_X1 port map( A1 => n7337, A2 => n7336, B1 => n7418, B2 => 
                           n7335, ZN => n7340);
   U8003 : OAI22_X1 port map( A1 => n7340, A2 => n7339, B1 => n7423, B2 => 
                           n7338, ZN => n7341);
   U8004 : AOI211_X1 port map( C1 => n7344, C2 => n7343, A => n7342, B => n7341
                           , ZN => n7352);
   U8005 : OR2_X1 port map( A1 => n7346, A2 => n7345, ZN => n7350);
   U8006 : AOI22_X1 port map( A1 => n7350, A2 => n7349, B1 => n7348, B2 => 
                           n7347, ZN => n7351);
   U8007 : NAND4_X1 port map( A1 => n7354, A2 => n7353, A3 => n7352, A4 => 
                           n7351, ZN => n7355);
   U8008 : AOI211_X1 port map( C1 => n7357, C2 => n7443, A => n7356, B => n7355
                           , ZN => n7359);
   U8009 : OAI22_X1 port map( A1 => n7359, A2 => n7529, B1 => n7358, B2 => 
                           n7435, ZN => IF_ISAxN10967);
   U8010 : OAI21_X1 port map( B1 => n7360, B2 => n7485, A => n7388, ZN => n7361
                           );
   U8011 : XOR2_X1 port map( A => n7546, B => n7361, Z => n7362);
   U8012 : XOR2_X1 port map( A => n7362, B => n7409, Z => n7363);
   U8013 : XOR2_X1 port map( A => DP_OP_719J1_125_1055xn2, B => n7363, Z => 
                           n7365);
   U8014 : NAND2_X1 port map( A1 => n7365, A2 => n7364, ZN => n7378);
   U8015 : NOR2_X1 port map( A1 => n7367, A2 => n7366, ZN => n7374);
   U8016 : NOR2_X1 port map( A1 => n7368, A2 => n7372, ZN => n7370);
   U8017 : AOI211_X1 port map( C1 => n7372, C2 => n7371, A => n7370, B => n7369
                           , ZN => n7373);
   U8018 : AOI211_X1 port map( C1 => n7376, C2 => n7375, A => n7374, B => n7373
                           , ZN => n7377);
   U8019 : OAI211_X1 port map( C1 => n7380, C2 => n7379, A => n7378, B => n7377
                           , ZN => n7433);
   U8020 : OAI21_X1 port map( B1 => n7388, B2 => n7382, A => n7381, ZN => n7387
                           );
   U8021 : OAI221_X1 port map( B1 => n7485, B2 => n7385, C1 => n7384, C2 => 
                           n7393, A => n7383, ZN => n7386);
   U8022 : AOI211_X1 port map( C1 => n7406, C2 => n7388, A => n7387, B => n7386
                           , ZN => n7430);
   U8023 : AOI22_X1 port map( A1 => n7392, A2 => n7391, B1 => n7390, B2 => 
                           n7389, ZN => n7429);
   U8024 : AOI211_X1 port map( C1 => n7394, C2 => n7393, A => n7409, B => n7485
                           , ZN => n7425);
   U8025 : AOI22_X1 port map( A1 => n7396, A2 => n7431, B1 => intadd_3xAx2x, B2
                           => n7395, ZN => n7398);
   U8026 : OAI221_X1 port map( B1 => n7164, B2 => n7400, C1 => n7399, C2 => 
                           n7398, A => n7397, ZN => n7401);
   U8027 : OAI21_X1 port map( B1 => n7403, B2 => n7402, A => n7401, ZN => n7404
                           );
   U8028 : AOI22_X1 port map( A1 => n7407, A2 => n7406, B1 => n7405, B2 => 
                           n7404, ZN => n7421);
   U8029 : AOI22_X1 port map( A1 => n7410, A2 => n7409, B1 => ashr_25xAx30x, B2
                           => n7408, ZN => n7415);
   U8030 : AOI221_X1 port map( B1 => n7415, B2 => n7414, C1 => n7413, C2 => 
                           n7412, A => n7411, ZN => n7419);
   U8031 : OAI221_X1 port map( B1 => n7419, B2 => n7418, C1 => n7419, C2 => 
                           n7417, A => n7416, ZN => n7420);
   U8032 : OAI211_X1 port map( C1 => n7423, C2 => n7422, A => n7421, B => n7420
                           , ZN => n7424);
   U8033 : AOI211_X1 port map( C1 => n7427, C2 => n7426, A => n7425, B => n7424
                           , ZN => n7428);
   U8034 : OAI211_X1 port map( C1 => n7431, C2 => n7430, A => n7429, B => n7428
                           , ZN => n7432);
   U8035 : AOI211_X1 port map( C1 => n7434, C2 => n7443, A => n7433, B => n7432
                           , ZN => n7437);
   U8036 : OAI22_X1 port map( A1 => n7437, A2 => n7529, B1 => n7436, B2 => 
                           n7435, ZN => IF_ISAxN10968);
   U8037 : NOR2_X1 port map( A1 => rst, A2 => n7438, ZN => IF_ISAxN10970);
   U8038 : NOR2_X1 port map( A1 => rst, A2 => n7439, ZN => IF_ISAxN10971);
   U8039 : AND2_X1 port map( A1 => n7505, A2 => fromMemoryPortxLOADEDDATAx(9), 
                           ZN => IF_ISAxN10972);
   U8040 : AND2_X1 port map( A1 => n7505, A2 => fromMemoryPortxLOADEDDATAx(10),
                           ZN => IF_ISAxN10973);
   U8041 : AND2_X1 port map( A1 => n7519, A2 => fromMemoryPortxLOADEDDATAx(11),
                           ZN => IF_ISAxN10974);
   U8042 : NAND3_X1 port map( A1 => n7534, A2 => n7531, A3 => n7451, ZN => 
                           n7488);
   U8043 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(2), A2 => 
                           fromMemoryPortxLOADEDDATAx(4), ZN => n7447);
   U8044 : INV_X1 port map( A => n7488, ZN => n7446);
   U8045 : NOR3_X1 port map( A1 => n7442, A2 => n7441, A3 => n7440, ZN => n7444
                           );
   U8046 : NAND2_X1 port map( A1 => n7444, A2 => n7443, ZN => n7445);
   U8047 : NAND2_X1 port map( A1 => n7446, A2 => n7445, ZN => n7487);
   U8048 : NOR2_X1 port map( A1 => n7447, A2 => n7487, ZN => n7452);
   U8049 : NOR2_X1 port map( A1 => rst, A2 => n7452, ZN => n7523);
   U8050 : OAI21_X1 port map( B1 => n7448, B2 => n7488, A => n7523, ZN => 
                           IF_ISAxN10969);
   U8051 : INV_X1 port map( A => n7449, ZN => n7450);
   U8052 : AOI21_X1 port map( B1 => n7451, B2 => n7450, A => rst, ZN => n7489);
   U8053 : INV_X1 port map( A => n7452, ZN => n7528);
   U8054 : OAI211_X1 port map( C1 => n7453, C2 => n7488, A => n7489, B => n7528
                           , ZN => IF_ISAxN10902);
   U8055 : NAND2_X1 port map( A1 => n7454, A2 => IF_ISAxsection_0_port, ZN => 
                           n7455);
   U8056 : NAND3_X1 port map( A1 => n7456, A2 => n7489, A3 => n7455, ZN => 
                           n7484);
   U8057 : CLKBUF_X1 port map( A => n7484, Z => n7482);
   U8058 : NOR2_X1 port map( A1 => n7457, A2 => n7482, ZN => IF_ISAxN10842);
   U8059 : NOR2_X1 port map( A1 => n7458, A2 => n7482, ZN => IF_ISAxN10843);
   U8060 : NOR2_X1 port map( A1 => n7459, A2 => n7482, ZN => IF_ISAxN10844);
   U8061 : NOR2_X1 port map( A1 => n7460, A2 => n7482, ZN => IF_ISAxN10845);
   U8062 : NOR2_X1 port map( A1 => n7461, A2 => n7482, ZN => IF_ISAxN10846);
   U8063 : NOR2_X1 port map( A1 => n7462, A2 => n7482, ZN => IF_ISAxN10847);
   U8064 : NOR2_X1 port map( A1 => n7463, A2 => n7482, ZN => IF_ISAxN10848);
   U8065 : NOR2_X1 port map( A1 => n7464, A2 => n7482, ZN => IF_ISAxN10849);
   U8066 : NOR2_X1 port map( A1 => n7465, A2 => n7482, ZN => IF_ISAxN10850);
   U8067 : NOR2_X1 port map( A1 => n7466, A2 => n7482, ZN => IF_ISAxN10851);
   U8068 : NOR2_X1 port map( A1 => n7467, A2 => n7482, ZN => IF_ISAxN10852);
   U8069 : NOR2_X1 port map( A1 => n7468, A2 => n7482, ZN => IF_ISAxN10853);
   U8070 : NOR2_X1 port map( A1 => n7469, A2 => n7484, ZN => IF_ISAxN10854);
   U8071 : NOR2_X1 port map( A1 => n7470, A2 => n7484, ZN => IF_ISAxN10855);
   U8072 : NOR2_X1 port map( A1 => n7471, A2 => n7484, ZN => IF_ISAxN10856);
   U8073 : NOR2_X1 port map( A1 => n7472, A2 => n7484, ZN => IF_ISAxN10857);
   U8074 : NOR2_X1 port map( A1 => n7473, A2 => n7484, ZN => IF_ISAxN10858);
   U8075 : NOR2_X1 port map( A1 => n7474, A2 => n7484, ZN => IF_ISAxN10859);
   U8076 : NOR2_X1 port map( A1 => n7475, A2 => n7484, ZN => IF_ISAxN10860);
   U8077 : NOR2_X1 port map( A1 => n7476, A2 => n7484, ZN => IF_ISAxN10861);
   U8078 : NOR2_X1 port map( A1 => n7477, A2 => n7484, ZN => IF_ISAxN10862);
   U8079 : NOR2_X1 port map( A1 => n7478, A2 => n7484, ZN => IF_ISAxN10863);
   U8080 : NOR2_X1 port map( A1 => n7479, A2 => n7484, ZN => IF_ISAxN10864);
   U8081 : NOR2_X1 port map( A1 => n7480, A2 => n7482, ZN => IF_ISAxN10865);
   U8082 : NOR2_X1 port map( A1 => n7481, A2 => n7484, ZN => IF_ISAxN10866);
   U8083 : NOR2_X1 port map( A1 => n7483, A2 => n7482, ZN => IF_ISAxN10867);
   U8084 : NOR2_X1 port map( A1 => n7485, A2 => n7484, ZN => IF_ISAxN10868);
   U8085 : OAI21_X1 port map( B1 => n7486, B2 => n7488, A => n7489, ZN => 
                           IF_ISAxN10832);
   U8086 : NAND2_X1 port map( A1 => n7489, A2 => n7487, ZN => IF_ISAxN10869);
   U8087 : OAI21_X1 port map( B1 => n7534, B2 => n7531, A => 
                           toMemoryPort_sync_port, ZN => n7490);
   U8088 : OAI211_X1 port map( C1 => IF_ISAxsection_0_port, C2 => n7490, A => 
                           n7489, B => n7488, ZN => IF_ISAxN10829);
   U8089 : NAND2_X1 port map( A1 => toRegsPortxDSTxx3x, A2 => 
                           toRegsPortxDSTxx2x, ZN => n7492);
   U8090 : NOR2_X1 port map( A1 => n7530, A2 => n7492, ZN => n7504);
   U8091 : INV_X1 port map( A => n7504, ZN => n7491);
   U8092 : NAND2_X1 port map( A1 => toRegsPortxDSTxx0x, A2 => 
                           toRegsPortxDSTxx4x, ZN => n7502);
   U8093 : OR2_X1 port map( A1 => n7536, A2 => n7502, ZN => n7493);
   U8094 : OAI21_X1 port map( B1 => n7491, B2 => n7493, A => n7505, ZN => 
                           IF_RegsxN659);
   U8095 : NAND2_X1 port map( A1 => toRegsPortxDSTxx4x, A2 => n7532, ZN => 
                           n7503);
   U8096 : OR2_X1 port map( A1 => n7536, A2 => n7503, ZN => n7501);
   U8097 : OAI21_X1 port map( B1 => n7491, B2 => n7501, A => n7516, ZN => 
                           IF_RegsxN692);
   U8098 : NOR2_X1 port map( A1 => toRegsPortxDSTxx1x, A2 => n7492, ZN => n7507
                           );
   U8099 : INV_X1 port map( A => n7507, ZN => n7494);
   U8100 : OAI21_X1 port map( B1 => n7494, B2 => n7493, A => n7519, ZN => 
                           IF_RegsxN693);
   U8101 : OAI21_X1 port map( B1 => n7494, B2 => n7501, A => n7516, ZN => 
                           IF_RegsxN694);
   U8102 : NAND4_X1 port map( A1 => toRegsPortxDSTxx1x, A2 => toRegsPort_notify
                           , A3 => toRegsPortxDSTxx3x, A4 => n7533, ZN => n7509
                           );
   U8103 : OAI21_X1 port map( B1 => n7502, B2 => n7509, A => n7505, ZN => 
                           IF_RegsxN695);
   U8104 : OAI21_X1 port map( B1 => n7503, B2 => n7509, A => n7519, ZN => 
                           IF_RegsxN696);
   U8105 : NAND2_X1 port map( A1 => toRegsPort_notify, A2 => toRegsPortxDSTxx0x
                           , ZN => n7499);
   U8106 : OAI21_X1 port map( B1 => n7499, B2 => n7495, A => n7519, ZN => 
                           IF_RegsxN697);
   U8107 : NAND2_X1 port map( A1 => toRegsPortxDSTxx2x, A2 => n7537, ZN => 
                           n7497);
   U8108 : NOR2_X1 port map( A1 => n7530, A2 => n7497, ZN => n7511);
   U8109 : NAND2_X1 port map( A1 => toRegsPort_notify, A2 => n7511, ZN => n7496
                           );
   U8110 : OAI21_X1 port map( B1 => n7502, B2 => n7496, A => n7505, ZN => 
                           IF_RegsxN699);
   U8111 : OAI21_X1 port map( B1 => n7496, B2 => n7503, A => n7505, ZN => 
                           IF_RegsxN700);
   U8112 : NOR2_X1 port map( A1 => toRegsPortxDSTxx1x, A2 => n7497, ZN => n7500
                           );
   U8113 : NAND2_X1 port map( A1 => toRegsPortxDSTxx4x, A2 => n7500, ZN => 
                           n7498);
   U8114 : OAI21_X1 port map( B1 => n7499, B2 => n7498, A => n7505, ZN => 
                           IF_RegsxN701);
   U8115 : INV_X1 port map( A => n7500, ZN => n7515);
   U8116 : OAI21_X1 port map( B1 => n7501, B2 => n7515, A => n7516, ZN => 
                           IF_RegsxN702);
   U8117 : NAND4_X1 port map( A1 => toRegsPortxDSTxx1x, A2 => toRegsPort_notify
                           , A3 => n7537, A4 => n7533, ZN => n7518);
   U8118 : OAI21_X1 port map( B1 => n7502, B2 => n7518, A => n7516, ZN => 
                           IF_RegsxN703);
   U8119 : OAI21_X1 port map( B1 => n7503, B2 => n7518, A => n7505, ZN => 
                           IF_RegsxN704);
   U8120 : NAND4_X1 port map( A1 => toRegsPort_notify, A2 => n7537, A3 => n7530
                           , A4 => n7533, ZN => n7521);
   U8121 : OAI21_X1 port map( B1 => n7502, B2 => n7521, A => n7516, ZN => 
                           IF_RegsxN705);
   U8122 : OAI21_X1 port map( B1 => n7503, B2 => n7521, A => n7519, ZN => 
                           IF_RegsxN706);
   U8123 : NAND3_X1 port map( A1 => toRegsPort_notify, A2 => n7504, A3 => n7535
                           , ZN => n7506);
   U8124 : OAI21_X1 port map( B1 => n7532, B2 => n7506, A => n7505, ZN => 
                           IF_RegsxN707);
   U8125 : OAI21_X1 port map( B1 => toRegsPortxDSTxx0x, B2 => n7506, A => n7516
                           , ZN => IF_RegsxN708);
   U8126 : NAND3_X1 port map( A1 => toRegsPort_notify, A2 => n7507, A3 => n7535
                           , ZN => n7508);
   U8127 : OAI21_X1 port map( B1 => n7532, B2 => n7508, A => n7516, ZN => 
                           IF_RegsxN709);
   U8128 : OAI21_X1 port map( B1 => toRegsPortxDSTxx0x, B2 => n7508, A => n7516
                           , ZN => IF_RegsxN710);
   U8129 : NAND2_X1 port map( A1 => toRegsPortxDSTxx0x, A2 => n7535, ZN => 
                           n7520);
   U8130 : OAI21_X1 port map( B1 => n7509, B2 => n7520, A => n7519, ZN => 
                           IF_RegsxN711);
   U8131 : NAND2_X1 port map( A1 => n7532, A2 => n7535, ZN => n7517);
   U8132 : OAI21_X1 port map( B1 => n7509, B2 => n7517, A => n7516, ZN => 
                           IF_RegsxN712);
   U8133 : OR2_X1 port map( A1 => n7536, A2 => n7520, ZN => n7513);
   U8134 : OAI21_X1 port map( B1 => n7510, B2 => n7513, A => n7516, ZN => 
                           IF_RegsxN713);
   U8135 : OR2_X1 port map( A1 => n7536, A2 => n7517, ZN => n7514);
   U8136 : OAI21_X1 port map( B1 => n7510, B2 => n7514, A => n7516, ZN => 
                           IF_RegsxN714);
   U8137 : INV_X1 port map( A => n7511, ZN => n7512);
   U8138 : OAI21_X1 port map( B1 => n7512, B2 => n7513, A => n7516, ZN => 
                           IF_RegsxN715);
   U8139 : OAI21_X1 port map( B1 => n7512, B2 => n7514, A => n7516, ZN => 
                           IF_RegsxN716);
   U8140 : OAI21_X1 port map( B1 => n7515, B2 => n7513, A => n7516, ZN => 
                           IF_RegsxN717);
   U8141 : OAI21_X1 port map( B1 => n7515, B2 => n7514, A => n7516, ZN => 
                           IF_RegsxN718);
   U8142 : OAI21_X1 port map( B1 => n7518, B2 => n7520, A => n7516, ZN => 
                           IF_RegsxN719);
   U8143 : OAI21_X1 port map( B1 => n7518, B2 => n7517, A => n7516, ZN => 
                           IF_RegsxN720);
   U8144 : OAI21_X1 port map( B1 => n7521, B2 => n7520, A => n7519, ZN => 
                           IF_RegsxN721);
   U8145 : NAND2_X1 port map( A1 => n7523, A2 => n7522, ZN => IF_ISAxN10935);
   U8146 : NAND2_X1 port map( A1 => n7534, A2 => n7531, ZN => n7525);
   U8147 : INV_X1 port map( A => IF_ISAxN10935, ZN => n7524);
   U8148 : OAI211_X1 port map( C1 => IF_ISAxsection_0_port, C2 => n7525, A => 
                           n7524, B => toRegsPort_notify, ZN => n7526);
   U8149 : OAI211_X1 port map( C1 => n7529, C2 => n7528, A => n7527, B => n7526
                           , ZN => n3458);
   clk_gate_IF_ISAxtoMemoryPort_notify_reg : SNPS_CLOCK_GATE_HIGH_CPU_0 port 
                           map( CLK => clk, EN => IF_ISAxN10829, ENCLK => 
                           net6523);
   clk_gate_IF_ISAxtoRegsPort_regxDSTDATAx : SNPS_CLOCK_GATE_HIGH_CPU_36 port 
                           map( CLK => clk, EN => IF_ISAxN10935, ENCLK => 
                           net6528);
   clk_gate_IF_ISAxtoRegsPort_regxDSTx : SNPS_CLOCK_GATE_HIGH_CPU_35 port map( 
                           CLK => clk, EN => IF_ISAxN10969, ENCLK => net6533);
   clk_gate_IF_ISAxpcReg_signal_reg : SNPS_CLOCK_GATE_HIGH_CPU_34 port map( CLK
                           => clk, EN => IF_ISAxN10902, ENCLK => net6538);
   clk_gate_IF_ISAxtoMemoryPort_regxREQx : SNPS_CLOCK_GATE_HIGH_CPU_33 port 
                           map( CLK => clk, EN => IF_ISAxN10832, ENCLK => 
                           net6543);
   clk_gate_IF_ISAxtoMemoryPort_regxADDRINx : SNPS_CLOCK_GATE_HIGH_CPU_32 port 
                           map( CLK => clk, EN => IF_ISAxN10869, ENCLK => 
                           net6548);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_31x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_31 port map( CLK => clk, EN
                           => IF_RegsxN659, ENCLK => net6553);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_30x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_30 port map( CLK => clk, EN
                           => IF_RegsxN692, ENCLK => net6558);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_29x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_29 port map( CLK => clk, EN
                           => IF_RegsxN693, ENCLK => net6563);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_28x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_28 port map( CLK => clk, EN
                           => IF_RegsxN694, ENCLK => net6568);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_27x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_27 port map( CLK => clk, EN
                           => IF_RegsxN695, ENCLK => net6573);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_26x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_26 port map( CLK => clk, EN
                           => IF_RegsxN696, ENCLK => net6578);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_25x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_25 port map( CLK => clk, EN
                           => IF_RegsxN697, ENCLK => net6583);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_24x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_24 port map( CLK => clk, EN
                           => IF_RegsxN698, ENCLK => net6588);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_23x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_23 port map( CLK => clk, EN
                           => IF_RegsxN699, ENCLK => net6593);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_22x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_22 port map( CLK => clk, EN
                           => IF_RegsxN700, ENCLK => net6598);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_21x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_21 port map( CLK => clk, EN
                           => IF_RegsxN701, ENCLK => net6603);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_20x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_20 port map( CLK => clk, EN
                           => IF_RegsxN702, ENCLK => net6608);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_19x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_19 port map( CLK => clk, EN
                           => IF_RegsxN703, ENCLK => net6613);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_18x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_18 port map( CLK => clk, EN
                           => IF_RegsxN704, ENCLK => net6618);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_17x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_17 port map( CLK => clk, EN
                           => IF_RegsxN705, ENCLK => net6623);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_16x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_16 port map( CLK => clk, EN
                           => IF_RegsxN706, ENCLK => net6628);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_15x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_15 port map( CLK => clk, EN
                           => IF_RegsxN707, ENCLK => net6633);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_14x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_14 port map( CLK => clk, EN
                           => IF_RegsxN708, ENCLK => net6638);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_13x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_13 port map( CLK => clk, EN
                           => IF_RegsxN709, ENCLK => net6643);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_12x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_12 port map( CLK => clk, EN
                           => IF_RegsxN710, ENCLK => net6648);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_11x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_11 port map( CLK => clk, EN
                           => IF_RegsxN711, ENCLK => net6653);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_10x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_10 port map( CLK => clk, EN
                           => IF_RegsxN712, ENCLK => net6658);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_09x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_9 port map( CLK => clk, EN 
                           => IF_RegsxN713, ENCLK => net6663);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_08x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_8 port map( CLK => clk, EN 
                           => IF_RegsxN714, ENCLK => net6668);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_07x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_7 port map( CLK => clk, EN 
                           => IF_RegsxN715, ENCLK => net6673);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_06x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_6 port map( CLK => clk, EN 
                           => IF_RegsxN716, ENCLK => net6678);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_05x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_5 port map( CLK => clk, EN 
                           => IF_RegsxN717, ENCLK => net6683);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_04x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_4 port map( CLK => clk, EN 
                           => IF_RegsxN718, ENCLK => net6688);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_03x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_3 port map( CLK => clk, EN 
                           => IF_RegsxN719, ENCLK => net6693);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_02x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_2 port map( CLK => clk, EN 
                           => IF_RegsxN720, ENCLK => net6698);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_01x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_1 port map( CLK => clk, EN 
                           => IF_RegsxN721, ENCLK => net6703);
   U3773 : INV_X1 port map( A => n7624, ZN => toMemoryPortxREQxx1x(0));
   n7624 <= '1';

end SYN_CPU_arch;
