package testbasic12_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic12_SECTIONS;

endpackage
