library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package ModuleStateName02_types is
-- No local datatypes implemented!


end package ModuleStateName02_types;