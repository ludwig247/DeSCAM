library ieee;
use IEEE.numeric_std.all;

package TestBasic11_types is
type TestBasic11_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic11_types;
