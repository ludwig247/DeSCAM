package testfunction1_types;

	import scam_model_types::*;
endpackage