package testbasic4_types;

endpackage