library ieee;
use IEEE.numeric_std.all;
use work.SCAM_Model_types.all;

package TestBasic20_types is
type Sections is (SECTION_A, SECTION_B);
type color_t is (GREEN, RED, YELLOW);
end package TestBasic20_types;