package testbasic19_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic19_SECTIONS;

endpackage
