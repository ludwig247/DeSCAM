library ieee;
use IEEE.numeric_std.all;
use work.SCAM_Model_types.all;

package TestBasic4_types is
end package TestBasic4_types;