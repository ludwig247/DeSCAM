package testmasterslave13_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave13_SECTIONS;

endpackage
