
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_CPU is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
subtype bool is BOOLEAN range FALSE to TRUE ;
   
   -- Declarations for conversion functions.
   function std_logic_to_bool(arg : in std_logic) return bool;
   function bool_to_std_logic(arg : in bool) return std_logic;

end CONV_PACK_CPU;

package body CONV_PACK_CPU is
   
   -- std_logic to enum type function
   function std_logic_to_bool(arg : in std_logic) return bool is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when '0' => return FALSE;
         when '1' => return TRUE;
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return FALSE;
      end case;
   end;
   
   -- enum type to std_logic function
   function bool_to_std_logic(arg : in bool) return std_logic is
   -- synopsys built_in SYN_FEED_THRU;
   begin
      case arg is
         when FALSE => return '0';
         when TRUE => return '1';
         when others => assert FALSE -- this should not happen.
               report "un-convertible value"
               severity warning;
               return '0';
      end case;
   end;

end CONV_PACK_CPU;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_35 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_35;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_34 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_34;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_33 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_33;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_32 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_32;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_31 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_31;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_30 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_30;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_29 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_29;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_28 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_28;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_27 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_27;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_26 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_26;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_25 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_25;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_24 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_24;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_23 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_23;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_22 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_22;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_21 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_21;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_20 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_20;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_19 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_19;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_18 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_18;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_17 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_17;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_16 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_16;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_15 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_15;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_14 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_14;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_13 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_13;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_12 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_12;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_11 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_11;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_10 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_10;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_9 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_9;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_8 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_8;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_7 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_7;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_6 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_6;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_5 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_5;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_4 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_4;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_3 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_3;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_2 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_2;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_1 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_1;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_36 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_36;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity SNPS_CLOCK_GATE_HIGH_CPU_0 is

   port( CLK, EN : in std_logic;  ENCLK : out std_logic);

end SNPS_CLOCK_GATE_HIGH_CPU_0;

architecture SYN_USE_DEFA_ARCH_NAME of SNPS_CLOCK_GATE_HIGH_CPU_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal net325220 : std_logic;

begin
   
   latch : DLL_X1 port map( D => EN, GN => CLK, Q => net325220);
   main_gate : AND2_X1 port map( A1 => net325220, A2 => CLK, ZN => ENCLK);

end SYN_USE_DEFA_ARCH_NAME;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CPU.all;

entity CPU is

   port( clk, rst : in std_logic;  fromMemoryPortxLOADEDDATAx : in 
         std_logic_vector (31 downto 0);  fromMemoryPort_sync : in bool;  
         fromMemoryPort_notify : out bool;  toMemoryPort_sync : in bool;  
         toMemoryPort_notify : out bool;  toMemoryPortxADDRINxx31x, 
         toMemoryPortxADDRINxx30x, toMemoryPortxADDRINxx29x, 
         toMemoryPortxADDRINxx28x, toMemoryPortxADDRINxx27x, 
         toMemoryPortxADDRINxx26x, toMemoryPortxADDRINxx25x, 
         toMemoryPortxADDRINxx24x, toMemoryPortxADDRINxx23x, 
         toMemoryPortxADDRINxx22x, toMemoryPortxADDRINxx21x, 
         toMemoryPortxADDRINxx20x, toMemoryPortxADDRINxx19x, 
         toMemoryPortxADDRINxx18x, toMemoryPortxADDRINxx17x, 
         toMemoryPortxADDRINxx16x, toMemoryPortxADDRINxx15x, 
         toMemoryPortxADDRINxx14x, toMemoryPortxADDRINxx13x, 
         toMemoryPortxADDRINxx12x, toMemoryPortxADDRINxx11x, 
         toMemoryPortxADDRINxx10x, toMemoryPortxADDRINxx9x, 
         toMemoryPortxADDRINxx8x, toMemoryPortxADDRINxx7x, 
         toMemoryPortxADDRINxx6x, toMemoryPortxADDRINxx5x, 
         toMemoryPortxADDRINxx4x, toMemoryPortxADDRINxx3x, 
         toMemoryPortxADDRINxx2x, toMemoryPortxADDRINxx1x, 
         toMemoryPortxADDRINxx0x, toMemoryPortxDATAINxx31x, 
         toMemoryPortxDATAINxx30x, toMemoryPortxDATAINxx29x, 
         toMemoryPortxDATAINxx28x, toMemoryPortxDATAINxx27x, 
         toMemoryPortxDATAINxx26x, toMemoryPortxDATAINxx25x, 
         toMemoryPortxDATAINxx24x, toMemoryPortxDATAINxx23x, 
         toMemoryPortxDATAINxx22x, toMemoryPortxDATAINxx21x, 
         toMemoryPortxDATAINxx20x, toMemoryPortxDATAINxx19x, 
         toMemoryPortxDATAINxx18x, toMemoryPortxDATAINxx17x, 
         toMemoryPortxDATAINxx16x, toMemoryPortxDATAINxx15x, 
         toMemoryPortxDATAINxx14x, toMemoryPortxDATAINxx13x, 
         toMemoryPortxDATAINxx12x, toMemoryPortxDATAINxx11x, 
         toMemoryPortxDATAINxx10x, toMemoryPortxDATAINxx9x, 
         toMemoryPortxDATAINxx8x, toMemoryPortxDATAINxx7x, 
         toMemoryPortxDATAINxx6x, toMemoryPortxDATAINxx5x, 
         toMemoryPortxDATAINxx4x, toMemoryPortxDATAINxx3x, 
         toMemoryPortxDATAINxx2x, toMemoryPortxDATAINxx1x, 
         toMemoryPortxDATAINxx0x, toMemoryPortxMASKxx2x, toMemoryPortxMASKxx1x,
         toMemoryPortxMASKxx0x, toMemoryPortxREQxx1x, toMemoryPortxREQxx0x : 
         out std_logic_vector (0 to 0));

end CPU;

architecture SYN_CPU_arch of CPU is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_1
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_2
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_3
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_4
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_5
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_6
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_7
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_8
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_9
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_10
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_11
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_12
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_13
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_14
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_15
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_16
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_17
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_18
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_19
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_20
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_21
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_22
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_23
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_24
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_25
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_26
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_27
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_28
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_29
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_30
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_31
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_32
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_33
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_34
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_35
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_36
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component SNPS_CLOCK_GATE_HIGH_CPU_0
      port( CLK, EN : in std_logic;  ENCLK : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X4
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal fromMemoryPort_sync_port, toMemoryPort_sync_port, 
      toMemoryPort_notify_port, toRegsPortxDSTxx4x, toRegsPortxDSTxx3x, 
      toRegsPortxDSTxx2x, toRegsPortxDSTxx1x, toRegsPortxDSTxx0x, 
      toRegsPortxDSTDATAxx31x, toRegsPortxDSTDATAxx30x, toRegsPortxDSTDATAxx29x
      , toRegsPortxDSTDATAxx28x, toRegsPortxDSTDATAxx27x, 
      toRegsPortxDSTDATAxx26x, toRegsPortxDSTDATAxx25x, toRegsPortxDSTDATAxx24x
      , toRegsPortxDSTDATAxx23x, toRegsPortxDSTDATAxx22x, 
      toRegsPortxDSTDATAxx21x, toRegsPortxDSTDATAxx20x, toRegsPortxDSTDATAxx19x
      , toRegsPortxDSTDATAxx18x, toRegsPortxDSTDATAxx17x, 
      toRegsPortxDSTDATAxx16x, toRegsPortxDSTDATAxx15x, toRegsPortxDSTDATAxx14x
      , toRegsPortxDSTDATAxx13x, toRegsPortxDSTDATAxx12x, 
      toRegsPortxDSTDATAxx11x, toRegsPortxDSTDATAxx10x, toRegsPortxDSTDATAxx9x,
      toRegsPortxDSTDATAxx8x, toRegsPortxDSTDATAxx7x, toRegsPortxDSTDATAxx6x, 
      toRegsPortxDSTDATAxx5x, toRegsPortxDSTDATAxx4x, toRegsPortxDSTDATAxx3x, 
      toRegsPortxDSTDATAxx2x, toRegsPortxDSTDATAxx1x, toRegsPortxDSTDATAxx0x, 
      toRegsPort_notify, fromRegsPortxREG_FILE_01xx31x, 
      fromRegsPortxREG_FILE_01xx30x, fromRegsPortxREG_FILE_01xx29x, 
      fromRegsPortxREG_FILE_01xx28x, fromRegsPortxREG_FILE_01xx27x, 
      fromRegsPortxREG_FILE_01xx26x, fromRegsPortxREG_FILE_01xx25x, 
      fromRegsPortxREG_FILE_01xx24x, fromRegsPortxREG_FILE_01xx23x, 
      fromRegsPortxREG_FILE_01xx22x, fromRegsPortxREG_FILE_01xx21x, 
      fromRegsPortxREG_FILE_01xx20x, fromRegsPortxREG_FILE_01xx19x, 
      fromRegsPortxREG_FILE_01xx18x, fromRegsPortxREG_FILE_01xx17x, 
      fromRegsPortxREG_FILE_01xx16x, fromRegsPortxREG_FILE_01xx15x, 
      fromRegsPortxREG_FILE_01xx14x, fromRegsPortxREG_FILE_01xx13x, 
      fromRegsPortxREG_FILE_01xx12x, fromRegsPortxREG_FILE_01xx11x, 
      fromRegsPortxREG_FILE_01xx10x, fromRegsPortxREG_FILE_01xx9x, 
      fromRegsPortxREG_FILE_01xx8x, fromRegsPortxREG_FILE_01xx7x, 
      fromRegsPortxREG_FILE_01xx6x, fromRegsPortxREG_FILE_01xx5x, 
      fromRegsPortxREG_FILE_01xx4x, fromRegsPortxREG_FILE_01xx3x, 
      fromRegsPortxREG_FILE_01xx2x, fromRegsPortxREG_FILE_01xx1x, 
      fromRegsPortxREG_FILE_01xx0x, fromRegsPortxREG_FILE_02xx31x, 
      fromRegsPortxREG_FILE_02xx30x, fromRegsPortxREG_FILE_02xx29x, 
      fromRegsPortxREG_FILE_02xx28x, fromRegsPortxREG_FILE_02xx27x, 
      fromRegsPortxREG_FILE_02xx26x, fromRegsPortxREG_FILE_02xx25x, 
      fromRegsPortxREG_FILE_02xx24x, fromRegsPortxREG_FILE_02xx23x, 
      fromRegsPortxREG_FILE_02xx22x, fromRegsPortxREG_FILE_02xx21x, 
      fromRegsPortxREG_FILE_02xx20x, fromRegsPortxREG_FILE_02xx19x, 
      fromRegsPortxREG_FILE_02xx18x, fromRegsPortxREG_FILE_02xx17x, 
      fromRegsPortxREG_FILE_02xx16x, fromRegsPortxREG_FILE_02xx15x, 
      fromRegsPortxREG_FILE_02xx14x, fromRegsPortxREG_FILE_02xx13x, 
      fromRegsPortxREG_FILE_02xx12x, fromRegsPortxREG_FILE_02xx11x, 
      fromRegsPortxREG_FILE_02xx10x, fromRegsPortxREG_FILE_02xx9x, 
      fromRegsPortxREG_FILE_02xx8x, fromRegsPortxREG_FILE_02xx7x, 
      fromRegsPortxREG_FILE_02xx6x, fromRegsPortxREG_FILE_02xx5x, 
      fromRegsPortxREG_FILE_02xx4x, fromRegsPortxREG_FILE_02xx3x, 
      fromRegsPortxREG_FILE_02xx2x, fromRegsPortxREG_FILE_02xx1x, 
      fromRegsPortxREG_FILE_02xx0x, fromRegsPortxREG_FILE_03xx31x, 
      fromRegsPortxREG_FILE_03xx30x, fromRegsPortxREG_FILE_03xx29x, 
      fromRegsPortxREG_FILE_03xx28x, fromRegsPortxREG_FILE_03xx27x, 
      fromRegsPortxREG_FILE_03xx26x, fromRegsPortxREG_FILE_03xx25x, 
      fromRegsPortxREG_FILE_03xx24x, fromRegsPortxREG_FILE_03xx23x, 
      fromRegsPortxREG_FILE_03xx22x, fromRegsPortxREG_FILE_03xx21x, 
      fromRegsPortxREG_FILE_03xx20x, fromRegsPortxREG_FILE_03xx19x, 
      fromRegsPortxREG_FILE_03xx18x, fromRegsPortxREG_FILE_03xx17x, 
      fromRegsPortxREG_FILE_03xx16x, fromRegsPortxREG_FILE_03xx15x, 
      fromRegsPortxREG_FILE_03xx14x, fromRegsPortxREG_FILE_03xx13x, 
      fromRegsPortxREG_FILE_03xx12x, fromRegsPortxREG_FILE_03xx11x, 
      fromRegsPortxREG_FILE_03xx10x, fromRegsPortxREG_FILE_03xx9x, 
      fromRegsPortxREG_FILE_03xx8x, fromRegsPortxREG_FILE_03xx7x, 
      fromRegsPortxREG_FILE_03xx6x, fromRegsPortxREG_FILE_03xx5x, 
      fromRegsPortxREG_FILE_03xx4x, fromRegsPortxREG_FILE_03xx3x, 
      fromRegsPortxREG_FILE_03xx2x, fromRegsPortxREG_FILE_03xx1x, 
      fromRegsPortxREG_FILE_03xx0x, fromRegsPortxREG_FILE_04xx31x, 
      fromRegsPortxREG_FILE_04xx30x, fromRegsPortxREG_FILE_04xx29x, 
      fromRegsPortxREG_FILE_04xx28x, fromRegsPortxREG_FILE_04xx27x, 
      fromRegsPortxREG_FILE_04xx26x, fromRegsPortxREG_FILE_04xx25x, 
      fromRegsPortxREG_FILE_04xx24x, fromRegsPortxREG_FILE_04xx23x, 
      fromRegsPortxREG_FILE_04xx22x, fromRegsPortxREG_FILE_04xx21x, 
      fromRegsPortxREG_FILE_04xx20x, fromRegsPortxREG_FILE_04xx19x, 
      fromRegsPortxREG_FILE_04xx18x, fromRegsPortxREG_FILE_04xx17x, 
      fromRegsPortxREG_FILE_04xx16x, fromRegsPortxREG_FILE_04xx15x, 
      fromRegsPortxREG_FILE_04xx14x, fromRegsPortxREG_FILE_04xx13x, 
      fromRegsPortxREG_FILE_04xx12x, fromRegsPortxREG_FILE_04xx11x, 
      fromRegsPortxREG_FILE_04xx10x, fromRegsPortxREG_FILE_04xx9x, 
      fromRegsPortxREG_FILE_04xx8x, fromRegsPortxREG_FILE_04xx7x, 
      fromRegsPortxREG_FILE_04xx6x, fromRegsPortxREG_FILE_04xx5x, 
      fromRegsPortxREG_FILE_04xx4x, fromRegsPortxREG_FILE_04xx3x, 
      fromRegsPortxREG_FILE_04xx2x, fromRegsPortxREG_FILE_04xx1x, 
      fromRegsPortxREG_FILE_04xx0x, fromRegsPortxREG_FILE_05xx31x, 
      fromRegsPortxREG_FILE_05xx30x, fromRegsPortxREG_FILE_05xx29x, 
      fromRegsPortxREG_FILE_05xx28x, fromRegsPortxREG_FILE_05xx27x, 
      fromRegsPortxREG_FILE_05xx26x, fromRegsPortxREG_FILE_05xx25x, 
      fromRegsPortxREG_FILE_05xx24x, fromRegsPortxREG_FILE_05xx23x, 
      fromRegsPortxREG_FILE_05xx22x, fromRegsPortxREG_FILE_05xx21x, 
      fromRegsPortxREG_FILE_05xx20x, fromRegsPortxREG_FILE_05xx19x, 
      fromRegsPortxREG_FILE_05xx18x, fromRegsPortxREG_FILE_05xx17x, 
      fromRegsPortxREG_FILE_05xx16x, fromRegsPortxREG_FILE_05xx15x, 
      fromRegsPortxREG_FILE_05xx14x, fromRegsPortxREG_FILE_05xx13x, 
      fromRegsPortxREG_FILE_05xx12x, fromRegsPortxREG_FILE_05xx11x, 
      fromRegsPortxREG_FILE_05xx10x, fromRegsPortxREG_FILE_05xx9x, 
      fromRegsPortxREG_FILE_05xx8x, fromRegsPortxREG_FILE_05xx7x, 
      fromRegsPortxREG_FILE_05xx6x, fromRegsPortxREG_FILE_05xx5x, 
      fromRegsPortxREG_FILE_05xx4x, fromRegsPortxREG_FILE_05xx3x, 
      fromRegsPortxREG_FILE_05xx2x, fromRegsPortxREG_FILE_05xx1x, 
      fromRegsPortxREG_FILE_05xx0x, fromRegsPortxREG_FILE_06xx31x, 
      fromRegsPortxREG_FILE_06xx30x, fromRegsPortxREG_FILE_06xx29x, 
      fromRegsPortxREG_FILE_06xx28x, fromRegsPortxREG_FILE_06xx27x, 
      fromRegsPortxREG_FILE_06xx26x, fromRegsPortxREG_FILE_06xx25x, 
      fromRegsPortxREG_FILE_06xx24x, fromRegsPortxREG_FILE_06xx23x, 
      fromRegsPortxREG_FILE_06xx22x, fromRegsPortxREG_FILE_06xx21x, 
      fromRegsPortxREG_FILE_06xx20x, fromRegsPortxREG_FILE_06xx19x, 
      fromRegsPortxREG_FILE_06xx18x, fromRegsPortxREG_FILE_06xx17x, 
      fromRegsPortxREG_FILE_06xx16x, fromRegsPortxREG_FILE_06xx15x, 
      fromRegsPortxREG_FILE_06xx14x, fromRegsPortxREG_FILE_06xx13x, 
      fromRegsPortxREG_FILE_06xx12x, fromRegsPortxREG_FILE_06xx11x, 
      fromRegsPortxREG_FILE_06xx10x, fromRegsPortxREG_FILE_06xx9x, 
      fromRegsPortxREG_FILE_06xx8x, fromRegsPortxREG_FILE_06xx7x, 
      fromRegsPortxREG_FILE_06xx6x, fromRegsPortxREG_FILE_06xx5x, 
      fromRegsPortxREG_FILE_06xx4x, fromRegsPortxREG_FILE_06xx3x, 
      fromRegsPortxREG_FILE_06xx2x, fromRegsPortxREG_FILE_06xx1x, 
      fromRegsPortxREG_FILE_06xx0x, fromRegsPortxREG_FILE_07xx31x, 
      fromRegsPortxREG_FILE_07xx30x, fromRegsPortxREG_FILE_07xx29x, 
      fromRegsPortxREG_FILE_07xx28x, fromRegsPortxREG_FILE_07xx27x, 
      fromRegsPortxREG_FILE_07xx26x, fromRegsPortxREG_FILE_07xx25x, 
      fromRegsPortxREG_FILE_07xx24x, fromRegsPortxREG_FILE_07xx23x, 
      fromRegsPortxREG_FILE_07xx22x, fromRegsPortxREG_FILE_07xx21x, 
      fromRegsPortxREG_FILE_07xx20x, fromRegsPortxREG_FILE_07xx19x, 
      fromRegsPortxREG_FILE_07xx18x, fromRegsPortxREG_FILE_07xx17x, 
      fromRegsPortxREG_FILE_07xx16x, fromRegsPortxREG_FILE_07xx15x, 
      fromRegsPortxREG_FILE_07xx14x, fromRegsPortxREG_FILE_07xx13x, 
      fromRegsPortxREG_FILE_07xx12x, fromRegsPortxREG_FILE_07xx11x, 
      fromRegsPortxREG_FILE_07xx10x, fromRegsPortxREG_FILE_07xx9x, 
      fromRegsPortxREG_FILE_07xx8x, fromRegsPortxREG_FILE_07xx7x, 
      fromRegsPortxREG_FILE_07xx6x, fromRegsPortxREG_FILE_07xx5x, 
      fromRegsPortxREG_FILE_07xx4x, fromRegsPortxREG_FILE_07xx3x, 
      fromRegsPortxREG_FILE_07xx2x, fromRegsPortxREG_FILE_07xx1x, 
      fromRegsPortxREG_FILE_07xx0x, fromRegsPortxREG_FILE_08xx31x, 
      fromRegsPortxREG_FILE_08xx30x, fromRegsPortxREG_FILE_08xx29x, 
      fromRegsPortxREG_FILE_08xx28x, fromRegsPortxREG_FILE_08xx27x, 
      fromRegsPortxREG_FILE_08xx26x, fromRegsPortxREG_FILE_08xx25x, 
      fromRegsPortxREG_FILE_08xx24x, fromRegsPortxREG_FILE_08xx23x, 
      fromRegsPortxREG_FILE_08xx22x, fromRegsPortxREG_FILE_08xx21x, 
      fromRegsPortxREG_FILE_08xx20x, fromRegsPortxREG_FILE_08xx19x, 
      fromRegsPortxREG_FILE_08xx18x, fromRegsPortxREG_FILE_08xx17x, 
      fromRegsPortxREG_FILE_08xx16x, fromRegsPortxREG_FILE_08xx15x, 
      fromRegsPortxREG_FILE_08xx14x, fromRegsPortxREG_FILE_08xx13x, 
      fromRegsPortxREG_FILE_08xx12x, fromRegsPortxREG_FILE_08xx11x, 
      fromRegsPortxREG_FILE_08xx10x, fromRegsPortxREG_FILE_08xx9x, 
      fromRegsPortxREG_FILE_08xx8x, fromRegsPortxREG_FILE_08xx7x, 
      fromRegsPortxREG_FILE_08xx6x, fromRegsPortxREG_FILE_08xx5x, 
      fromRegsPortxREG_FILE_08xx4x, fromRegsPortxREG_FILE_08xx3x, 
      fromRegsPortxREG_FILE_08xx2x, fromRegsPortxREG_FILE_08xx1x, 
      fromRegsPortxREG_FILE_08xx0x, fromRegsPortxREG_FILE_09xx31x, 
      fromRegsPortxREG_FILE_09xx30x, fromRegsPortxREG_FILE_09xx29x, 
      fromRegsPortxREG_FILE_09xx28x, fromRegsPortxREG_FILE_09xx27x, 
      fromRegsPortxREG_FILE_09xx26x, fromRegsPortxREG_FILE_09xx25x, 
      fromRegsPortxREG_FILE_09xx24x, fromRegsPortxREG_FILE_09xx23x, 
      fromRegsPortxREG_FILE_09xx22x, fromRegsPortxREG_FILE_09xx21x, 
      fromRegsPortxREG_FILE_09xx20x, fromRegsPortxREG_FILE_09xx19x, 
      fromRegsPortxREG_FILE_09xx18x, fromRegsPortxREG_FILE_09xx17x, 
      fromRegsPortxREG_FILE_09xx16x, fromRegsPortxREG_FILE_09xx15x, 
      fromRegsPortxREG_FILE_09xx14x, fromRegsPortxREG_FILE_09xx13x, 
      fromRegsPortxREG_FILE_09xx12x, fromRegsPortxREG_FILE_09xx11x, 
      fromRegsPortxREG_FILE_09xx10x, fromRegsPortxREG_FILE_09xx9x, 
      fromRegsPortxREG_FILE_09xx8x, fromRegsPortxREG_FILE_09xx7x, 
      fromRegsPortxREG_FILE_09xx6x, fromRegsPortxREG_FILE_09xx5x, 
      fromRegsPortxREG_FILE_09xx4x, fromRegsPortxREG_FILE_09xx3x, 
      fromRegsPortxREG_FILE_09xx2x, fromRegsPortxREG_FILE_09xx1x, 
      fromRegsPortxREG_FILE_09xx0x, fromRegsPortxREG_FILE_10xx31x, 
      fromRegsPortxREG_FILE_10xx30x, fromRegsPortxREG_FILE_10xx29x, 
      fromRegsPortxREG_FILE_10xx28x, fromRegsPortxREG_FILE_10xx27x, 
      fromRegsPortxREG_FILE_10xx26x, fromRegsPortxREG_FILE_10xx25x, 
      fromRegsPortxREG_FILE_10xx24x, fromRegsPortxREG_FILE_10xx23x, 
      fromRegsPortxREG_FILE_10xx22x, fromRegsPortxREG_FILE_10xx21x, 
      fromRegsPortxREG_FILE_10xx20x, fromRegsPortxREG_FILE_10xx19x, 
      fromRegsPortxREG_FILE_10xx18x, fromRegsPortxREG_FILE_10xx17x, 
      fromRegsPortxREG_FILE_10xx16x, fromRegsPortxREG_FILE_10xx15x, 
      fromRegsPortxREG_FILE_10xx14x, fromRegsPortxREG_FILE_10xx13x, 
      fromRegsPortxREG_FILE_10xx12x, fromRegsPortxREG_FILE_10xx11x, 
      fromRegsPortxREG_FILE_10xx10x, fromRegsPortxREG_FILE_10xx9x, 
      fromRegsPortxREG_FILE_10xx8x, fromRegsPortxREG_FILE_10xx7x, 
      fromRegsPortxREG_FILE_10xx6x, fromRegsPortxREG_FILE_10xx5x, 
      fromRegsPortxREG_FILE_10xx4x, fromRegsPortxREG_FILE_10xx3x, 
      fromRegsPortxREG_FILE_10xx2x, fromRegsPortxREG_FILE_10xx1x, 
      fromRegsPortxREG_FILE_10xx0x, fromRegsPortxREG_FILE_11xx31x, 
      fromRegsPortxREG_FILE_11xx30x, fromRegsPortxREG_FILE_11xx29x, 
      fromRegsPortxREG_FILE_11xx28x, fromRegsPortxREG_FILE_11xx27x, 
      fromRegsPortxREG_FILE_11xx26x, fromRegsPortxREG_FILE_11xx25x, 
      fromRegsPortxREG_FILE_11xx24x, fromRegsPortxREG_FILE_11xx23x, 
      fromRegsPortxREG_FILE_11xx22x, fromRegsPortxREG_FILE_11xx21x, 
      fromRegsPortxREG_FILE_11xx20x, fromRegsPortxREG_FILE_11xx19x, 
      fromRegsPortxREG_FILE_11xx18x, fromRegsPortxREG_FILE_11xx17x, 
      fromRegsPortxREG_FILE_11xx16x, fromRegsPortxREG_FILE_11xx15x, 
      fromRegsPortxREG_FILE_11xx14x, fromRegsPortxREG_FILE_11xx13x, 
      fromRegsPortxREG_FILE_11xx12x, fromRegsPortxREG_FILE_11xx11x, 
      fromRegsPortxREG_FILE_11xx10x, fromRegsPortxREG_FILE_11xx9x, 
      fromRegsPortxREG_FILE_11xx8x, fromRegsPortxREG_FILE_11xx7x, 
      fromRegsPortxREG_FILE_11xx6x, fromRegsPortxREG_FILE_11xx5x, 
      fromRegsPortxREG_FILE_11xx4x, fromRegsPortxREG_FILE_11xx3x, 
      fromRegsPortxREG_FILE_11xx2x, fromRegsPortxREG_FILE_11xx1x, 
      fromRegsPortxREG_FILE_11xx0x, fromRegsPortxREG_FILE_12xx31x, 
      fromRegsPortxREG_FILE_12xx30x, fromRegsPortxREG_FILE_12xx29x, 
      fromRegsPortxREG_FILE_12xx28x, fromRegsPortxREG_FILE_12xx27x, 
      fromRegsPortxREG_FILE_12xx26x, fromRegsPortxREG_FILE_12xx25x, 
      fromRegsPortxREG_FILE_12xx24x, fromRegsPortxREG_FILE_12xx23x, 
      fromRegsPortxREG_FILE_12xx22x, fromRegsPortxREG_FILE_12xx21x, 
      fromRegsPortxREG_FILE_12xx20x, fromRegsPortxREG_FILE_12xx19x, 
      fromRegsPortxREG_FILE_12xx18x, fromRegsPortxREG_FILE_12xx17x, 
      fromRegsPortxREG_FILE_12xx16x, fromRegsPortxREG_FILE_12xx15x, 
      fromRegsPortxREG_FILE_12xx14x, fromRegsPortxREG_FILE_12xx13x, 
      fromRegsPortxREG_FILE_12xx12x, fromRegsPortxREG_FILE_12xx11x, 
      fromRegsPortxREG_FILE_12xx10x, fromRegsPortxREG_FILE_12xx9x, 
      fromRegsPortxREG_FILE_12xx8x, fromRegsPortxREG_FILE_12xx7x, 
      fromRegsPortxREG_FILE_12xx6x, fromRegsPortxREG_FILE_12xx5x, 
      fromRegsPortxREG_FILE_12xx4x, fromRegsPortxREG_FILE_12xx3x, 
      fromRegsPortxREG_FILE_12xx2x, fromRegsPortxREG_FILE_12xx1x, 
      fromRegsPortxREG_FILE_12xx0x, fromRegsPortxREG_FILE_13xx31x, 
      fromRegsPortxREG_FILE_13xx30x, fromRegsPortxREG_FILE_13xx29x, 
      fromRegsPortxREG_FILE_13xx28x, fromRegsPortxREG_FILE_13xx27x, 
      fromRegsPortxREG_FILE_13xx26x, fromRegsPortxREG_FILE_13xx25x, 
      fromRegsPortxREG_FILE_13xx24x, fromRegsPortxREG_FILE_13xx23x, 
      fromRegsPortxREG_FILE_13xx22x, fromRegsPortxREG_FILE_13xx21x, 
      fromRegsPortxREG_FILE_13xx20x, fromRegsPortxREG_FILE_13xx19x, 
      fromRegsPortxREG_FILE_13xx18x, fromRegsPortxREG_FILE_13xx17x, 
      fromRegsPortxREG_FILE_13xx16x, fromRegsPortxREG_FILE_13xx15x, 
      fromRegsPortxREG_FILE_13xx14x, fromRegsPortxREG_FILE_13xx13x, 
      fromRegsPortxREG_FILE_13xx12x, fromRegsPortxREG_FILE_13xx11x, 
      fromRegsPortxREG_FILE_13xx10x, fromRegsPortxREG_FILE_13xx9x, 
      fromRegsPortxREG_FILE_13xx8x, fromRegsPortxREG_FILE_13xx7x, 
      fromRegsPortxREG_FILE_13xx6x, fromRegsPortxREG_FILE_13xx5x, 
      fromRegsPortxREG_FILE_13xx4x, fromRegsPortxREG_FILE_13xx3x, 
      fromRegsPortxREG_FILE_13xx2x, fromRegsPortxREG_FILE_13xx1x, 
      fromRegsPortxREG_FILE_13xx0x, fromRegsPortxREG_FILE_14xx31x, 
      fromRegsPortxREG_FILE_14xx30x, fromRegsPortxREG_FILE_14xx29x, 
      fromRegsPortxREG_FILE_14xx28x, fromRegsPortxREG_FILE_14xx27x, 
      fromRegsPortxREG_FILE_14xx26x, fromRegsPortxREG_FILE_14xx25x, 
      fromRegsPortxREG_FILE_14xx24x, fromRegsPortxREG_FILE_14xx23x, 
      fromRegsPortxREG_FILE_14xx22x, fromRegsPortxREG_FILE_14xx21x, 
      fromRegsPortxREG_FILE_14xx20x, fromRegsPortxREG_FILE_14xx19x, 
      fromRegsPortxREG_FILE_14xx18x, fromRegsPortxREG_FILE_14xx17x, 
      fromRegsPortxREG_FILE_14xx16x, fromRegsPortxREG_FILE_14xx15x, 
      fromRegsPortxREG_FILE_14xx14x, fromRegsPortxREG_FILE_14xx13x, 
      fromRegsPortxREG_FILE_14xx12x, fromRegsPortxREG_FILE_14xx11x, 
      fromRegsPortxREG_FILE_14xx10x, fromRegsPortxREG_FILE_14xx9x, 
      fromRegsPortxREG_FILE_14xx8x, fromRegsPortxREG_FILE_14xx7x, 
      fromRegsPortxREG_FILE_14xx6x, fromRegsPortxREG_FILE_14xx5x, 
      fromRegsPortxREG_FILE_14xx4x, fromRegsPortxREG_FILE_14xx3x, 
      fromRegsPortxREG_FILE_14xx2x, fromRegsPortxREG_FILE_14xx1x, 
      fromRegsPortxREG_FILE_14xx0x, fromRegsPortxREG_FILE_15xx31x, 
      fromRegsPortxREG_FILE_15xx30x, fromRegsPortxREG_FILE_15xx29x, 
      fromRegsPortxREG_FILE_15xx28x, fromRegsPortxREG_FILE_15xx27x, 
      fromRegsPortxREG_FILE_15xx26x, fromRegsPortxREG_FILE_15xx25x, 
      fromRegsPortxREG_FILE_15xx24x, fromRegsPortxREG_FILE_15xx23x, 
      fromRegsPortxREG_FILE_15xx22x, fromRegsPortxREG_FILE_15xx21x, 
      fromRegsPortxREG_FILE_15xx20x, fromRegsPortxREG_FILE_15xx19x, 
      fromRegsPortxREG_FILE_15xx18x, fromRegsPortxREG_FILE_15xx17x, 
      fromRegsPortxREG_FILE_15xx16x, fromRegsPortxREG_FILE_15xx15x, 
      fromRegsPortxREG_FILE_15xx14x, fromRegsPortxREG_FILE_15xx13x, 
      fromRegsPortxREG_FILE_15xx12x, fromRegsPortxREG_FILE_15xx11x, 
      fromRegsPortxREG_FILE_15xx10x, fromRegsPortxREG_FILE_15xx9x, 
      fromRegsPortxREG_FILE_15xx8x, fromRegsPortxREG_FILE_15xx7x, 
      fromRegsPortxREG_FILE_15xx6x, fromRegsPortxREG_FILE_15xx5x, 
      fromRegsPortxREG_FILE_15xx4x, fromRegsPortxREG_FILE_15xx3x, 
      fromRegsPortxREG_FILE_15xx2x, fromRegsPortxREG_FILE_15xx1x, 
      fromRegsPortxREG_FILE_15xx0x, fromRegsPortxREG_FILE_16xx31x, 
      fromRegsPortxREG_FILE_16xx30x, fromRegsPortxREG_FILE_16xx29x, 
      fromRegsPortxREG_FILE_16xx28x, fromRegsPortxREG_FILE_16xx27x, 
      fromRegsPortxREG_FILE_16xx26x, fromRegsPortxREG_FILE_16xx25x, 
      fromRegsPortxREG_FILE_16xx24x, fromRegsPortxREG_FILE_16xx23x, 
      fromRegsPortxREG_FILE_16xx22x, fromRegsPortxREG_FILE_16xx21x, 
      fromRegsPortxREG_FILE_16xx20x, fromRegsPortxREG_FILE_16xx19x, 
      fromRegsPortxREG_FILE_16xx18x, fromRegsPortxREG_FILE_16xx17x, 
      fromRegsPortxREG_FILE_16xx16x, fromRegsPortxREG_FILE_16xx15x, 
      fromRegsPortxREG_FILE_16xx14x, fromRegsPortxREG_FILE_16xx13x, 
      fromRegsPortxREG_FILE_16xx12x, fromRegsPortxREG_FILE_16xx11x, 
      fromRegsPortxREG_FILE_16xx10x, fromRegsPortxREG_FILE_16xx9x, 
      fromRegsPortxREG_FILE_16xx8x, fromRegsPortxREG_FILE_16xx7x, 
      fromRegsPortxREG_FILE_16xx6x, fromRegsPortxREG_FILE_16xx5x, 
      fromRegsPortxREG_FILE_16xx4x, fromRegsPortxREG_FILE_16xx3x, 
      fromRegsPortxREG_FILE_16xx2x, fromRegsPortxREG_FILE_16xx1x, 
      fromRegsPortxREG_FILE_16xx0x, fromRegsPortxREG_FILE_17xx31x, 
      fromRegsPortxREG_FILE_17xx30x, fromRegsPortxREG_FILE_17xx29x, 
      fromRegsPortxREG_FILE_17xx28x, fromRegsPortxREG_FILE_17xx27x, 
      fromRegsPortxREG_FILE_17xx26x, fromRegsPortxREG_FILE_17xx25x, 
      fromRegsPortxREG_FILE_17xx24x, fromRegsPortxREG_FILE_17xx23x, 
      fromRegsPortxREG_FILE_17xx22x, fromRegsPortxREG_FILE_17xx21x, 
      fromRegsPortxREG_FILE_17xx20x, fromRegsPortxREG_FILE_17xx19x, 
      fromRegsPortxREG_FILE_17xx18x, fromRegsPortxREG_FILE_17xx17x, 
      fromRegsPortxREG_FILE_17xx16x, fromRegsPortxREG_FILE_17xx15x, 
      fromRegsPortxREG_FILE_17xx14x, fromRegsPortxREG_FILE_17xx13x, 
      fromRegsPortxREG_FILE_17xx12x, fromRegsPortxREG_FILE_17xx11x, 
      fromRegsPortxREG_FILE_17xx10x, fromRegsPortxREG_FILE_17xx9x, 
      fromRegsPortxREG_FILE_17xx8x, fromRegsPortxREG_FILE_17xx7x, 
      fromRegsPortxREG_FILE_17xx6x, fromRegsPortxREG_FILE_17xx5x, 
      fromRegsPortxREG_FILE_17xx4x, fromRegsPortxREG_FILE_17xx3x, 
      fromRegsPortxREG_FILE_17xx2x, fromRegsPortxREG_FILE_17xx1x, 
      fromRegsPortxREG_FILE_17xx0x, fromRegsPortxREG_FILE_18xx31x, 
      fromRegsPortxREG_FILE_18xx30x, fromRegsPortxREG_FILE_18xx29x, 
      fromRegsPortxREG_FILE_18xx28x, fromRegsPortxREG_FILE_18xx27x, 
      fromRegsPortxREG_FILE_18xx26x, fromRegsPortxREG_FILE_18xx25x, 
      fromRegsPortxREG_FILE_18xx24x, fromRegsPortxREG_FILE_18xx23x, 
      fromRegsPortxREG_FILE_18xx22x, fromRegsPortxREG_FILE_18xx21x, 
      fromRegsPortxREG_FILE_18xx20x, fromRegsPortxREG_FILE_18xx19x, 
      fromRegsPortxREG_FILE_18xx18x, fromRegsPortxREG_FILE_18xx17x, 
      fromRegsPortxREG_FILE_18xx16x, fromRegsPortxREG_FILE_18xx15x, 
      fromRegsPortxREG_FILE_18xx14x, fromRegsPortxREG_FILE_18xx13x, 
      fromRegsPortxREG_FILE_18xx12x, fromRegsPortxREG_FILE_18xx11x, 
      fromRegsPortxREG_FILE_18xx10x, fromRegsPortxREG_FILE_18xx9x, 
      fromRegsPortxREG_FILE_18xx8x, fromRegsPortxREG_FILE_18xx7x, 
      fromRegsPortxREG_FILE_18xx6x, fromRegsPortxREG_FILE_18xx5x, 
      fromRegsPortxREG_FILE_18xx4x, fromRegsPortxREG_FILE_18xx3x, 
      fromRegsPortxREG_FILE_18xx2x, fromRegsPortxREG_FILE_18xx1x, 
      fromRegsPortxREG_FILE_18xx0x, fromRegsPortxREG_FILE_19xx31x, 
      fromRegsPortxREG_FILE_19xx30x, fromRegsPortxREG_FILE_19xx29x, 
      fromRegsPortxREG_FILE_19xx28x, fromRegsPortxREG_FILE_19xx27x, 
      fromRegsPortxREG_FILE_19xx26x, fromRegsPortxREG_FILE_19xx25x, 
      fromRegsPortxREG_FILE_19xx24x, fromRegsPortxREG_FILE_19xx23x, 
      fromRegsPortxREG_FILE_19xx22x, fromRegsPortxREG_FILE_19xx21x, 
      fromRegsPortxREG_FILE_19xx20x, fromRegsPortxREG_FILE_19xx19x, 
      fromRegsPortxREG_FILE_19xx18x, fromRegsPortxREG_FILE_19xx17x, 
      fromRegsPortxREG_FILE_19xx16x, fromRegsPortxREG_FILE_19xx15x, 
      fromRegsPortxREG_FILE_19xx14x, fromRegsPortxREG_FILE_19xx13x, 
      fromRegsPortxREG_FILE_19xx12x, fromRegsPortxREG_FILE_19xx11x, 
      fromRegsPortxREG_FILE_19xx10x, fromRegsPortxREG_FILE_19xx9x, 
      fromRegsPortxREG_FILE_19xx8x, fromRegsPortxREG_FILE_19xx7x, 
      fromRegsPortxREG_FILE_19xx6x, fromRegsPortxREG_FILE_19xx5x, 
      fromRegsPortxREG_FILE_19xx4x, fromRegsPortxREG_FILE_19xx3x, 
      fromRegsPortxREG_FILE_19xx2x, fromRegsPortxREG_FILE_19xx1x, 
      fromRegsPortxREG_FILE_19xx0x, fromRegsPortxREG_FILE_20xx31x, 
      fromRegsPortxREG_FILE_20xx30x, fromRegsPortxREG_FILE_20xx29x, 
      fromRegsPortxREG_FILE_20xx28x, fromRegsPortxREG_FILE_20xx27x, 
      fromRegsPortxREG_FILE_20xx26x, fromRegsPortxREG_FILE_20xx25x, 
      fromRegsPortxREG_FILE_20xx24x, fromRegsPortxREG_FILE_20xx23x, 
      fromRegsPortxREG_FILE_20xx22x, fromRegsPortxREG_FILE_20xx21x, 
      fromRegsPortxREG_FILE_20xx20x, fromRegsPortxREG_FILE_20xx19x, 
      fromRegsPortxREG_FILE_20xx18x, fromRegsPortxREG_FILE_20xx17x, 
      fromRegsPortxREG_FILE_20xx16x, fromRegsPortxREG_FILE_20xx15x, 
      fromRegsPortxREG_FILE_20xx14x, fromRegsPortxREG_FILE_20xx13x, 
      fromRegsPortxREG_FILE_20xx12x, fromRegsPortxREG_FILE_20xx11x, 
      fromRegsPortxREG_FILE_20xx10x, fromRegsPortxREG_FILE_20xx9x, 
      fromRegsPortxREG_FILE_20xx8x, fromRegsPortxREG_FILE_20xx7x, 
      fromRegsPortxREG_FILE_20xx6x, fromRegsPortxREG_FILE_20xx5x, 
      fromRegsPortxREG_FILE_20xx4x, fromRegsPortxREG_FILE_20xx3x, 
      fromRegsPortxREG_FILE_20xx2x, fromRegsPortxREG_FILE_20xx1x, 
      fromRegsPortxREG_FILE_20xx0x, fromRegsPortxREG_FILE_21xx31x, 
      fromRegsPortxREG_FILE_21xx30x, fromRegsPortxREG_FILE_21xx29x, 
      fromRegsPortxREG_FILE_21xx28x, fromRegsPortxREG_FILE_21xx27x, 
      fromRegsPortxREG_FILE_21xx26x, fromRegsPortxREG_FILE_21xx25x, 
      fromRegsPortxREG_FILE_21xx24x, fromRegsPortxREG_FILE_21xx23x, 
      fromRegsPortxREG_FILE_21xx22x, fromRegsPortxREG_FILE_21xx21x, 
      fromRegsPortxREG_FILE_21xx20x, fromRegsPortxREG_FILE_21xx19x, 
      fromRegsPortxREG_FILE_21xx18x, fromRegsPortxREG_FILE_21xx17x, 
      fromRegsPortxREG_FILE_21xx16x, fromRegsPortxREG_FILE_21xx15x, 
      fromRegsPortxREG_FILE_21xx14x, fromRegsPortxREG_FILE_21xx13x, 
      fromRegsPortxREG_FILE_21xx12x, fromRegsPortxREG_FILE_21xx11x, 
      fromRegsPortxREG_FILE_21xx10x, fromRegsPortxREG_FILE_21xx9x, 
      fromRegsPortxREG_FILE_21xx8x, fromRegsPortxREG_FILE_21xx7x, 
      fromRegsPortxREG_FILE_21xx6x, fromRegsPortxREG_FILE_21xx5x, 
      fromRegsPortxREG_FILE_21xx4x, fromRegsPortxREG_FILE_21xx3x, 
      fromRegsPortxREG_FILE_21xx2x, fromRegsPortxREG_FILE_21xx1x, 
      fromRegsPortxREG_FILE_21xx0x, fromRegsPortxREG_FILE_22xx31x, 
      fromRegsPortxREG_FILE_22xx30x, fromRegsPortxREG_FILE_22xx29x, 
      fromRegsPortxREG_FILE_22xx28x, fromRegsPortxREG_FILE_22xx27x, 
      fromRegsPortxREG_FILE_22xx26x, fromRegsPortxREG_FILE_22xx25x, 
      fromRegsPortxREG_FILE_22xx24x, fromRegsPortxREG_FILE_22xx23x, 
      fromRegsPortxREG_FILE_22xx22x, fromRegsPortxREG_FILE_22xx21x, 
      fromRegsPortxREG_FILE_22xx20x, fromRegsPortxREG_FILE_22xx19x, 
      fromRegsPortxREG_FILE_22xx18x, fromRegsPortxREG_FILE_22xx17x, 
      fromRegsPortxREG_FILE_22xx16x, fromRegsPortxREG_FILE_22xx15x, 
      fromRegsPortxREG_FILE_22xx14x, fromRegsPortxREG_FILE_22xx13x, 
      fromRegsPortxREG_FILE_22xx12x, fromRegsPortxREG_FILE_22xx11x, 
      fromRegsPortxREG_FILE_22xx10x, fromRegsPortxREG_FILE_22xx9x, 
      fromRegsPortxREG_FILE_22xx8x, fromRegsPortxREG_FILE_22xx7x, 
      fromRegsPortxREG_FILE_22xx6x, fromRegsPortxREG_FILE_22xx5x, 
      fromRegsPortxREG_FILE_22xx4x, fromRegsPortxREG_FILE_22xx3x, 
      fromRegsPortxREG_FILE_22xx2x, fromRegsPortxREG_FILE_22xx1x, 
      fromRegsPortxREG_FILE_22xx0x, fromRegsPortxREG_FILE_23xx31x, 
      fromRegsPortxREG_FILE_23xx30x, fromRegsPortxREG_FILE_23xx29x, 
      fromRegsPortxREG_FILE_23xx28x, fromRegsPortxREG_FILE_23xx27x, 
      fromRegsPortxREG_FILE_23xx26x, fromRegsPortxREG_FILE_23xx25x, 
      fromRegsPortxREG_FILE_23xx24x, fromRegsPortxREG_FILE_23xx23x, 
      fromRegsPortxREG_FILE_23xx22x, fromRegsPortxREG_FILE_23xx21x, 
      fromRegsPortxREG_FILE_23xx20x, fromRegsPortxREG_FILE_23xx19x, 
      fromRegsPortxREG_FILE_23xx18x, fromRegsPortxREG_FILE_23xx17x, 
      fromRegsPortxREG_FILE_23xx16x, fromRegsPortxREG_FILE_23xx15x, 
      fromRegsPortxREG_FILE_23xx14x, fromRegsPortxREG_FILE_23xx13x, 
      fromRegsPortxREG_FILE_23xx12x, fromRegsPortxREG_FILE_23xx11x, 
      fromRegsPortxREG_FILE_23xx10x, fromRegsPortxREG_FILE_23xx9x, 
      fromRegsPortxREG_FILE_23xx8x, fromRegsPortxREG_FILE_23xx7x, 
      fromRegsPortxREG_FILE_23xx6x, fromRegsPortxREG_FILE_23xx5x, 
      fromRegsPortxREG_FILE_23xx4x, fromRegsPortxREG_FILE_23xx3x, 
      fromRegsPortxREG_FILE_23xx2x, fromRegsPortxREG_FILE_23xx1x, 
      fromRegsPortxREG_FILE_23xx0x, fromRegsPortxREG_FILE_24xx31x, 
      fromRegsPortxREG_FILE_24xx30x, fromRegsPortxREG_FILE_24xx29x, 
      fromRegsPortxREG_FILE_24xx28x, fromRegsPortxREG_FILE_24xx27x, 
      fromRegsPortxREG_FILE_24xx26x, fromRegsPortxREG_FILE_24xx25x, 
      fromRegsPortxREG_FILE_24xx24x, fromRegsPortxREG_FILE_24xx23x, 
      fromRegsPortxREG_FILE_24xx22x, fromRegsPortxREG_FILE_24xx21x, 
      fromRegsPortxREG_FILE_24xx20x, fromRegsPortxREG_FILE_24xx19x, 
      fromRegsPortxREG_FILE_24xx18x, fromRegsPortxREG_FILE_24xx17x, 
      fromRegsPortxREG_FILE_24xx16x, fromRegsPortxREG_FILE_24xx15x, 
      fromRegsPortxREG_FILE_24xx14x, fromRegsPortxREG_FILE_24xx13x, 
      fromRegsPortxREG_FILE_24xx12x, fromRegsPortxREG_FILE_24xx11x, 
      fromRegsPortxREG_FILE_24xx10x, fromRegsPortxREG_FILE_24xx9x, 
      fromRegsPortxREG_FILE_24xx8x, fromRegsPortxREG_FILE_24xx7x, 
      fromRegsPortxREG_FILE_24xx6x, fromRegsPortxREG_FILE_24xx5x, 
      fromRegsPortxREG_FILE_24xx4x, fromRegsPortxREG_FILE_24xx3x, 
      fromRegsPortxREG_FILE_24xx2x, fromRegsPortxREG_FILE_24xx1x, 
      fromRegsPortxREG_FILE_24xx0x, fromRegsPortxREG_FILE_25xx31x, 
      fromRegsPortxREG_FILE_25xx30x, fromRegsPortxREG_FILE_25xx29x, 
      fromRegsPortxREG_FILE_25xx28x, fromRegsPortxREG_FILE_25xx27x, 
      fromRegsPortxREG_FILE_25xx26x, fromRegsPortxREG_FILE_25xx25x, 
      fromRegsPortxREG_FILE_25xx24x, fromRegsPortxREG_FILE_25xx23x, 
      fromRegsPortxREG_FILE_25xx22x, fromRegsPortxREG_FILE_25xx21x, 
      fromRegsPortxREG_FILE_25xx20x, fromRegsPortxREG_FILE_25xx19x, 
      fromRegsPortxREG_FILE_25xx18x, fromRegsPortxREG_FILE_25xx17x, 
      fromRegsPortxREG_FILE_25xx16x, fromRegsPortxREG_FILE_25xx15x, 
      fromRegsPortxREG_FILE_25xx14x, fromRegsPortxREG_FILE_25xx13x, 
      fromRegsPortxREG_FILE_25xx12x, fromRegsPortxREG_FILE_25xx11x, 
      fromRegsPortxREG_FILE_25xx10x, fromRegsPortxREG_FILE_25xx9x, 
      fromRegsPortxREG_FILE_25xx8x, fromRegsPortxREG_FILE_25xx7x, 
      fromRegsPortxREG_FILE_25xx6x, fromRegsPortxREG_FILE_25xx5x, 
      fromRegsPortxREG_FILE_25xx4x, fromRegsPortxREG_FILE_25xx3x, 
      fromRegsPortxREG_FILE_25xx2x, fromRegsPortxREG_FILE_25xx1x, 
      fromRegsPortxREG_FILE_25xx0x, fromRegsPortxREG_FILE_26xx31x, 
      fromRegsPortxREG_FILE_26xx30x, fromRegsPortxREG_FILE_26xx29x, 
      fromRegsPortxREG_FILE_26xx28x, fromRegsPortxREG_FILE_26xx27x, 
      fromRegsPortxREG_FILE_26xx26x, fromRegsPortxREG_FILE_26xx25x, 
      fromRegsPortxREG_FILE_26xx24x, fromRegsPortxREG_FILE_26xx23x, 
      fromRegsPortxREG_FILE_26xx22x, fromRegsPortxREG_FILE_26xx21x, 
      fromRegsPortxREG_FILE_26xx20x, fromRegsPortxREG_FILE_26xx19x, 
      fromRegsPortxREG_FILE_26xx18x, fromRegsPortxREG_FILE_26xx17x, 
      fromRegsPortxREG_FILE_26xx16x, fromRegsPortxREG_FILE_26xx15x, 
      fromRegsPortxREG_FILE_26xx14x, fromRegsPortxREG_FILE_26xx13x, 
      fromRegsPortxREG_FILE_26xx12x, fromRegsPortxREG_FILE_26xx11x, 
      fromRegsPortxREG_FILE_26xx10x, fromRegsPortxREG_FILE_26xx9x, 
      fromRegsPortxREG_FILE_26xx8x, fromRegsPortxREG_FILE_26xx7x, 
      fromRegsPortxREG_FILE_26xx6x, fromRegsPortxREG_FILE_26xx5x, 
      fromRegsPortxREG_FILE_26xx4x, fromRegsPortxREG_FILE_26xx3x, 
      fromRegsPortxREG_FILE_26xx2x, fromRegsPortxREG_FILE_26xx1x, 
      fromRegsPortxREG_FILE_26xx0x, fromRegsPortxREG_FILE_27xx31x, 
      fromRegsPortxREG_FILE_27xx30x, fromRegsPortxREG_FILE_27xx29x, 
      fromRegsPortxREG_FILE_27xx28x, fromRegsPortxREG_FILE_27xx27x, 
      fromRegsPortxREG_FILE_27xx26x, fromRegsPortxREG_FILE_27xx25x, 
      fromRegsPortxREG_FILE_27xx24x, fromRegsPortxREG_FILE_27xx23x, 
      fromRegsPortxREG_FILE_27xx22x, fromRegsPortxREG_FILE_27xx21x, 
      fromRegsPortxREG_FILE_27xx20x, fromRegsPortxREG_FILE_27xx19x, 
      fromRegsPortxREG_FILE_27xx18x, fromRegsPortxREG_FILE_27xx17x, 
      fromRegsPortxREG_FILE_27xx16x, fromRegsPortxREG_FILE_27xx15x, 
      fromRegsPortxREG_FILE_27xx14x, fromRegsPortxREG_FILE_27xx13x, 
      fromRegsPortxREG_FILE_27xx12x, fromRegsPortxREG_FILE_27xx11x, 
      fromRegsPortxREG_FILE_27xx10x, fromRegsPortxREG_FILE_27xx9x, 
      fromRegsPortxREG_FILE_27xx8x, fromRegsPortxREG_FILE_27xx7x, 
      fromRegsPortxREG_FILE_27xx6x, fromRegsPortxREG_FILE_27xx5x, 
      fromRegsPortxREG_FILE_27xx4x, fromRegsPortxREG_FILE_27xx3x, 
      fromRegsPortxREG_FILE_27xx2x, fromRegsPortxREG_FILE_27xx1x, 
      fromRegsPortxREG_FILE_27xx0x, fromRegsPortxREG_FILE_28xx31x, 
      fromRegsPortxREG_FILE_28xx30x, fromRegsPortxREG_FILE_28xx29x, 
      fromRegsPortxREG_FILE_28xx28x, fromRegsPortxREG_FILE_28xx27x, 
      fromRegsPortxREG_FILE_28xx26x, fromRegsPortxREG_FILE_28xx25x, 
      fromRegsPortxREG_FILE_28xx24x, fromRegsPortxREG_FILE_28xx23x, 
      fromRegsPortxREG_FILE_28xx22x, fromRegsPortxREG_FILE_28xx21x, 
      fromRegsPortxREG_FILE_28xx20x, fromRegsPortxREG_FILE_28xx19x, 
      fromRegsPortxREG_FILE_28xx18x, fromRegsPortxREG_FILE_28xx17x, 
      fromRegsPortxREG_FILE_28xx16x, fromRegsPortxREG_FILE_28xx15x, 
      fromRegsPortxREG_FILE_28xx14x, fromRegsPortxREG_FILE_28xx13x, 
      fromRegsPortxREG_FILE_28xx12x, fromRegsPortxREG_FILE_28xx11x, 
      fromRegsPortxREG_FILE_28xx10x, fromRegsPortxREG_FILE_28xx9x, 
      fromRegsPortxREG_FILE_28xx8x, fromRegsPortxREG_FILE_28xx7x, 
      fromRegsPortxREG_FILE_28xx6x, fromRegsPortxREG_FILE_28xx5x, 
      fromRegsPortxREG_FILE_28xx4x, fromRegsPortxREG_FILE_28xx3x, 
      fromRegsPortxREG_FILE_28xx2x, fromRegsPortxREG_FILE_28xx1x, 
      fromRegsPortxREG_FILE_28xx0x, fromRegsPortxREG_FILE_29xx31x, 
      fromRegsPortxREG_FILE_29xx30x, fromRegsPortxREG_FILE_29xx29x, 
      fromRegsPortxREG_FILE_29xx28x, fromRegsPortxREG_FILE_29xx27x, 
      fromRegsPortxREG_FILE_29xx26x, fromRegsPortxREG_FILE_29xx25x, 
      fromRegsPortxREG_FILE_29xx24x, fromRegsPortxREG_FILE_29xx23x, 
      fromRegsPortxREG_FILE_29xx22x, fromRegsPortxREG_FILE_29xx21x, 
      fromRegsPortxREG_FILE_29xx20x, fromRegsPortxREG_FILE_29xx19x, 
      fromRegsPortxREG_FILE_29xx18x, fromRegsPortxREG_FILE_29xx17x, 
      fromRegsPortxREG_FILE_29xx16x, fromRegsPortxREG_FILE_29xx15x, 
      fromRegsPortxREG_FILE_29xx14x, fromRegsPortxREG_FILE_29xx13x, 
      fromRegsPortxREG_FILE_29xx12x, fromRegsPortxREG_FILE_29xx11x, 
      fromRegsPortxREG_FILE_29xx10x, fromRegsPortxREG_FILE_29xx9x, 
      fromRegsPortxREG_FILE_29xx8x, fromRegsPortxREG_FILE_29xx7x, 
      fromRegsPortxREG_FILE_29xx6x, fromRegsPortxREG_FILE_29xx5x, 
      fromRegsPortxREG_FILE_29xx4x, fromRegsPortxREG_FILE_29xx3x, 
      fromRegsPortxREG_FILE_29xx2x, fromRegsPortxREG_FILE_29xx1x, 
      fromRegsPortxREG_FILE_29xx0x, fromRegsPortxREG_FILE_30xx31x, 
      fromRegsPortxREG_FILE_30xx30x, fromRegsPortxREG_FILE_30xx29x, 
      fromRegsPortxREG_FILE_30xx28x, fromRegsPortxREG_FILE_30xx27x, 
      fromRegsPortxREG_FILE_30xx26x, fromRegsPortxREG_FILE_30xx25x, 
      fromRegsPortxREG_FILE_30xx24x, fromRegsPortxREG_FILE_30xx23x, 
      fromRegsPortxREG_FILE_30xx22x, fromRegsPortxREG_FILE_30xx21x, 
      fromRegsPortxREG_FILE_30xx20x, fromRegsPortxREG_FILE_30xx19x, 
      fromRegsPortxREG_FILE_30xx18x, fromRegsPortxREG_FILE_30xx17x, 
      fromRegsPortxREG_FILE_30xx16x, fromRegsPortxREG_FILE_30xx15x, 
      fromRegsPortxREG_FILE_30xx14x, fromRegsPortxREG_FILE_30xx13x, 
      fromRegsPortxREG_FILE_30xx12x, fromRegsPortxREG_FILE_30xx11x, 
      fromRegsPortxREG_FILE_30xx10x, fromRegsPortxREG_FILE_30xx9x, 
      fromRegsPortxREG_FILE_30xx8x, fromRegsPortxREG_FILE_30xx7x, 
      fromRegsPortxREG_FILE_30xx6x, fromRegsPortxREG_FILE_30xx5x, 
      fromRegsPortxREG_FILE_30xx4x, fromRegsPortxREG_FILE_30xx3x, 
      fromRegsPortxREG_FILE_30xx2x, fromRegsPortxREG_FILE_30xx1x, 
      fromRegsPortxREG_FILE_30xx0x, fromRegsPortxREG_FILE_31xx31x, 
      fromRegsPortxREG_FILE_31xx30x, fromRegsPortxREG_FILE_31xx29x, 
      fromRegsPortxREG_FILE_31xx28x, fromRegsPortxREG_FILE_31xx27x, 
      fromRegsPortxREG_FILE_31xx26x, fromRegsPortxREG_FILE_31xx25x, 
      fromRegsPortxREG_FILE_31xx24x, fromRegsPortxREG_FILE_31xx23x, 
      fromRegsPortxREG_FILE_31xx22x, fromRegsPortxREG_FILE_31xx21x, 
      fromRegsPortxREG_FILE_31xx20x, fromRegsPortxREG_FILE_31xx19x, 
      fromRegsPortxREG_FILE_31xx18x, fromRegsPortxREG_FILE_31xx17x, 
      fromRegsPortxREG_FILE_31xx16x, fromRegsPortxREG_FILE_31xx15x, 
      fromRegsPortxREG_FILE_31xx14x, fromRegsPortxREG_FILE_31xx13x, 
      fromRegsPortxREG_FILE_31xx12x, fromRegsPortxREG_FILE_31xx11x, 
      fromRegsPortxREG_FILE_31xx10x, fromRegsPortxREG_FILE_31xx9x, 
      fromRegsPortxREG_FILE_31xx8x, fromRegsPortxREG_FILE_31xx7x, 
      fromRegsPortxREG_FILE_31xx6x, fromRegsPortxREG_FILE_31xx5x, 
      fromRegsPortxREG_FILE_31xx4x, fromRegsPortxREG_FILE_31xx3x, 
      fromRegsPortxREG_FILE_31xx2x, fromRegsPortxREG_FILE_31xx1x, 
      fromRegsPortxREG_FILE_31xx0x, IF_ISAxN10974, IF_ISAxN10973, IF_ISAxN10972
      , IF_ISAxN10971, IF_ISAxN10970, IF_ISAxN10969, IF_ISAxN10968, 
      IF_ISAxN10967, IF_ISAxN10966, IF_ISAxN10965, IF_ISAxN10964, IF_ISAxN10963
      , IF_ISAxN10962, IF_ISAxN10961, IF_ISAxN10960, IF_ISAxN10959, 
      IF_ISAxN10958, IF_ISAxN10957, IF_ISAxN10956, IF_ISAxN10955, IF_ISAxN10954
      , IF_ISAxN10953, IF_ISAxN10952, IF_ISAxN10951, IF_ISAxN10950, 
      IF_ISAxN10949, IF_ISAxN10948, IF_ISAxN10947, IF_ISAxN10946, IF_ISAxN10945
      , IF_ISAxN10944, IF_ISAxN10943, IF_ISAxN10942, IF_ISAxN10941, 
      IF_ISAxN10940, IF_ISAxN10939, IF_ISAxN10938, IF_ISAxN10936, IF_ISAxN10935
      , IF_ISAxN10904, IF_ISAxN10902, IF_ISAxN10869, IF_ISAxN10868, 
      IF_ISAxN10867, IF_ISAxN10866, IF_ISAxN10865, IF_ISAxN10864, IF_ISAxN10863
      , IF_ISAxN10862, IF_ISAxN10861, IF_ISAxN10860, IF_ISAxN10859, 
      IF_ISAxN10858, IF_ISAxN10857, IF_ISAxN10856, IF_ISAxN10855, IF_ISAxN10854
      , IF_ISAxN10853, IF_ISAxN10852, IF_ISAxN10851, IF_ISAxN10850, 
      IF_ISAxN10849, IF_ISAxN10848, IF_ISAxN10847, IF_ISAxN10846, IF_ISAxN10845
      , IF_ISAxN10844, IF_ISAxN10843, IF_ISAxN10842, IF_ISAxN10832, 
      IF_ISAxN10829, IF_ISAxN2460, IF_ISAxN2459, IF_ISAxpcReg_signal_2_port, 
      IF_ISAxpcReg_signal_3_port, IF_ISAxpcReg_signal_4_port, 
      IF_ISAxpcReg_signal_5_port, IF_ISAxpcReg_signal_6_port, 
      IF_ISAxpcReg_signal_7_port, IF_ISAxpcReg_signal_8_port, 
      IF_ISAxpcReg_signal_9_port, IF_ISAxpcReg_signal_10_port, 
      IF_ISAxpcReg_signal_11_port, IF_ISAxpcReg_signal_12_port, 
      IF_ISAxpcReg_signal_13_port, IF_ISAxpcReg_signal_14_port, 
      IF_ISAxpcReg_signal_15_port, IF_ISAxpcReg_signal_16_port, 
      IF_ISAxpcReg_signal_17_port, IF_ISAxpcReg_signal_18_port, 
      IF_ISAxpcReg_signal_19_port, IF_ISAxpcReg_signal_20_port, 
      IF_ISAxpcReg_signal_21_port, IF_ISAxpcReg_signal_22_port, 
      IF_ISAxpcReg_signal_23_port, IF_ISAxpcReg_signal_24_port, 
      IF_ISAxpcReg_signal_25_port, IF_ISAxpcReg_signal_26_port, 
      IF_ISAxpcReg_signal_27_port, IF_ISAxpcReg_signal_28_port, 
      IF_ISAxpcReg_signal_29_port, IF_ISAxpcReg_signal_30_port, 
      IF_ISAxpcReg_signal_31_port, IF_ISAxsection_0_port, IF_ISAxsection_2_port
      , IF_RegsxN721, IF_RegsxN720, IF_RegsxN719, IF_RegsxN718, IF_RegsxN717, 
      IF_RegsxN716, IF_RegsxN715, IF_RegsxN714, IF_RegsxN713, IF_RegsxN712, 
      IF_RegsxN711, IF_RegsxN710, IF_RegsxN709, IF_RegsxN708, IF_RegsxN707, 
      IF_RegsxN706, IF_RegsxN705, IF_RegsxN704, IF_RegsxN703, IF_RegsxN702, 
      IF_RegsxN701, IF_RegsxN700, IF_RegsxN699, IF_RegsxN698, IF_RegsxN697, 
      IF_RegsxN696, IF_RegsxN695, IF_RegsxN694, IF_RegsxN693, IF_RegsxN692, 
      IF_RegsxN691, IF_RegsxN690, IF_RegsxN689, IF_RegsxN688, IF_RegsxN687, 
      IF_RegsxN686, IF_RegsxN685, IF_RegsxN684, IF_RegsxN683, IF_RegsxN682, 
      IF_RegsxN681, IF_RegsxN680, IF_RegsxN679, IF_RegsxN678, IF_RegsxN677, 
      IF_RegsxN676, IF_RegsxN675, IF_RegsxN674, IF_RegsxN673, IF_RegsxN672, 
      IF_RegsxN671, IF_RegsxN670, IF_RegsxN669, IF_RegsxN668, IF_RegsxN667, 
      IF_RegsxN666, IF_RegsxN665, IF_RegsxN664, IF_RegsxN663, IF_RegsxN662, 
      IF_RegsxN661, IF_RegsxN660, IF_RegsxN659, net325226, net325231, net325236
      , net325241, net325246, net325251, net325256, net325261, net325266, 
      net325271, net325276, net325281, net325286, net325291, net325296, 
      net325301, net325306, net325311, net325316, net325321, net325326, 
      net325331, net325336, net325341, net325346, net325351, net325356, 
      net325361, net325366, net325371, net325376, net325381, net325386, 
      net325391, net325396, net325401, net325406, ashr_25xAx30x, ashr_25xAx29x,
      ashr_25xAx28x, ashr_25xAx27x, ashr_25xAx26x, ashr_25xAx25x, ashr_25xAx24x
      , ashr_25xAx23x, ashr_25xAx22x, ashr_25xAx21x, ashr_25xAx20x, 
      ashr_25xAx19x, ashr_25xAx18x, ashr_25xAx17x, ashr_25xAx16x, ashr_25xAx15x
      , ashr_25xAx14x, ashr_25xAx13x, ashr_25xAx12x, ashr_25xAx11x, 
      ashr_25xAx10x, ashr_25xAx9x, ashr_25xAx8x, ashr_25xAx7x, ashr_25xAx6x, 
      ashr_25xAx5x, ashr_25xAx4x, ashr_25xAx3x, ashr_25xAx2x, ashr_25xAx1x, 
      ashr_25xAx0x, ashr_25xSHx4x, ashr_25xSHx3x, n3458, add_x_26xBx30x, 
      add_x_26xBx29x, add_x_26xBx28x, add_x_26xBx27x, add_x_26xBx26x, 
      add_x_26xBx25x, add_x_26xBx24x, add_x_26xBx23x, add_x_26xBx22x, 
      add_x_26xBx21x, add_x_26xBx20x, add_x_26xBx19x, add_x_26xBx18x, 
      add_x_26xBx17x, add_x_26xBx16x, add_x_26xBx15x, add_x_26xBx14x, 
      add_x_26xBx13x, add_x_26xBx12x, add_x_26xBx11x, add_x_26xBx10x, 
      add_x_26xBx9x, add_x_26xBx8x, add_x_26xBx7x, add_x_26xBx6x, add_x_26xBx5x
      , DP_OP_679J14_122_3096xn99, DP_OP_679J14_122_3096xn98, 
      DP_OP_679J14_122_3096xn97, DP_OP_679J14_122_3096xn96, 
      DP_OP_679J14_122_3096xn95, DP_OP_679J14_122_3096xn94, 
      DP_OP_679J14_122_3096xn93, DP_OP_679J14_122_3096xn92, 
      DP_OP_679J14_122_3096xn91, DP_OP_679J14_122_3096xn90, 
      DP_OP_679J14_122_3096xn89, DP_OP_679J14_122_3096xn88, 
      DP_OP_679J14_122_3096xn87, DP_OP_679J14_122_3096xn86, 
      DP_OP_679J14_122_3096xn85, DP_OP_679J14_122_3096xn84, 
      DP_OP_679J14_122_3096xn83, DP_OP_679J14_122_3096xn82, 
      DP_OP_679J14_122_3096xn81, DP_OP_679J14_122_3096xn80, 
      DP_OP_679J14_122_3096xn79, DP_OP_679J14_122_3096xn78, 
      DP_OP_679J14_122_3096xn77, DP_OP_679J14_122_3096xn76, 
      DP_OP_679J14_122_3096xn75, DP_OP_679J14_122_3096xn74, 
      DP_OP_679J14_122_3096xn73, DP_OP_679J14_122_3096xn72, 
      DP_OP_679J14_122_3096xn71, DP_OP_679J14_122_3096xn70, 
      DP_OP_679J14_122_3096xn69, DP_OP_679J14_122_3096xn68, 
      DP_OP_679J14_122_3096xn67, DP_OP_679J14_122_3096xn66, 
      DP_OP_679J14_122_3096xn65, DP_OP_679J14_122_3096xn64, 
      DP_OP_679J14_122_3096xn63, DP_OP_679J14_122_3096xn62, 
      DP_OP_679J14_122_3096xn61, DP_OP_679J14_122_3096xn60, 
      DP_OP_679J14_122_3096xn59, DP_OP_679J14_122_3096xn58, 
      DP_OP_679J14_122_3096xn57, DP_OP_679J14_122_3096xn56, 
      DP_OP_679J14_122_3096xn55, DP_OP_679J14_122_3096xn54, 
      DP_OP_679J14_122_3096xn53, DP_OP_679J14_122_3096xn52, 
      DP_OP_679J14_122_3096xn51, DP_OP_679J14_122_3096xn50, 
      DP_OP_679J14_122_3096xn49, DP_OP_679J14_122_3096xn48, 
      DP_OP_679J14_122_3096xn47, DP_OP_679J14_122_3096xn46, 
      DP_OP_679J14_122_3096xn45, DP_OP_679J14_122_3096xn44, 
      DP_OP_679J14_122_3096xn43, DP_OP_679J14_122_3096xn42, 
      DP_OP_679J14_122_3096xn41, DP_OP_679J14_122_3096xn40, 
      DP_OP_679J14_122_3096xn39, DP_OP_679J14_122_3096xn38, 
      DP_OP_679J14_122_3096xn32, DP_OP_679J14_122_3096xn31, 
      DP_OP_679J14_122_3096xn30, DP_OP_679J14_122_3096xn29, 
      DP_OP_679J14_122_3096xn28, DP_OP_679J14_122_3096xn27, 
      DP_OP_679J14_122_3096xn26, DP_OP_679J14_122_3096xn25, 
      DP_OP_679J14_122_3096xn24, DP_OP_679J14_122_3096xn23, 
      DP_OP_679J14_122_3096xn22, DP_OP_679J14_122_3096xn21, 
      DP_OP_679J14_122_3096xn20, DP_OP_679J14_122_3096xn19, 
      DP_OP_679J14_122_3096xn18, DP_OP_679J14_122_3096xn17, 
      DP_OP_679J14_122_3096xn16, DP_OP_679J14_122_3096xn15, 
      DP_OP_679J14_122_3096xn14, DP_OP_679J14_122_3096xn13, 
      DP_OP_679J14_122_3096xn12, DP_OP_679J14_122_3096xn11, 
      DP_OP_679J14_122_3096xn10, DP_OP_679J14_122_3096xn9, 
      DP_OP_679J14_122_3096xn8, DP_OP_679J14_122_3096xn7, 
      DP_OP_679J14_122_3096xn6, DP_OP_679J14_122_3096xn5, 
      DP_OP_679J14_122_3096xn4, DP_OP_679J14_122_3096xn3, 
      DP_OP_679J14_122_3096xn2, DP_OP_719J14_125_1055xn164, 
      DP_OP_719J14_125_1055xn163, DP_OP_719J14_125_1055xn162, 
      DP_OP_719J14_125_1055xn161, DP_OP_719J14_125_1055xn160, 
      DP_OP_719J14_125_1055xn159, DP_OP_719J14_125_1055xn158, 
      DP_OP_719J14_125_1055xn157, DP_OP_719J14_125_1055xn156, 
      DP_OP_719J14_125_1055xn155, DP_OP_719J14_125_1055xn154, 
      DP_OP_719J14_125_1055xn153, DP_OP_719J14_125_1055xn152, 
      DP_OP_719J14_125_1055xn151, DP_OP_719J14_125_1055xn150, 
      DP_OP_719J14_125_1055xn149, DP_OP_719J14_125_1055xn148, 
      DP_OP_719J14_125_1055xn147, DP_OP_719J14_125_1055xn146, 
      DP_OP_719J14_125_1055xn145, DP_OP_719J14_125_1055xn144, 
      DP_OP_719J14_125_1055xn143, DP_OP_719J14_125_1055xn142, 
      DP_OP_719J14_125_1055xn141, DP_OP_719J14_125_1055xn140, 
      DP_OP_719J14_125_1055xn139, DP_OP_719J14_125_1055xn138, 
      DP_OP_719J14_125_1055xn137, DP_OP_719J14_125_1055xn136, 
      DP_OP_719J14_125_1055xn135, DP_OP_719J14_125_1055xn134, 
      DP_OP_719J14_125_1055xn99, DP_OP_719J14_125_1055xn98, 
      DP_OP_719J14_125_1055xn97, DP_OP_719J14_125_1055xn96, 
      DP_OP_719J14_125_1055xn95, DP_OP_719J14_125_1055xn94, 
      DP_OP_719J14_125_1055xn93, DP_OP_719J14_125_1055xn92, 
      DP_OP_719J14_125_1055xn91, DP_OP_719J14_125_1055xn90, 
      DP_OP_719J14_125_1055xn89, DP_OP_719J14_125_1055xn88, 
      DP_OP_719J14_125_1055xn87, DP_OP_719J14_125_1055xn86, 
      DP_OP_719J14_125_1055xn85, DP_OP_719J14_125_1055xn84, 
      DP_OP_719J14_125_1055xn83, DP_OP_719J14_125_1055xn82, 
      DP_OP_719J14_125_1055xn81, DP_OP_719J14_125_1055xn80, 
      DP_OP_719J14_125_1055xn79, DP_OP_719J14_125_1055xn78, 
      DP_OP_719J14_125_1055xn77, DP_OP_719J14_125_1055xn76, 
      DP_OP_719J14_125_1055xn75, DP_OP_719J14_125_1055xn74, 
      DP_OP_719J14_125_1055xn73, DP_OP_719J14_125_1055xn72, 
      DP_OP_719J14_125_1055xn71, DP_OP_719J14_125_1055xn70, 
      DP_OP_719J14_125_1055xn69, DP_OP_719J14_125_1055xn68, 
      DP_OP_719J14_125_1055xn67, DP_OP_719J14_125_1055xn66, 
      DP_OP_719J14_125_1055xn65, DP_OP_719J14_125_1055xn64, 
      DP_OP_719J14_125_1055xn63, DP_OP_719J14_125_1055xn62, 
      DP_OP_719J14_125_1055xn61, DP_OP_719J14_125_1055xn60, 
      DP_OP_719J14_125_1055xn59, DP_OP_719J14_125_1055xn58, 
      DP_OP_719J14_125_1055xn57, DP_OP_719J14_125_1055xn56, 
      DP_OP_719J14_125_1055xn55, DP_OP_719J14_125_1055xn54, 
      DP_OP_719J14_125_1055xn53, DP_OP_719J14_125_1055xn52, 
      DP_OP_719J14_125_1055xn51, DP_OP_719J14_125_1055xn50, 
      DP_OP_719J14_125_1055xn49, DP_OP_719J14_125_1055xn48, 
      DP_OP_719J14_125_1055xn47, DP_OP_719J14_125_1055xn46, 
      DP_OP_719J14_125_1055xn45, DP_OP_719J14_125_1055xn44, 
      DP_OP_719J14_125_1055xn43, DP_OP_719J14_125_1055xn42, 
      DP_OP_719J14_125_1055xn41, DP_OP_719J14_125_1055xn40, 
      DP_OP_719J14_125_1055xn39, DP_OP_719J14_125_1055xn38, 
      DP_OP_719J14_125_1055xn32, DP_OP_719J14_125_1055xn31, 
      DP_OP_719J14_125_1055xn30, DP_OP_719J14_125_1055xn29, 
      DP_OP_719J14_125_1055xn28, DP_OP_719J14_125_1055xn27, 
      DP_OP_719J14_125_1055xn26, DP_OP_719J14_125_1055xn25, 
      DP_OP_719J14_125_1055xn24, DP_OP_719J14_125_1055xn23, 
      DP_OP_719J14_125_1055xn22, DP_OP_719J14_125_1055xn21, 
      DP_OP_719J14_125_1055xn20, DP_OP_719J14_125_1055xn19, 
      DP_OP_719J14_125_1055xn18, DP_OP_719J14_125_1055xn17, 
      DP_OP_719J14_125_1055xn16, DP_OP_719J14_125_1055xn15, 
      DP_OP_719J14_125_1055xn14, DP_OP_719J14_125_1055xn13, 
      DP_OP_719J14_125_1055xn12, DP_OP_719J14_125_1055xn11, 
      DP_OP_719J14_125_1055xn10, DP_OP_719J14_125_1055xn9, 
      DP_OP_719J14_125_1055xn8, DP_OP_719J14_125_1055xn7, 
      DP_OP_719J14_125_1055xn6, DP_OP_719J14_125_1055xn5, 
      DP_OP_719J14_125_1055xn4, DP_OP_719J14_125_1055xn3, 
      DP_OP_719J14_125_1055xn2, intadd_25xBx0x, intadd_25xCI, intadd_25xSUMx28x
      , intadd_25xSUMx27x, intadd_25xSUMx26x, intadd_25xSUMx25x, 
      intadd_25xSUMx24x, intadd_25xSUMx23x, intadd_25xSUMx22x, 
      intadd_25xSUMx21x, intadd_25xSUMx20x, intadd_25xSUMx19x, 
      intadd_25xSUMx18x, intadd_25xSUMx17x, intadd_25xSUMx16x, 
      intadd_25xSUMx15x, intadd_25xSUMx14x, intadd_25xSUMx13x, 
      intadd_25xSUMx12x, intadd_25xSUMx11x, intadd_25xSUMx10x, intadd_25xSUMx9x
      , intadd_25xSUMx8x, intadd_25xSUMx7x, intadd_25xSUMx6x, intadd_25xSUMx5x,
      intadd_25xSUMx4x, intadd_25xSUMx3x, intadd_25xSUMx2x, intadd_25xSUMx1x, 
      intadd_25xSUMx0x, intadd_25xn29, intadd_25xn28, intadd_25xn27, 
      intadd_25xn26, intadd_25xn25, intadd_25xn24, intadd_25xn23, intadd_25xn22
      , intadd_25xn21, intadd_25xn20, intadd_25xn19, intadd_25xn18, 
      intadd_25xn17, intadd_25xn16, intadd_25xn15, intadd_25xn14, intadd_25xn13
      , intadd_25xn12, intadd_25xn11, intadd_25xn10, intadd_25xn9, intadd_25xn8
      , intadd_25xn7, intadd_25xn6, intadd_25xn5, intadd_25xn4, intadd_25xn3, 
      intadd_25xn2, intadd_25xn1, intadd_26xAx7x, intadd_26xAx6x, 
      intadd_26xAx5x, intadd_26xAx4x, intadd_26xAx3x, intadd_26xAx2x, 
      intadd_26xAx1x, intadd_26xAx0x, intadd_26xBx7x, intadd_26xBx6x, 
      intadd_26xBx5x, intadd_26xBx4x, intadd_26xBx3x, intadd_26xBx2x, 
      intadd_26xBx1x, intadd_26xBx0x, intadd_26xCI, intadd_26xSUMx7x, 
      intadd_26xSUMx6x, intadd_26xSUMx5x, intadd_26xSUMx4x, intadd_26xSUMx3x, 
      intadd_26xSUMx2x, intadd_26xSUMx1x, intadd_26xSUMx0x, intadd_26xn8, 
      intadd_26xn7, intadd_26xn6, intadd_26xn5, intadd_26xn4, intadd_26xn3, 
      intadd_26xn2, intadd_26xn1, intadd_27xAx3x, intadd_27xAx2x, 
      intadd_27xAx1x, intadd_27xAx0x, intadd_27xBx3x, intadd_27xBx2x, 
      intadd_27xBx1x, intadd_27xBx0x, intadd_27xCI, intadd_27xSUMx3x, 
      intadd_27xSUMx2x, intadd_27xSUMx1x, intadd_27xSUMx0x, intadd_27xn4, 
      intadd_27xn3, intadd_27xn2, intadd_27xn1, intadd_28xAx2x, intadd_28xAx1x,
      intadd_28xAx0x, intadd_28xBx2x, intadd_28xBx1x, intadd_28xBx0x, 
      intadd_28xCI, intadd_28xSUMx2x, intadd_28xSUMx1x, intadd_28xSUMx0x, 
      intadd_28xn3, intadd_28xn2, intadd_28xn1, intadd_29xAx2x, intadd_29xAx1x,
      intadd_29xAx0x, intadd_29xBx2x, intadd_29xBx1x, intadd_29xBx0x, 
      intadd_29xCI, intadd_29xSUMx2x, intadd_29xSUMx1x, intadd_29xSUMx0x, 
      intadd_29xn3, intadd_29xn2, intadd_29xn1, n3558, n3559, n3560, n3561, 
      n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, 
      n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, 
      n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, 
      n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, 
      n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, 
      n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, 
      n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, 
      n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, 
      n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, 
      n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, 
      n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, 
      n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, 
      n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, 
      n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, 
      n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, 
      n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, 
      n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, 
      n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, 
      n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, 
      n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, 
      n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, 
      n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, 
      n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, 
      n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, 
      n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, 
      n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, 
      n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, 
      n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, 
      n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, 
      n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, 
      n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, 
      n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, 
      n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, 
      n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, 
      n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, 
      n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, 
      n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, 
      n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, 
      n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, 
      n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, 
      n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, 
      n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, 
      n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, 
      n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, 
      n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, 
      n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, 
      n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, 
      n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, 
      n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, 
      n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, 
      n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, 
      n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, 
      n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, 
      n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, 
      n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, 
      n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, 
      n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, 
      n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, 
      n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, 
      n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, 
      n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, 
      n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, 
      n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, 
      n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, 
      n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, 
      n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, 
      n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, 
      n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, 
      n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, 
      n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, 
      n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, 
      n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, 
      n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, 
      n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, 
      n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, 
      n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, 
      n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, 
      n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, 
      n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, 
      n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, 
      n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, 
      n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, 
      n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, 
      n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, 
      n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, 
      n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, 
      n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, 
      n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, 
      n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, 
      n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, 
      n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, 
      n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, 
      n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, 
      n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, 
      n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, 
      n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, 
      n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, 
      n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, 
      n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, 
      n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, 
      n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, 
      n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, 
      n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, 
      n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, 
      n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, 
      n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, 
      n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, 
      n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, 
      n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, 
      n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, 
      n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, 
      n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, 
      n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, 
      n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, 
      n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, 
      n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, 
      n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, 
      n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, 
      n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, 
      n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, 
      n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, 
      n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, 
      n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, 
      n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, 
      n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, 
      n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, 
      n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, 
      n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, 
      n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, 
      n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, 
      n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, 
      n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, 
      n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, 
      n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, 
      n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, 
      n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, 
      n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, 
      n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, 
      n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, 
      n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, 
      n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, 
      n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, 
      n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, 
      n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, 
      n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, 
      n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, 
      n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, 
      n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, 
      n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, 
      n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, 
      n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, 
      n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, 
      n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, 
      n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, 
      n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, 
      n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, 
      n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, 
      n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, 
      n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, 
      n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, 
      n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, 
      n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, 
      n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, 
      n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, 
      n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, 
      n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, 
      n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, 
      n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, 
      n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, 
      n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, 
      n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, 
      n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, 
      n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, 
      n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, 
      n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, 
      n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, 
      n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, 
      n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, 
      n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, 
      n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, 
      n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, 
      n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, 
      n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, 
      n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, 
      n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, 
      n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, 
      n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, 
      n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, 
      n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, 
      n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, 
      n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, 
      n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, 
      n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, 
      n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, 
      n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, 
      n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, 
      n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, 
      n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, 
      n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, 
      n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, 
      n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, 
      n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, 
      n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, 
      n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, 
      n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, 
      n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, 
      n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, 
      n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, 
      n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, 
      n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, 
      n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, 
      n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, 
      n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, 
      n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, 
      n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, 
      n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, 
      n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, 
      n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, 
      n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, 
      n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, 
      n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, 
      n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, 
      n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, 
      n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, 
      n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, 
      n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, 
      n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, 
      n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, 
      n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, 
      n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, 
      n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, 
      n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, 
      n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, 
      n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, 
      n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, 
      n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, 
      n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, 
      n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, 
      n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, 
      n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, 
      n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, 
      n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, 
      n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, 
      n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, 
      n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, 
      n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, 
      n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, 
      n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, 
      n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, 
      n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, 
      n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, 
      n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, 
      n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, 
      n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, 
      n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, 
      n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, 
      n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, 
      n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, 
      n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, 
      n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, 
      n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, 
      n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, 
      n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, 
      n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, 
      n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, 
      n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, 
      n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, 
      n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, 
      n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, 
      n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, 
      n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, 
      n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, 
      n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, 
      n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, 
      n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, 
      n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, 
      n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, 
      n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, 
      n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, 
      n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, 
      n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, 
      n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, 
      n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, 
      n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, 
      n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, 
      n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, 
      n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, 
      n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, 
      n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, 
      n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, 
      n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, 
      n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, 
      n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, 
      n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, 
      n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, 
      n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, 
      n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, 
      n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, 
      n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, 
      n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, 
      n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, 
      n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, 
      n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, 
      n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, 
      n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, 
      n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, 
      n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, 
      n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, 
      n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, 
      n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, 
      n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, 
      n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, 
      n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, 
      n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, 
      n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, 
      n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, 
      n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, 
      n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, 
      n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, 
      n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, 
      n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, 
      n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, 
      n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, 
      n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, 
      n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, 
      n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, 
      n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, 
      n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, 
      n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, 
      n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, 
      n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, 
      n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, 
      n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, 
      n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, 
      n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, 
      n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, 
      n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, 
      n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, 
      n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, 
      n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, 
      n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, 
      n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, 
      n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, 
      n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, 
      n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, 
      n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, 
      n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, 
      n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, 
      n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, 
      n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, 
      n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, 
      n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, 
      n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, 
      n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, 
      n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, 
      n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, 
      n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, 
      n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, 
      n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, 
      n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, 
      n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, 
      n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, 
      n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, 
      n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, 
      n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, 
      n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, 
      n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, 
      n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, 
      n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, 
      n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, 
      n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, 
      n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, 
      n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, 
      n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, 
      n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, 
      n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, 
      n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, 
      n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, 
      n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, 
      n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, 
      n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, 
      n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, 
      n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, 
      n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, 
      n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, 
      n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, 
      n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, 
      n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, 
      n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, 
      n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, 
      n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, 
      n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, 
      n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, 
      n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, 
      n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, 
      n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, 
      n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, 
      n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, 
      n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, 
      n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, 
      n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, 
      n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, 
      n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, 
      n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, 
      n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, 
      n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, 
      n7622, n7623, n7624, n7625, n7626, n7628, n_1000, n_1001, n_1002, n_1003,
      n_1004, n_1005, n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, 
      n_1013, n_1014, n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, 
      n_1022, n_1023, n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, 
      n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, 
      n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, 
      n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, 
      n_1058, n_1059, n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, 
      n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, 
      n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, 
      n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, 
      n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, 
      n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, 
      n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, 
      n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, 
      n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, 
      n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, 
      n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, 
      n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, 
      n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, 
      n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, 
      n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, 
      n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, 
      n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, 
      n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, 
      n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, 
      n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, 
      n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, 
      n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, 
      n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, 
      n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, 
      n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, 
      n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, 
      n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, 
      n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, 
      n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, 
      n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, 
      n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, 
      n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, 
      n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, 
      n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, 
      n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, 
      n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, 
      n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, 
      n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, 
      n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, 
      n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, 
      n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, 
      n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, 
      n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, 
      n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, 
      n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, 
      n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, 
      n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, 
      n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, 
      n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, 
      n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, 
      n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, 
      n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, 
      n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, 
      n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, 
      n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, 
      n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, 
      n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, 
      n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, 
      n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, 
      n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, 
      n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, 
      n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, 
      n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, 
      n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, 
      n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, 
      n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, 
      n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, 
      n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, 
      n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, 
      n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, 
      n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, 
      n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, 
      n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, 
      n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, 
      n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, 
      n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, 
      n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, 
      n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, 
      n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, 
      n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, 
      n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, 
      n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, 
      n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, 
      n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, 
      n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, 
      n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, 
      n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, 
      n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, 
      n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, 
      n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, 
      n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, 
      n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, 
      n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, 
      n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, 
      n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, 
      n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, 
      n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, 
      n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, 
      n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, 
      n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, 
      n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, 
      n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, 
      n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, 
      n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, 
      n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, 
      n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, 
      n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, 
      n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, 
      n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, 
      n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, 
      n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, 
      n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, 
      n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, 
      n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, 
      n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, 
      n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, 
      n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, 
      n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118 : 
      std_logic;

begin
   fromMemoryPort_sync_port <= bool_to_std_logic(fromMemoryPort_sync);
   fromMemoryPort_notify <= std_logic_to_bool(IF_ISAxsection_0_port);
   toMemoryPort_sync_port <= bool_to_std_logic(toMemoryPort_sync);
   toMemoryPort_notify <= std_logic_to_bool(toMemoryPort_notify_port);
   
   IF_ISAxsection_regx2x : DFF_X1 port map( D => n7555, CK => net325226, Q => 
                           IF_ISAxsection_2_port, QN => n7535);
   IF_ISAxsection_regx1x : DFF_X1 port map( D => n7554, CK => net325226, Q => 
                           n_1000, QN => n7538);
   IF_ISAxtoRegsPort_regxDSTxx0x : DFF_X1 port map( D => IF_ISAxN10970, CK => 
                           net325236, Q => toRegsPortxDSTxx0x, QN => n7536);
   IF_ISAxtoRegsPort_regxDSTxx1x : DFF_X1 port map( D => IF_ISAxN10971, CK => 
                           net325236, Q => toRegsPortxDSTxx1x, QN => n7534);
   IF_ISAxtoRegsPort_regxDSTxx2x : DFF_X1 port map( D => IF_ISAxN10972, CK => 
                           net325236, Q => toRegsPortxDSTxx2x, QN => n7537);
   IF_ISAxtoRegsPort_regxDSTxx3x : DFF_X1 port map( D => IF_ISAxN10973, CK => 
                           net325236, Q => toRegsPortxDSTxx3x, QN => n7541);
   IF_ISAxtoRegsPort_regxDSTxx4x : DFF_X1 port map( D => IF_ISAxN10974, CK => 
                           net325236, Q => toRegsPortxDSTxx4x, QN => n7539);
   IF_ISAxsection_regx0x : DFF_X1 port map( D => n7556, CK => net325226, Q => 
                           IF_ISAxsection_0_port, QN => n_1001);
   IF_ISAxpcReg_signal_regx0x : DFF_X1 port map( D => n7552, CK => net325241, Q
                           => IF_ISAxN2459, QN => n7549);
   IF_ISAxpcReg_signal_regx1x : DFF_X1 port map( D => IF_ISAxN10904, CK => 
                           net325241, Q => IF_ISAxN2460, QN => n7542);
   IF_ISAxpcReg_signal_regx2x : DFF_X1 port map( D => n7586, CK => net325241, Q
                           => IF_ISAxpcReg_signal_2_port, QN => n7546);
   IF_ISAxpcReg_signal_regx3x : DFF_X1 port map( D => n7585, CK => net325241, Q
                           => IF_ISAxpcReg_signal_3_port, QN => n_1002);
   IF_ISAxpcReg_signal_regx4x : DFF_X1 port map( D => n7584, CK => net325241, Q
                           => IF_ISAxpcReg_signal_4_port, QN => n_1003);
   IF_ISAxpcReg_signal_regx5x : DFF_X1 port map( D => n7583, CK => net325241, Q
                           => IF_ISAxpcReg_signal_5_port, QN => n_1004);
   IF_ISAxpcReg_signal_regx6x : DFF_X1 port map( D => n7582, CK => net325241, Q
                           => IF_ISAxpcReg_signal_6_port, QN => n7543);
   IF_ISAxpcReg_signal_regx7x : DFF_X1 port map( D => n7581, CK => net325241, Q
                           => IF_ISAxpcReg_signal_7_port, QN => n_1005);
   IF_ISAxpcReg_signal_regx8x : DFF_X1 port map( D => n7580, CK => net325241, Q
                           => IF_ISAxpcReg_signal_8_port, QN => n7544);
   IF_ISAxpcReg_signal_regx9x : DFF_X1 port map( D => n7579, CK => net325241, Q
                           => IF_ISAxpcReg_signal_9_port, QN => n_1006);
   IF_ISAxpcReg_signal_regx10x : DFF_X1 port map( D => n7578, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_10_port, QN => n7545);
   IF_ISAxpcReg_signal_regx11x : DFF_X1 port map( D => n7577, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_11_port, QN => n_1007);
   IF_ISAxpcReg_signal_regx12x : DFF_X1 port map( D => n7576, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_12_port, QN => n7547);
   IF_ISAxpcReg_signal_regx13x : DFF_X1 port map( D => n7575, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_13_port, QN => n_1008);
   IF_ISAxpcReg_signal_regx14x : DFF_X1 port map( D => n7574, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_14_port, QN => n_1009);
   IF_ISAxpcReg_signal_regx15x : DFF_X1 port map( D => n7573, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_15_port, QN => n_1010);
   IF_ISAxpcReg_signal_regx16x : DFF_X1 port map( D => n7572, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_16_port, QN => n_1011);
   IF_ISAxpcReg_signal_regx17x : DFF_X1 port map( D => n7571, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_17_port, QN => n_1012);
   IF_ISAxpcReg_signal_regx18x : DFF_X1 port map( D => n7570, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_18_port, QN => n_1013);
   IF_ISAxpcReg_signal_regx19x : DFF_X1 port map( D => n7569, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_19_port, QN => n_1014);
   IF_ISAxpcReg_signal_regx20x : DFF_X1 port map( D => n7568, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_20_port, QN => n_1015);
   IF_ISAxpcReg_signal_regx21x : DFF_X1 port map( D => n7567, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_21_port, QN => n_1016);
   IF_ISAxpcReg_signal_regx22x : DFF_X1 port map( D => n7566, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_22_port, QN => n_1017);
   IF_ISAxpcReg_signal_regx23x : DFF_X1 port map( D => n7565, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_23_port, QN => n_1018);
   IF_ISAxpcReg_signal_regx24x : DFF_X1 port map( D => n7564, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_24_port, QN => n_1019);
   IF_ISAxpcReg_signal_regx25x : DFF_X1 port map( D => n7563, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_25_port, QN => n_1020);
   IF_ISAxpcReg_signal_regx26x : DFF_X1 port map( D => n7562, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_26_port, QN => n_1021);
   IF_ISAxpcReg_signal_regx27x : DFF_X1 port map( D => n7561, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_27_port, QN => n_1022);
   IF_ISAxpcReg_signal_regx28x : DFF_X1 port map( D => n7560, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_28_port, QN => n_1023);
   IF_ISAxpcReg_signal_regx29x : DFF_X1 port map( D => n7559, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_29_port, QN => n_1024);
   IF_ISAxpcReg_signal_regx30x : DFF_X1 port map( D => n7558, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_30_port, QN => n_1025);
   IF_ISAxpcReg_signal_regx31x : DFF_X1 port map( D => n7557, CK => net325241, 
                           Q => IF_ISAxpcReg_signal_31_port, QN => n7548);
   IF_ISAxtoMemoryPort_regxREQxx0x : DFF_X1 port map( D => n7595, CK => 
                           net325246, Q => toMemoryPortxREQxx0x(0), QN => 
                           n_1026);
   IF_ISAxtoMemoryPort_regxMASKxx0x : DFF_X1 port map( D => n7594, CK => 
                           net325246, Q => toMemoryPortxMASKxx0x(0), QN => 
                           n_1027);
   IF_ISAxtoMemoryPort_regxMASKxx1x : DFF_X1 port map( D => n7593, CK => 
                           net325246, Q => toMemoryPortxMASKxx1x(0), QN => 
                           n_1028);
   IF_ISAxtoMemoryPort_regxMASKxx2x : DFF_X1 port map( D => n7592, CK => 
                           net325246, Q => toMemoryPortxMASKxx2x(0), QN => 
                           n_1029);
   IF_ISAxtoMemoryPort_regxADDRINxx0x : DFF_X1 port map( D => n7552, CK => 
                           net325251, Q => toMemoryPortxADDRINxx0x(0), QN => 
                           n_1030);
   IF_ISAxtoMemoryPort_regxADDRINxx1x : DFF_X1 port map( D => n7626, CK => 
                           net325251, Q => toMemoryPortxADDRINxx1x(0), QN => 
                           n_1031);
   IF_ISAxtoMemoryPort_regxADDRINxx2x : DFF_X1 port map( D => n7625, CK => 
                           net325251, Q => toMemoryPortxADDRINxx2x(0), QN => 
                           n_1032);
   IF_ISAxtoMemoryPort_regxADDRINxx3x : DFF_X1 port map( D => n7624, CK => 
                           net325251, Q => toMemoryPortxADDRINxx3x(0), QN => 
                           n_1033);
   IF_ISAxtoMemoryPort_regxADDRINxx4x : DFF_X1 port map( D => n7623, CK => 
                           net325251, Q => toMemoryPortxADDRINxx4x(0), QN => 
                           n_1034);
   IF_ISAxtoMemoryPort_regxADDRINxx5x : DFF_X1 port map( D => n7622, CK => 
                           net325251, Q => toMemoryPortxADDRINxx5x(0), QN => 
                           n_1035);
   IF_ISAxtoMemoryPort_regxADDRINxx6x : DFF_X1 port map( D => n7621, CK => 
                           net325251, Q => toMemoryPortxADDRINxx6x(0), QN => 
                           n_1036);
   IF_ISAxtoMemoryPort_regxADDRINxx7x : DFF_X1 port map( D => n7620, CK => 
                           net325251, Q => toMemoryPortxADDRINxx7x(0), QN => 
                           n_1037);
   IF_ISAxtoMemoryPort_regxADDRINxx8x : DFF_X1 port map( D => n7619, CK => 
                           net325251, Q => toMemoryPortxADDRINxx8x(0), QN => 
                           n_1038);
   IF_ISAxtoMemoryPort_regxADDRINxx9x : DFF_X1 port map( D => n7618, CK => 
                           net325251, Q => toMemoryPortxADDRINxx9x(0), QN => 
                           n_1039);
   IF_ISAxtoMemoryPort_regxADDRINxx10x : DFF_X1 port map( D => n7617, CK => 
                           net325251, Q => toMemoryPortxADDRINxx10x(0), QN => 
                           n_1040);
   IF_ISAxtoMemoryPort_regxADDRINxx11x : DFF_X1 port map( D => n7616, CK => 
                           net325251, Q => toMemoryPortxADDRINxx11x(0), QN => 
                           n_1041);
   IF_ISAxtoMemoryPort_regxADDRINxx12x : DFF_X1 port map( D => n7615, CK => 
                           net325251, Q => toMemoryPortxADDRINxx12x(0), QN => 
                           n_1042);
   IF_ISAxtoMemoryPort_regxADDRINxx13x : DFF_X1 port map( D => n7614, CK => 
                           net325251, Q => toMemoryPortxADDRINxx13x(0), QN => 
                           n_1043);
   IF_ISAxtoMemoryPort_regxADDRINxx14x : DFF_X1 port map( D => n7613, CK => 
                           net325251, Q => toMemoryPortxADDRINxx14x(0), QN => 
                           n_1044);
   IF_ISAxtoMemoryPort_regxADDRINxx15x : DFF_X1 port map( D => n7612, CK => 
                           net325251, Q => toMemoryPortxADDRINxx15x(0), QN => 
                           n_1045);
   IF_ISAxtoMemoryPort_regxADDRINxx16x : DFF_X1 port map( D => n7611, CK => 
                           net325251, Q => toMemoryPortxADDRINxx16x(0), QN => 
                           n_1046);
   IF_ISAxtoMemoryPort_regxADDRINxx17x : DFF_X1 port map( D => n7610, CK => 
                           net325251, Q => toMemoryPortxADDRINxx17x(0), QN => 
                           n_1047);
   IF_ISAxtoMemoryPort_regxADDRINxx18x : DFF_X1 port map( D => n7609, CK => 
                           net325251, Q => toMemoryPortxADDRINxx18x(0), QN => 
                           n_1048);
   IF_ISAxtoMemoryPort_regxADDRINxx19x : DFF_X1 port map( D => n7608, CK => 
                           net325251, Q => toMemoryPortxADDRINxx19x(0), QN => 
                           n_1049);
   IF_ISAxtoMemoryPort_regxADDRINxx20x : DFF_X1 port map( D => n7607, CK => 
                           net325251, Q => toMemoryPortxADDRINxx20x(0), QN => 
                           n_1050);
   IF_ISAxtoMemoryPort_regxADDRINxx21x : DFF_X1 port map( D => n7606, CK => 
                           net325251, Q => toMemoryPortxADDRINxx21x(0), QN => 
                           n_1051);
   IF_ISAxtoMemoryPort_regxADDRINxx22x : DFF_X1 port map( D => n7605, CK => 
                           net325251, Q => toMemoryPortxADDRINxx22x(0), QN => 
                           n_1052);
   IF_ISAxtoMemoryPort_regxADDRINxx23x : DFF_X1 port map( D => n7604, CK => 
                           net325251, Q => toMemoryPortxADDRINxx23x(0), QN => 
                           n_1053);
   IF_ISAxtoMemoryPort_regxADDRINxx24x : DFF_X1 port map( D => n7603, CK => 
                           net325251, Q => toMemoryPortxADDRINxx24x(0), QN => 
                           n_1054);
   IF_ISAxtoMemoryPort_regxADDRINxx25x : DFF_X1 port map( D => n7602, CK => 
                           net325251, Q => toMemoryPortxADDRINxx25x(0), QN => 
                           n_1055);
   IF_ISAxtoMemoryPort_regxADDRINxx26x : DFF_X1 port map( D => n7601, CK => 
                           net325251, Q => toMemoryPortxADDRINxx26x(0), QN => 
                           n_1056);
   IF_ISAxtoMemoryPort_regxADDRINxx27x : DFF_X1 port map( D => n7600, CK => 
                           net325251, Q => toMemoryPortxADDRINxx27x(0), QN => 
                           n_1057);
   IF_ISAxtoMemoryPort_regxADDRINxx28x : DFF_X1 port map( D => n7599, CK => 
                           net325251, Q => toMemoryPortxADDRINxx28x(0), QN => 
                           n_1058);
   IF_ISAxtoMemoryPort_regxADDRINxx29x : DFF_X1 port map( D => n7598, CK => 
                           net325251, Q => toMemoryPortxADDRINxx29x(0), QN => 
                           n_1059);
   IF_ISAxtoMemoryPort_regxADDRINxx30x : DFF_X1 port map( D => n7597, CK => 
                           net325251, Q => toMemoryPortxADDRINxx30x(0), QN => 
                           n_1060);
   IF_ISAxtoMemoryPort_regxADDRINxx31x : DFF_X1 port map( D => n7596, CK => 
                           net325251, Q => toMemoryPortxADDRINxx31x(0), QN => 
                           n_1061);
   IF_ISAxtoMemoryPort_notify_reg : DFF_X1 port map( D => n7553, CK => 
                           net325226, Q => toMemoryPort_notify_port, QN => 
                           n_1062);
   IF_ISAxtoRegsPort_notify_reg : DFF_X1 port map( D => n3458, CK => clk, Q => 
                           toRegsPort_notify, QN => n7540);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx31x, QN => n_1063);
   IF_ISAxtoRegsPort_regxDSTDATAxx31x : DFF_X1 port map( D => IF_ISAxN10968, CK
                           => net325231, Q => toRegsPortxDSTDATAxx31x, QN => 
                           n_1064);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx31x, QN => n_1065);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx31x, QN => n_1066);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx31x, QN => n_1067);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx31x, QN => n_1068);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx31x, QN => n_1069);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx31x, QN => n_1070);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx31x, QN => n_1071);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx31x, QN => n_1072);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx31x, QN => n_1073);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx31x, QN => n_1074);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx31x, QN => n_1075);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx31x, QN => n_1076);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx31x, QN => n_1077);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx31x, QN => n_1078);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx31x, QN => n_1079);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx31x, QN => n_1080);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx31x, QN => n_1081);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx31x, QN => n_1082);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx31x, QN => n_1083);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx31x, QN => n_1084);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx31x, QN => n_1085);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx31x, QN => n_1086);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx31x, QN => n_1087);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx31x, QN => n_1088);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx31x, QN => n_1089);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx31x, QN => n_1090);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx31x, QN => n_1091);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx31x, QN => n_1092);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx31x, QN => n_1093);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx31x : DFF_X1 port map( D => 
                           IF_RegsxN691, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx31x, QN => n_1094);
   IF_ISAxtoRegsPort_regxDSTDATAxx15x : DFF_X1 port map( D => IF_ISAxN10952, CK
                           => net325231, Q => toRegsPortxDSTDATAxx15x, QN => 
                           n_1095);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx15x, QN => n_1096);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx15x, QN => n_1097);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx15x, QN => n_1098);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx15x, QN => n_1099);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx15x, QN => n_1100);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx15x, QN => n_1101);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx15x, QN => n_1102);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx15x, QN => n_1103);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx15x, QN => n_1104);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx15x, QN => n_1105);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx15x, QN => n_1106);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx15x, QN => n_1107);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx15x, QN => n_1108);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx15x, QN => n_1109);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx15x, QN => n_1110);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx15x, QN => n_1111);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx15x, QN => n_1112);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx15x, QN => n_1113);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx15x, QN => n_1114);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx15x, QN => n_1115);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx15x, QN => n_1116);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx15x, QN => n_1117);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx15x, QN => n_1118);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx15x, QN => n_1119);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx15x, QN => n_1120);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx15x, QN => n_1121);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx15x, QN => n_1122);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx15x, QN => n_1123);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx15x, QN => n_1124);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx15x, QN => n_1125);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx15x : DFF_X1 port map( D => 
                           IF_RegsxN675, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx15x, QN => n_1126);
   IF_ISAxtoRegsPort_regxDSTDATAxx23x : DFF_X1 port map( D => IF_ISAxN10960, CK
                           => net325231, Q => toRegsPortxDSTDATAxx23x, QN => 
                           n_1127);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx23x, QN => n_1128);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx23x, QN => n_1129);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx23x, QN => n_1130);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx23x, QN => n_1131);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx23x, QN => n_1132);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx23x, QN => n_1133);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx23x, QN => n_1134);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx23x, QN => n_1135);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx23x, QN => n_1136);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx23x, QN => n_1137);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx23x, QN => n_1138);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx23x, QN => n_1139);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx23x, QN => n_1140);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx23x, QN => n_1141);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx23x, QN => n_1142);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx23x, QN => n_1143);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx23x, QN => n_1144);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx23x, QN => n_1145);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx23x, QN => n_1146);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx23x, QN => n_1147);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx23x, QN => n_1148);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx23x, QN => n_1149);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx23x, QN => n_1150);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx23x, QN => n_1151);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx23x, QN => n_1152);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx23x, QN => n_1153);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx23x, QN => n_1154);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx23x, QN => n_1155);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx23x, QN => n_1156);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx23x, QN => n_1157);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx23x : DFF_X1 port map( D => 
                           IF_RegsxN683, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx23x, QN => n_1158);
   IF_ISAxtoRegsPort_regxDSTDATAxx27x : DFF_X1 port map( D => IF_ISAxN10964, CK
                           => net325231, Q => toRegsPortxDSTDATAxx27x, QN => 
                           n_1159);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx27x, QN => n_1160);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx27x, QN => n_1161);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx27x, QN => n_1162);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx27x, QN => n_1163);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx27x, QN => n_1164);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx27x, QN => n_1165);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx27x, QN => n_1166);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx27x, QN => n_1167);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx27x, QN => n_1168);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx27x, QN => n_1169);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx27x, QN => n_1170);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx27x, QN => n_1171);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx27x, QN => n_1172);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx27x, QN => n_1173);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx27x, QN => n_1174);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx27x, QN => n_1175);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx27x, QN => n_1176);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx27x, QN => n_1177);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx27x, QN => n_1178);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx27x, QN => n_1179);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx27x, QN => n_1180);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx27x, QN => n_1181);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx27x, QN => n_1182);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx27x, QN => n_1183);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx27x, QN => n_1184);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx27x, QN => n_1185);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx27x, QN => n_1186);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx27x, QN => n_1187);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx27x, QN => n_1188);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx27x, QN => n_1189);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx27x : DFF_X1 port map( D => 
                           IF_RegsxN687, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx27x, QN => n_1190);
   IF_ISAxtoRegsPort_regxDSTDATAxx29x : DFF_X1 port map( D => IF_ISAxN10966, CK
                           => net325231, Q => toRegsPortxDSTDATAxx29x, QN => 
                           n_1191);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx29x, QN => n_1192);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx29x, QN => n_1193);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx29x, QN => n_1194);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx29x, QN => n_1195);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx29x, QN => n_1196);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx29x, QN => n_1197);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx29x, QN => n_1198);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx29x, QN => n_1199);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx29x, QN => n_1200);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx29x, QN => n_1201);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx29x, QN => n_1202);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx29x, QN => n_1203);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx29x, QN => n_1204);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx29x, QN => n_1205);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx29x, QN => n_1206);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx29x, QN => n_1207);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx29x, QN => n_1208);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx29x, QN => n_1209);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx29x, QN => n_1210);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx29x, QN => n_1211);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx29x, QN => n_1212);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx29x, QN => n_1213);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx29x, QN => n_1214);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx29x, QN => n_1215);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx29x, QN => n_1216);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx29x, QN => n_1217);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx29x, QN => n_1218);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx29x, QN => n_1219);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx29x, QN => n_1220);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx29x, QN => n_1221);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx29x : DFF_X1 port map( D => 
                           IF_RegsxN689, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx29x, QN => n_1222);
   IF_ISAxtoRegsPort_regxDSTDATAxx30x : DFF_X1 port map( D => IF_ISAxN10967, CK
                           => net325231, Q => toRegsPortxDSTDATAxx30x, QN => 
                           n_1223);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx30x, QN => n_1224);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx30x, QN => n_1225);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx30x, QN => n_1226);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx30x, QN => n_1227);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx30x, QN => n_1228);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx30x, QN => n_1229);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx30x, QN => n_1230);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx30x, QN => n_1231);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx30x, QN => n_1232);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx30x, QN => n_1233);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx30x, QN => n_1234);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx30x, QN => n_1235);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx30x, QN => n_1236);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx30x, QN => n_1237);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx30x, QN => n_1238);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx30x, QN => n_1239);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx30x, QN => n_1240);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx30x, QN => n_1241);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx30x, QN => n_1242);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx30x, QN => n_1243);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx30x, QN => n_1244);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx30x, QN => n_1245);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx30x, QN => n_1246);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx30x, QN => n_1247);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx30x, QN => n_1248);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx30x, QN => n_1249);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx30x, QN => n_1250);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx30x, QN => n_1251);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx30x, QN => n_1252);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx30x, QN => n_1253);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx30x : DFF_X1 port map( D => 
                           IF_RegsxN690, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx30x, QN => n_1254);
   IF_ISAxtoRegsPort_regxDSTDATAxx0x : DFF_X1 port map( D => IF_ISAxN10936, CK 
                           => net325231, Q => toRegsPortxDSTDATAxx0x, QN => 
                           n_1255);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx0x, QN => n_1256);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx0x, QN => n_1257);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx0x, QN => n_1258);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx0x, QN => n_1259);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx0x, QN => n_1260);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx0x, QN => n_1261);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx0x, QN => n_1262);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx0x, QN => n_1263);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx0x, QN => n_1264);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx0x, QN => n_1265);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx0x, QN => n_1266);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx0x, QN => n_1267);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx0x, QN => n_1268);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx0x, QN => n_1269);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx0x, QN => n_1270);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx0x, QN => n_1271);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx0x, QN => n_1272);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx0x, QN => n_1273);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx0x, QN => n_1274);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx0x, QN => n_1275);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx0x, QN => n_1276);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx0x, QN => n_1277);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx0x, QN => n_1278);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx0x, QN => n_1279);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx0x, QN => n_1280);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx0x, QN => n_1281);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx0x, QN => n_1282);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx0x, QN => n_1283);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx0x, QN => n_1284);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx0x, QN => n_1285);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx0x : DFF_X1 port map( D => 
                           IF_RegsxN660, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx0x, QN => n_1286);
   IF_ISAxtoMemoryPort_regxDATAINxx0x : DFF_X1 port map( D => n7591, CK => 
                           net325246, Q => toMemoryPortxDATAINxx0x(0), QN => 
                           n_1287);
   IF_ISAxtoRegsPort_regxDSTDATAxx16x : DFF_X1 port map( D => IF_ISAxN10953, CK
                           => net325231, Q => toRegsPortxDSTDATAxx16x, QN => 
                           n_1288);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx16x, QN => n_1289);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx16x, QN => n_1290);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx16x, QN => n_1291);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx16x, QN => n_1292);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx16x, QN => n_1293);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx16x, QN => n_1294);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx16x, QN => n_1295);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx16x, QN => n_1296);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx16x, QN => n_1297);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx16x, QN => n_1298);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx16x, QN => n_1299);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx16x, QN => n_1300);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx16x, QN => n_1301);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx16x, QN => n_1302);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx16x, QN => n_1303);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx16x, QN => n_1304);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx16x, QN => n_1305);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx16x, QN => n_1306);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx16x, QN => n_1307);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx16x, QN => n_1308);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx16x, QN => n_1309);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx16x, QN => n_1310);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx16x, QN => n_1311);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx16x, QN => n_1312);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx16x, QN => n_1313);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx16x, QN => n_1314);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx16x, QN => n_1315);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx16x, QN => n_1316);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx16x, QN => n_1317);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx16x, QN => n_1318);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx16x : DFF_X1 port map( D => 
                           IF_RegsxN676, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx16x, QN => n_1319);
   IF_ISAxtoRegsPort_regxDSTDATAxx24x : DFF_X1 port map( D => IF_ISAxN10961, CK
                           => net325231, Q => toRegsPortxDSTDATAxx24x, QN => 
                           n_1320);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx24x, QN => n_1321);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx24x, QN => n_1322);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx24x, QN => n_1323);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx24x, QN => n_1324);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx24x, QN => n_1325);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx24x, QN => n_1326);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx24x, QN => n_1327);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx24x, QN => n_1328);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx24x, QN => n_1329);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx24x, QN => n_1330);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx24x, QN => n_1331);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx24x, QN => n_1332);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx24x, QN => n_1333);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx24x, QN => n_1334);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx24x, QN => n_1335);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx24x, QN => n_1336);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx24x, QN => n_1337);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx24x, QN => n_1338);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx24x, QN => n_1339);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx24x, QN => n_1340);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx24x, QN => n_1341);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx24x, QN => n_1342);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx24x, QN => n_1343);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx24x, QN => n_1344);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx24x, QN => n_1345);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx24x, QN => n_1346);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx24x, QN => n_1347);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx24x, QN => n_1348);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx24x, QN => n_1349);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx24x, QN => n_1350);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx24x : DFF_X1 port map( D => 
                           IF_RegsxN684, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx24x, QN => n_1351);
   IF_ISAxtoRegsPort_regxDSTDATAxx28x : DFF_X1 port map( D => IF_ISAxN10965, CK
                           => net325231, Q => toRegsPortxDSTDATAxx28x, QN => 
                           n_1352);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx28x, QN => n_1353);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx28x, QN => n_1354);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx28x, QN => n_1355);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx28x, QN => n_1356);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx28x, QN => n_1357);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx28x, QN => n_1358);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx28x, QN => n_1359);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx28x, QN => n_1360);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx28x, QN => n_1361);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx28x, QN => n_1362);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx28x, QN => n_1363);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx28x, QN => n_1364);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx28x, QN => n_1365);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx28x, QN => n_1366);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx28x, QN => n_1367);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx28x, QN => n_1368);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx28x, QN => n_1369);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx28x, QN => n_1370);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx28x, QN => n_1371);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx28x, QN => n_1372);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx28x, QN => n_1373);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx28x, QN => n_1374);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx28x, QN => n_1375);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx28x, QN => n_1376);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx28x, QN => n_1377);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx28x, QN => n_1378);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx28x, QN => n_1379);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx28x, QN => n_1380);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx28x, QN => n_1381);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx28x, QN => n_1382);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx28x : DFF_X1 port map( D => 
                           IF_RegsxN688, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx28x, QN => n_1383);
   IF_ISAxtoRegsPort_regxDSTDATAxx10x : DFF_X1 port map( D => IF_ISAxN10947, CK
                           => net325231, Q => toRegsPortxDSTDATAxx10x, QN => 
                           n_1384);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx10x, QN => n_1385);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx10x, QN => n_1386);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx10x, QN => n_1387);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx10x, QN => n_1388);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx10x, QN => n_1389);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx10x, QN => n_1390);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx10x, QN => n_1391);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx10x, QN => n_1392);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx10x, QN => n_1393);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx10x, QN => n_1394);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx10x, QN => n_1395);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx10x, QN => n_1396);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx10x, QN => n_1397);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx10x, QN => n_1398);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx10x, QN => n_1399);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx10x, QN => n_1400);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx10x, QN => n_1401);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx10x, QN => n_1402);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx10x, QN => n_1403);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx10x, QN => n_1404);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx10x, QN => n_1405);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx10x, QN => n_1406);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx10x, QN => n_1407);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx10x, QN => n_1408);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx10x, QN => n_1409);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx10x, QN => n_1410);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx10x, QN => n_1411);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx10x, QN => n_1412);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx10x, QN => n_1413);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx10x, QN => n_1414);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx10x : DFF_X1 port map( D => 
                           IF_RegsxN670, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx10x, QN => n_1415);
   IF_ISAxtoRegsPort_regxDSTDATAxx26x : DFF_X1 port map( D => IF_ISAxN10963, CK
                           => net325231, Q => toRegsPortxDSTDATAxx26x, QN => 
                           n_1416);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx26x, QN => n_1417);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx26x, QN => n_1418);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx26x, QN => n_1419);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx26x, QN => n_1420);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx26x, QN => n_1421);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx26x, QN => n_1422);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx26x, QN => n_1423);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx26x, QN => n_1424);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx26x, QN => n_1425);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx26x, QN => n_1426);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx26x, QN => n_1427);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx26x, QN => n_1428);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx26x, QN => n_1429);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx26x, QN => n_1430);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx26x, QN => n_1431);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx26x, QN => n_1432);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx26x, QN => n_1433);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx26x, QN => n_1434);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx26x, QN => n_1435);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx26x, QN => n_1436);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx26x, QN => n_1437);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx26x, QN => n_1438);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx26x, QN => n_1439);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx26x, QN => n_1440);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx26x, QN => n_1441);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx26x, QN => n_1442);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx26x, QN => n_1443);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx26x, QN => n_1444);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx26x, QN => n_1445);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx26x, QN => n_1446);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx26x : DFF_X1 port map( D => 
                           IF_RegsxN686, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx26x, QN => n_1447);
   IF_ISAxtoRegsPort_regxDSTDATAxx12x : DFF_X1 port map( D => IF_ISAxN10949, CK
                           => net325231, Q => toRegsPortxDSTDATAxx12x, QN => 
                           n_1448);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx12x, QN => n_1449);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx12x, QN => n_1450);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx12x, QN => n_1451);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx12x, QN => n_1452);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx12x, QN => n_1453);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx12x, QN => n_1454);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx12x, QN => n_1455);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx12x, QN => n_1456);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx12x, QN => n_1457);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx12x, QN => n_1458);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx12x, QN => n_1459);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx12x, QN => n_1460);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx12x, QN => n_1461);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx12x, QN => n_1462);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx12x, QN => n_1463);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx12x, QN => n_1464);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx12x, QN => n_1465);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx12x, QN => n_1466);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx12x, QN => n_1467);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx12x, QN => n_1468);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx12x, QN => n_1469);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx12x, QN => n_1470);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx12x, QN => n_1471);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx12x, QN => n_1472);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx12x, QN => n_1473);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx12x, QN => n_1474);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx12x, QN => n_1475);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx12x, QN => n_1476);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx12x, QN => n_1477);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx12x, QN => n_1478);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx12x : DFF_X1 port map( D => 
                           IF_RegsxN672, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx12x, QN => n_1479);
   IF_ISAxtoRegsPort_regxDSTDATAxx20x : DFF_X1 port map( D => IF_ISAxN10957, CK
                           => net325231, Q => toRegsPortxDSTDATAxx20x, QN => 
                           n_1480);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx20x, QN => n_1481);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx20x, QN => n_1482);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx20x, QN => n_1483);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx20x, QN => n_1484);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx20x, QN => n_1485);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx20x, QN => n_1486);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx20x, QN => n_1487);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx20x, QN => n_1488);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx20x, QN => n_1489);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx20x, QN => n_1490);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx20x, QN => n_1491);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx20x, QN => n_1492);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx20x, QN => n_1493);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx20x, QN => n_1494);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx20x, QN => n_1495);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx20x, QN => n_1496);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx20x, QN => n_1497);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx20x, QN => n_1498);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx20x, QN => n_1499);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx20x, QN => n_1500);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx20x, QN => n_1501);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx20x, QN => n_1502);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx20x, QN => n_1503);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx20x, QN => n_1504);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx20x, QN => n_1505);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx20x, QN => n_1506);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx20x, QN => n_1507);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx20x, QN => n_1508);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx20x, QN => n_1509);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx20x, QN => n_1510);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx20x : DFF_X1 port map( D => 
                           IF_RegsxN680, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx20x, QN => n_1511);
   IF_ISAxtoRegsPort_regxDSTDATAxx22x : DFF_X1 port map( D => IF_ISAxN10959, CK
                           => net325231, Q => toRegsPortxDSTDATAxx22x, QN => 
                           n_1512);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx22x, QN => n_1513);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx22x, QN => n_1514);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx22x, QN => n_1515);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx22x, QN => n_1516);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx22x, QN => n_1517);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx22x, QN => n_1518);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx22x, QN => n_1519);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx22x, QN => n_1520);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx22x, QN => n_1521);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx22x, QN => n_1522);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx22x, QN => n_1523);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx22x, QN => n_1524);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx22x, QN => n_1525);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx22x, QN => n_1526);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx22x, QN => n_1527);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx22x, QN => n_1528);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx22x, QN => n_1529);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx22x, QN => n_1530);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx22x, QN => n_1531);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx22x, QN => n_1532);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx22x, QN => n_1533);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx22x, QN => n_1534);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx22x, QN => n_1535);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx22x, QN => n_1536);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx22x, QN => n_1537);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx22x, QN => n_1538);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx22x, QN => n_1539);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx22x, QN => n_1540);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx22x, QN => n_1541);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx22x, QN => n_1542);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx22x : DFF_X1 port map( D => 
                           IF_RegsxN682, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx22x, QN => n_1543);
   IF_ISAxtoRegsPort_regxDSTDATAxx8x : DFF_X1 port map( D => IF_ISAxN10945, CK 
                           => net325231, Q => toRegsPortxDSTDATAxx8x, QN => 
                           n_1544);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx8x, QN => n_1545);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx8x, QN => n_1546);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx8x, QN => n_1547);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx8x, QN => n_1548);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx8x, QN => n_1549);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx8x, QN => n_1550);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx8x, QN => n_1551);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx8x, QN => n_1552);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx8x, QN => n_1553);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx8x, QN => n_1554);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx8x, QN => n_1555);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx8x, QN => n_1556);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx8x, QN => n_1557);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx8x, QN => n_1558);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx8x, QN => n_1559);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx8x, QN => n_1560);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx8x, QN => n_1561);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx8x, QN => n_1562);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx8x, QN => n_1563);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx8x, QN => n_1564);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx8x, QN => n_1565);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx8x, QN => n_1566);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx8x, QN => n_1567);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx8x, QN => n_1568);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx8x, QN => n_1569);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx8x, QN => n_1570);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx8x, QN => n_1571);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx8x, QN => n_1572);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx8x, QN => n_1573);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx8x, QN => n_1574);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx8x : DFF_X1 port map( D => 
                           IF_RegsxN668, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx8x, QN => n_1575);
   IF_ISAxtoRegsPort_regxDSTDATAxx11x : DFF_X1 port map( D => IF_ISAxN10948, CK
                           => net325231, Q => toRegsPortxDSTDATAxx11x, QN => 
                           n_1576);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx11x, QN => n_1577);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx11x, QN => n_1578);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx11x, QN => n_1579);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx11x, QN => n_1580);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx11x, QN => n_1581);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx11x, QN => n_1582);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx11x, QN => n_1583);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx11x, QN => n_1584);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx11x, QN => n_1585);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx11x, QN => n_1586);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx11x, QN => n_1587);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx11x, QN => n_1588);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx11x, QN => n_1589);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx11x, QN => n_1590);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx11x, QN => n_1591);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx11x, QN => n_1592);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx11x, QN => n_1593);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx11x, QN => n_1594);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx11x, QN => n_1595);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx11x, QN => n_1596);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx11x, QN => n_1597);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx11x, QN => n_1598);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx11x, QN => n_1599);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx11x, QN => n_1600);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx11x, QN => n_1601);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx11x, QN => n_1602);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx11x, QN => n_1603);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx11x, QN => n_1604);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx11x, QN => n_1605);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx11x, QN => n_1606);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx11x : DFF_X1 port map( D => 
                           IF_RegsxN671, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx11x, QN => n_1607);
   IF_ISAxtoRegsPort_regxDSTDATAxx13x : DFF_X1 port map( D => IF_ISAxN10950, CK
                           => net325231, Q => toRegsPortxDSTDATAxx13x, QN => 
                           n_1608);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx13x, QN => n_1609);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx13x, QN => n_1610);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx13x, QN => n_1611);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx13x, QN => n_1612);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx13x, QN => n_1613);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx13x, QN => n_1614);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx13x, QN => n_1615);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx13x, QN => n_1616);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx13x, QN => n_1617);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx13x, QN => n_1618);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx13x, QN => n_1619);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx13x, QN => n_1620);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx13x, QN => n_1621);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx13x, QN => n_1622);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx13x, QN => n_1623);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx13x, QN => n_1624);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx13x, QN => n_1625);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx13x, QN => n_1626);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx13x, QN => n_1627);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx13x, QN => n_1628);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx13x, QN => n_1629);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx13x, QN => n_1630);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx13x, QN => n_1631);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx13x, QN => n_1632);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx13x, QN => n_1633);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx13x, QN => n_1634);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx13x, QN => n_1635);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx13x, QN => n_1636);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx13x, QN => n_1637);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx13x, QN => n_1638);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx13x : DFF_X1 port map( D => 
                           IF_RegsxN673, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx13x, QN => n_1639);
   IF_ISAxtoRegsPort_regxDSTDATAxx14x : DFF_X1 port map( D => IF_ISAxN10951, CK
                           => net325231, Q => toRegsPortxDSTDATAxx14x, QN => 
                           n_1640);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx14x, QN => n_1641);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx14x, QN => n_1642);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx14x, QN => n_1643);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx14x, QN => n_1644);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx14x, QN => n_1645);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx14x, QN => n_1646);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx14x, QN => n_1647);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx14x, QN => n_1648);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx14x, QN => n_1649);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx14x, QN => n_1650);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx14x, QN => n_1651);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx14x, QN => n_1652);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx14x, QN => n_1653);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx14x, QN => n_1654);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx14x, QN => n_1655);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx14x, QN => n_1656);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx14x, QN => n_1657);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx14x, QN => n_1658);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx14x, QN => n_1659);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx14x, QN => n_1660);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx14x, QN => n_1661);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx14x, QN => n_1662);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx14x, QN => n_1663);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx14x, QN => n_1664);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx14x, QN => n_1665);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx14x, QN => n_1666);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx14x, QN => n_1667);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx14x, QN => n_1668);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx14x, QN => n_1669);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx14x, QN => n_1670);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx14x : DFF_X1 port map( D => 
                           IF_RegsxN674, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx14x, QN => n_1671);
   IF_ISAxtoRegsPort_regxDSTDATAxx4x : DFF_X1 port map( D => IF_ISAxN10941, CK 
                           => net325231, Q => toRegsPortxDSTDATAxx4x, QN => 
                           n_1672);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx4x, QN => n_1673);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx4x, QN => n_1674);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx4x, QN => n_1675);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx4x, QN => n_1676);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx4x, QN => n_1677);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx4x, QN => n_1678);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx4x, QN => n_1679);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx4x, QN => n_1680);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx4x, QN => n_1681);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx4x, QN => n_1682);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx4x, QN => n_1683);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx4x, QN => n_1684);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx4x, QN => n_1685);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx4x, QN => n_1686);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx4x, QN => n_1687);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx4x, QN => n_1688);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx4x, QN => n_1689);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx4x, QN => n_1690);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx4x, QN => n_1691);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx4x, QN => n_1692);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx4x, QN => n_1693);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx4x, QN => n_1694);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx4x, QN => n_1695);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx4x, QN => n_1696);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx4x, QN => n_1697);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx4x, QN => n_1698);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx4x, QN => n_1699);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx4x, QN => n_1700);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx4x, QN => n_1701);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx4x, QN => n_1702);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx4x : DFF_X1 port map( D => 
                           IF_RegsxN664, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx4x, QN => n_1703);
   IF_ISAxtoMemoryPort_regxDATAINxx4x : DFF_X1 port map( D => n7590, CK => 
                           net325246, Q => toMemoryPortxDATAINxx4x(0), QN => 
                           n_1704);
   IF_ISAxtoRegsPort_regxDSTDATAxx17x : DFF_X1 port map( D => IF_ISAxN10954, CK
                           => net325231, Q => toRegsPortxDSTDATAxx17x, QN => 
                           n_1705);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx17x, QN => n_1706);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx17x, QN => n_1707);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx17x, QN => n_1708);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx17x, QN => n_1709);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx17x, QN => n_1710);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx17x, QN => n_1711);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx17x, QN => n_1712);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx17x, QN => n_1713);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx17x, QN => n_1714);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx17x, QN => n_1715);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx17x, QN => n_1716);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx17x, QN => n_1717);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx17x, QN => n_1718);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx17x, QN => n_1719);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx17x, QN => n_1720);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx17x, QN => n_1721);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx17x, QN => n_1722);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx17x, QN => n_1723);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx17x, QN => n_1724);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx17x, QN => n_1725);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx17x, QN => n_1726);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx17x, QN => n_1727);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx17x, QN => n_1728);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx17x, QN => n_1729);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx17x, QN => n_1730);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx17x, QN => n_1731);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx17x, QN => n_1732);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx17x, QN => n_1733);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx17x, QN => n_1734);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx17x, QN => n_1735);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx17x : DFF_X1 port map( D => 
                           IF_RegsxN677, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx17x, QN => n_1736);
   IF_ISAxtoRegsPort_regxDSTDATAxx25x : DFF_X1 port map( D => IF_ISAxN10962, CK
                           => net325231, Q => toRegsPortxDSTDATAxx25x, QN => 
                           n_1737);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx25x, QN => n_1738);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx25x, QN => n_1739);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx25x, QN => n_1740);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx25x, QN => n_1741);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx25x, QN => n_1742);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx25x, QN => n_1743);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx25x, QN => n_1744);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx25x, QN => n_1745);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx25x, QN => n_1746);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx25x, QN => n_1747);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx25x, QN => n_1748);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx25x, QN => n_1749);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx25x, QN => n_1750);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx25x, QN => n_1751);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx25x, QN => n_1752);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx25x, QN => n_1753);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx25x, QN => n_1754);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx25x, QN => n_1755);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx25x, QN => n_1756);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx25x, QN => n_1757);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx25x, QN => n_1758);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx25x, QN => n_1759);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx25x, QN => n_1760);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx25x, QN => n_1761);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx25x, QN => n_1762);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx25x, QN => n_1763);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx25x, QN => n_1764);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx25x, QN => n_1765);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx25x, QN => n_1766);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx25x, QN => n_1767);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx25x : DFF_X1 port map( D => 
                           IF_RegsxN685, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx25x, QN => n_1768);
   IF_ISAxtoRegsPort_regxDSTDATAxx18x : DFF_X1 port map( D => IF_ISAxN10955, CK
                           => net325231, Q => toRegsPortxDSTDATAxx18x, QN => 
                           n_1769);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx18x, QN => n_1770);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx18x, QN => n_1771);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx18x, QN => n_1772);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx18x, QN => n_1773);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx18x, QN => n_1774);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx18x, QN => n_1775);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx18x, QN => n_1776);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx18x, QN => n_1777);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx18x, QN => n_1778);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx18x, QN => n_1779);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx18x, QN => n_1780);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx18x, QN => n_1781);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx18x, QN => n_1782);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx18x, QN => n_1783);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx18x, QN => n_1784);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx18x, QN => n_1785);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx18x, QN => n_1786);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx18x, QN => n_1787);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx18x, QN => n_1788);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx18x, QN => n_1789);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx18x, QN => n_1790);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx18x, QN => n_1791);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx18x, QN => n_1792);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx18x, QN => n_1793);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx18x, QN => n_1794);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx18x, QN => n_1795);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx18x, QN => n_1796);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx18x, QN => n_1797);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx18x, QN => n_1798);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx18x, QN => n_1799);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx18x : DFF_X1 port map( D => 
                           IF_RegsxN678, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx18x, QN => n_1800);
   IF_ISAxtoRegsPort_regxDSTDATAxx19x : DFF_X1 port map( D => IF_ISAxN10956, CK
                           => net325231, Q => toRegsPortxDSTDATAxx19x, QN => 
                           n_1801);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx19x, QN => n_1802);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx19x, QN => n_1803);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx19x, QN => n_1804);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx19x, QN => n_1805);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx19x, QN => n_1806);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx19x, QN => n_1807);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx19x, QN => n_1808);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx19x, QN => n_1809);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx19x, QN => n_1810);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx19x, QN => n_1811);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx19x, QN => n_1812);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx19x, QN => n_1813);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx19x, QN => n_1814);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx19x, QN => n_1815);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx19x, QN => n_1816);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx19x, QN => n_1817);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx19x, QN => n_1818);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx19x, QN => n_1819);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx19x, QN => n_1820);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx19x, QN => n_1821);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx19x, QN => n_1822);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx19x, QN => n_1823);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx19x, QN => n_1824);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx19x, QN => n_1825);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx19x, QN => n_1826);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx19x, QN => n_1827);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx19x, QN => n_1828);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx19x, QN => n_1829);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx19x, QN => n_1830);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx19x, QN => n_1831);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx19x : DFF_X1 port map( D => 
                           IF_RegsxN679, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx19x, QN => n_1832);
   IF_ISAxtoRegsPort_regxDSTDATAxx6x : DFF_X1 port map( D => IF_ISAxN10943, CK 
                           => net325231, Q => toRegsPortxDSTDATAxx6x, QN => 
                           n_1833);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx6x, QN => n_1834);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx6x, QN => n_1835);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx6x, QN => n_1836);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx6x, QN => n_1837);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx6x, QN => n_1838);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx6x, QN => n_1839);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx6x, QN => n_1840);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx6x, QN => n_1841);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx6x, QN => n_1842);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx6x, QN => n_1843);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx6x, QN => n_1844);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx6x, QN => n_1845);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx6x, QN => n_1846);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx6x, QN => n_1847);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx6x, QN => n_1848);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx6x, QN => n_1849);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx6x, QN => n_1850);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx6x, QN => n_1851);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx6x, QN => n_1852);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx6x, QN => n_1853);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx6x, QN => n_1854);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx6x, QN => n_1855);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx6x, QN => n_1856);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx6x, QN => n_1857);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx6x, QN => n_1858);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx6x, QN => n_1859);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx6x, QN => n_1860);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx6x, QN => n_1861);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx6x, QN => n_1862);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx6x, QN => n_1863);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx6x : DFF_X1 port map( D => 
                           IF_RegsxN666, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx6x, QN => n_1864);
   IF_ISAxtoRegsPort_regxDSTDATAxx7x : DFF_X1 port map( D => IF_ISAxN10944, CK 
                           => net325231, Q => toRegsPortxDSTDATAxx7x, QN => 
                           n_1865);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx7x, QN => n_1866);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx7x, QN => n_1867);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx7x, QN => n_1868);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx7x, QN => n_1869);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx7x, QN => n_1870);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx7x, QN => n_1871);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx7x, QN => n_1872);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx7x, QN => n_1873);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx7x, QN => n_1874);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx7x, QN => n_1875);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx7x, QN => n_1876);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx7x, QN => n_1877);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx7x, QN => n_1878);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx7x, QN => n_1879);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx7x, QN => n_1880);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx7x, QN => n_1881);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx7x, QN => n_1882);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx7x, QN => n_1883);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx7x, QN => n_1884);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx7x, QN => n_1885);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx7x, QN => n_1886);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx7x, QN => n_1887);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx7x, QN => n_1888);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx7x, QN => n_1889);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx7x, QN => n_1890);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx7x, QN => n_1891);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx7x, QN => n_1892);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx7x, QN => n_1893);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx7x, QN => n_1894);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx7x, QN => n_1895);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx7x : DFF_X1 port map( D => 
                           IF_RegsxN667, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx7x, QN => n_1896);
   IF_ISAxtoRegsPort_regxDSTDATAxx2x : DFF_X1 port map( D => IF_ISAxN10939, CK 
                           => net325231, Q => toRegsPortxDSTDATAxx2x, QN => 
                           n_1897);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx2x, QN => n_1898);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx2x, QN => n_1899);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx2x, QN => n_1900);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx2x, QN => n_1901);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx2x, QN => n_1902);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx2x, QN => n_1903);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx2x, QN => n_1904);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx2x, QN => n_1905);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx2x, QN => n_1906);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx2x, QN => n_1907);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx2x, QN => n_1908);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx2x, QN => n_1909);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx2x, QN => n_1910);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx2x, QN => n_1911);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx2x, QN => n_1912);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx2x, QN => n_1913);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx2x, QN => n_1914);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx2x, QN => n_1915);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx2x, QN => n_1916);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx2x, QN => n_1917);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx2x, QN => n_1918);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx2x, QN => n_1919);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx2x, QN => n_1920);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx2x, QN => n_1921);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx2x, QN => n_1922);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx2x, QN => n_1923);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx2x, QN => n_1924);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx2x, QN => n_1925);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx2x, QN => n_1926);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx2x, QN => n_1927);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx2x : DFF_X1 port map( D => 
                           IF_RegsxN662, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx2x, QN => n_1928);
   IF_ISAxtoMemoryPort_regxDATAINxx2x : DFF_X1 port map( D => n7589, CK => 
                           net325246, Q => toMemoryPortxDATAINxx2x(0), QN => 
                           n_1929);
   IF_ISAxtoRegsPort_regxDSTDATAxx3x : DFF_X1 port map( D => IF_ISAxN10940, CK 
                           => net325231, Q => toRegsPortxDSTDATAxx3x, QN => 
                           n_1930);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx3x, QN => n_1931);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx3x, QN => n_1932);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx3x, QN => n_1933);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx3x, QN => n_1934);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx3x, QN => n_1935);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx3x, QN => n_1936);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx3x, QN => n_1937);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx3x, QN => n_1938);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx3x, QN => n_1939);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx3x, QN => n_1940);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx3x, QN => n_1941);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx3x, QN => n_1942);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx3x, QN => n_1943);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx3x, QN => n_1944);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx3x, QN => n_1945);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx3x, QN => n_1946);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx3x, QN => n_1947);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx3x, QN => n_1948);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx3x, QN => n_1949);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx3x, QN => n_1950);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx3x, QN => n_1951);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx3x, QN => n_1952);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx3x, QN => n_1953);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx3x, QN => n_1954);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx3x, QN => n_1955);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx3x, QN => n_1956);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx3x, QN => n_1957);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx3x, QN => n_1958);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx3x, QN => n_1959);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx3x, QN => n_1960);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx3x : DFF_X1 port map( D => 
                           IF_RegsxN663, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx3x, QN => n_1961);
   IF_ISAxtoMemoryPort_regxDATAINxx3x : DFF_X1 port map( D => n7588, CK => 
                           net325246, Q => toMemoryPortxDATAINxx3x(0), QN => 
                           n_1962);
   IF_ISAxtoRegsPort_regxDSTDATAxx21x : DFF_X1 port map( D => IF_ISAxN10958, CK
                           => net325231, Q => toRegsPortxDSTDATAxx21x, QN => 
                           n_1963);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx21x, QN => n_1964);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx21x, QN => n_1965);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx21x, QN => n_1966);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx21x, QN => n_1967);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx21x, QN => n_1968);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx21x, QN => n_1969);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx21x, QN => n_1970);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx21x, QN => n_1971);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx21x, QN => n_1972);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx21x, QN => n_1973);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx21x, QN => n_1974);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx21x, QN => n_1975);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx21x, QN => n_1976);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx21x, QN => n_1977);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx21x, QN => n_1978);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx21x, QN => n_1979);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx21x, QN => n_1980);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx21x, QN => n_1981);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx21x, QN => n_1982);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx21x, QN => n_1983);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx21x, QN => n_1984);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx21x, QN => n_1985);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx21x, QN => n_1986);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx21x, QN => n_1987);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx21x, QN => n_1988);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx21x, QN => n_1989);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx21x, QN => n_1990);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx21x, QN => n_1991);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx21x, QN => n_1992);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx21x, QN => n_1993);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx21x : DFF_X1 port map( D => 
                           IF_RegsxN681, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx21x, QN => n_1994);
   IF_ISAxtoRegsPort_regxDSTDATAxx5x : DFF_X1 port map( D => IF_ISAxN10942, CK 
                           => net325231, Q => toRegsPortxDSTDATAxx5x, QN => 
                           n_1995);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx5x, QN => n_1996);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx5x, QN => n_1997);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx5x, QN => n_1998);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx5x, QN => n_1999);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx5x, QN => n_2000);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx5x, QN => n_2001);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx5x, QN => n_2002);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx5x, QN => n_2003);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx5x, QN => n_2004);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx5x, QN => n_2005);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx5x, QN => n_2006);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx5x, QN => n_2007);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx5x, QN => n_2008);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx5x, QN => n_2009);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx5x, QN => n_2010);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx5x, QN => n_2011);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx5x, QN => n_2012);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx5x, QN => n_2013);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx5x, QN => n_2014);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx5x, QN => n_2015);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx5x, QN => n_2016);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx5x, QN => n_2017);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx5x, QN => n_2018);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx5x, QN => n_2019);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx5x, QN => n_2020);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx5x, QN => n_2021);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx5x, QN => n_2022);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx5x, QN => n_2023);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx5x, QN => n_2024);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx5x, QN => n_2025);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx5x : DFF_X1 port map( D => 
                           IF_RegsxN665, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx5x, QN => n_2026);
   IF_ISAxtoRegsPort_regxDSTDATAxx9x : DFF_X1 port map( D => IF_ISAxN10946, CK 
                           => net325231, Q => toRegsPortxDSTDATAxx9x, QN => 
                           n_2027);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx9x, QN => n_2028);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx9x, QN => n_2029);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx9x, QN => n_2030);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx9x, QN => n_2031);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx9x, QN => n_2032);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx9x, QN => n_2033);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx9x, QN => n_2034);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx9x, QN => n_2035);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx9x, QN => n_2036);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx9x, QN => n_2037);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx9x, QN => n_2038);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx9x, QN => n_2039);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx9x, QN => n_2040);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx9x, QN => n_2041);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx9x, QN => n_2042);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx9x, QN => n_2043);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx9x, QN => n_2044);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx9x, QN => n_2045);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx9x, QN => n_2046);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx9x, QN => n_2047);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx9x, QN => n_2048);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx9x, QN => n_2049);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx9x, QN => n_2050);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx9x, QN => n_2051);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx9x, QN => n_2052);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx9x, QN => n_2053);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx9x, QN => n_2054);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx9x, QN => n_2055);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx9x, QN => n_2056);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx9x, QN => n_2057);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx9x : DFF_X1 port map( D => 
                           IF_RegsxN669, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx9x, QN => n_2058);
   IF_ISAxtoRegsPort_regxDSTDATAxx1x : DFF_X1 port map( D => IF_ISAxN10938, CK 
                           => net325231, Q => toRegsPortxDSTDATAxx1x, QN => 
                           n_2059);
   IF_RegsxRegsToCtl_port_regxREG_FILE_31xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325256, Q => 
                           fromRegsPortxREG_FILE_31xx1x, QN => n_2060);
   IF_RegsxRegsToCtl_port_regxREG_FILE_01xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325406, Q => 
                           fromRegsPortxREG_FILE_01xx1x, QN => n_2061);
   IF_RegsxRegsToCtl_port_regxREG_FILE_02xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325401, Q => 
                           fromRegsPortxREG_FILE_02xx1x, QN => n_2062);
   IF_RegsxRegsToCtl_port_regxREG_FILE_03xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325396, Q => 
                           fromRegsPortxREG_FILE_03xx1x, QN => n_2063);
   IF_RegsxRegsToCtl_port_regxREG_FILE_04xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325391, Q => 
                           fromRegsPortxREG_FILE_04xx1x, QN => n_2064);
   IF_RegsxRegsToCtl_port_regxREG_FILE_05xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325386, Q => 
                           fromRegsPortxREG_FILE_05xx1x, QN => n_2065);
   IF_RegsxRegsToCtl_port_regxREG_FILE_06xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325381, Q => 
                           fromRegsPortxREG_FILE_06xx1x, QN => n_2066);
   IF_RegsxRegsToCtl_port_regxREG_FILE_07xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325376, Q => 
                           fromRegsPortxREG_FILE_07xx1x, QN => n_2067);
   IF_RegsxRegsToCtl_port_regxREG_FILE_08xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325371, Q => 
                           fromRegsPortxREG_FILE_08xx1x, QN => n_2068);
   IF_RegsxRegsToCtl_port_regxREG_FILE_09xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325366, Q => 
                           fromRegsPortxREG_FILE_09xx1x, QN => n_2069);
   IF_RegsxRegsToCtl_port_regxREG_FILE_10xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325361, Q => 
                           fromRegsPortxREG_FILE_10xx1x, QN => n_2070);
   IF_RegsxRegsToCtl_port_regxREG_FILE_11xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325356, Q => 
                           fromRegsPortxREG_FILE_11xx1x, QN => n_2071);
   IF_RegsxRegsToCtl_port_regxREG_FILE_12xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325351, Q => 
                           fromRegsPortxREG_FILE_12xx1x, QN => n_2072);
   IF_RegsxRegsToCtl_port_regxREG_FILE_13xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325346, Q => 
                           fromRegsPortxREG_FILE_13xx1x, QN => n_2073);
   IF_RegsxRegsToCtl_port_regxREG_FILE_14xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325341, Q => 
                           fromRegsPortxREG_FILE_14xx1x, QN => n_2074);
   IF_RegsxRegsToCtl_port_regxREG_FILE_15xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325336, Q => 
                           fromRegsPortxREG_FILE_15xx1x, QN => n_2075);
   IF_RegsxRegsToCtl_port_regxREG_FILE_16xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325331, Q => 
                           fromRegsPortxREG_FILE_16xx1x, QN => n_2076);
   IF_RegsxRegsToCtl_port_regxREG_FILE_17xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325326, Q => 
                           fromRegsPortxREG_FILE_17xx1x, QN => n_2077);
   IF_RegsxRegsToCtl_port_regxREG_FILE_18xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325321, Q => 
                           fromRegsPortxREG_FILE_18xx1x, QN => n_2078);
   IF_RegsxRegsToCtl_port_regxREG_FILE_19xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325316, Q => 
                           fromRegsPortxREG_FILE_19xx1x, QN => n_2079);
   IF_RegsxRegsToCtl_port_regxREG_FILE_20xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325311, Q => 
                           fromRegsPortxREG_FILE_20xx1x, QN => n_2080);
   IF_RegsxRegsToCtl_port_regxREG_FILE_21xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325306, Q => 
                           fromRegsPortxREG_FILE_21xx1x, QN => n_2081);
   IF_RegsxRegsToCtl_port_regxREG_FILE_22xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325301, Q => 
                           fromRegsPortxREG_FILE_22xx1x, QN => n_2082);
   IF_RegsxRegsToCtl_port_regxREG_FILE_23xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325296, Q => 
                           fromRegsPortxREG_FILE_23xx1x, QN => n_2083);
   IF_RegsxRegsToCtl_port_regxREG_FILE_24xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325291, Q => 
                           fromRegsPortxREG_FILE_24xx1x, QN => n_2084);
   IF_RegsxRegsToCtl_port_regxREG_FILE_25xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325286, Q => 
                           fromRegsPortxREG_FILE_25xx1x, QN => n_2085);
   IF_RegsxRegsToCtl_port_regxREG_FILE_26xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325281, Q => 
                           fromRegsPortxREG_FILE_26xx1x, QN => n_2086);
   IF_RegsxRegsToCtl_port_regxREG_FILE_27xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325276, Q => 
                           fromRegsPortxREG_FILE_27xx1x, QN => n_2087);
   IF_RegsxRegsToCtl_port_regxREG_FILE_28xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325271, Q => 
                           fromRegsPortxREG_FILE_28xx1x, QN => n_2088);
   IF_RegsxRegsToCtl_port_regxREG_FILE_29xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325266, Q => 
                           fromRegsPortxREG_FILE_29xx1x, QN => n_2089);
   IF_RegsxRegsToCtl_port_regxREG_FILE_30xx1x : DFF_X1 port map( D => 
                           IF_RegsxN661, CK => net325261, Q => 
                           fromRegsPortxREG_FILE_30xx1x, QN => n_2090);
   IF_ISAxtoMemoryPort_regxDATAINxx1x : DFF_X1 port map( D => n7587, CK => 
                           net325246, Q => toMemoryPortxDATAINxx1x(0), QN => 
                           n_2091);
   IF_ISAxtoMemoryPort_regxDATAINxx9x : DFF_X1 port map( D => IF_ISAxN10846, CK
                           => net325246, Q => toMemoryPortxDATAINxx9x(0), QN =>
                           n_2092);
   IF_ISAxtoMemoryPort_regxDATAINxx5x : DFF_X1 port map( D => IF_ISAxN10842, CK
                           => net325246, Q => toMemoryPortxDATAINxx5x(0), QN =>
                           n_2093);
   IF_ISAxtoMemoryPort_regxDATAINxx21x : DFF_X1 port map( D => IF_ISAxN10858, 
                           CK => net325246, Q => toMemoryPortxDATAINxx21x(0), 
                           QN => n_2094);
   IF_ISAxtoMemoryPort_regxDATAINxx7x : DFF_X1 port map( D => IF_ISAxN10844, CK
                           => net325246, Q => toMemoryPortxDATAINxx7x(0), QN =>
                           n_2095);
   IF_ISAxtoMemoryPort_regxDATAINxx6x : DFF_X1 port map( D => IF_ISAxN10843, CK
                           => net325246, Q => toMemoryPortxDATAINxx6x(0), QN =>
                           n_2096);
   IF_ISAxtoMemoryPort_regxDATAINxx19x : DFF_X1 port map( D => IF_ISAxN10856, 
                           CK => net325246, Q => toMemoryPortxDATAINxx19x(0), 
                           QN => n_2097);
   IF_ISAxtoMemoryPort_regxDATAINxx18x : DFF_X1 port map( D => IF_ISAxN10855, 
                           CK => net325246, Q => toMemoryPortxDATAINxx18x(0), 
                           QN => n_2098);
   IF_ISAxtoMemoryPort_regxDATAINxx25x : DFF_X1 port map( D => IF_ISAxN10862, 
                           CK => net325246, Q => toMemoryPortxDATAINxx25x(0), 
                           QN => n_2099);
   IF_ISAxtoMemoryPort_regxDATAINxx17x : DFF_X1 port map( D => IF_ISAxN10854, 
                           CK => net325246, Q => toMemoryPortxDATAINxx17x(0), 
                           QN => n_2100);
   IF_ISAxtoMemoryPort_regxDATAINxx14x : DFF_X1 port map( D => IF_ISAxN10851, 
                           CK => net325246, Q => toMemoryPortxDATAINxx14x(0), 
                           QN => n_2101);
   IF_ISAxtoMemoryPort_regxDATAINxx13x : DFF_X1 port map( D => IF_ISAxN10850, 
                           CK => net325246, Q => toMemoryPortxDATAINxx13x(0), 
                           QN => n_2102);
   IF_ISAxtoMemoryPort_regxDATAINxx11x : DFF_X1 port map( D => IF_ISAxN10848, 
                           CK => net325246, Q => toMemoryPortxDATAINxx11x(0), 
                           QN => n_2103);
   IF_ISAxtoMemoryPort_regxDATAINxx8x : DFF_X1 port map( D => IF_ISAxN10845, CK
                           => net325246, Q => toMemoryPortxDATAINxx8x(0), QN =>
                           n_2104);
   IF_ISAxtoMemoryPort_regxDATAINxx22x : DFF_X1 port map( D => IF_ISAxN10859, 
                           CK => net325246, Q => toMemoryPortxDATAINxx22x(0), 
                           QN => n_2105);
   IF_ISAxtoMemoryPort_regxDATAINxx20x : DFF_X1 port map( D => IF_ISAxN10857, 
                           CK => net325246, Q => toMemoryPortxDATAINxx20x(0), 
                           QN => n_2106);
   IF_ISAxtoMemoryPort_regxDATAINxx12x : DFF_X1 port map( D => IF_ISAxN10849, 
                           CK => net325246, Q => toMemoryPortxDATAINxx12x(0), 
                           QN => n_2107);
   IF_ISAxtoMemoryPort_regxDATAINxx26x : DFF_X1 port map( D => IF_ISAxN10863, 
                           CK => net325246, Q => toMemoryPortxDATAINxx26x(0), 
                           QN => n_2108);
   IF_ISAxtoMemoryPort_regxDATAINxx10x : DFF_X1 port map( D => IF_ISAxN10847, 
                           CK => net325246, Q => toMemoryPortxDATAINxx10x(0), 
                           QN => n_2109);
   IF_ISAxtoMemoryPort_regxDATAINxx28x : DFF_X1 port map( D => IF_ISAxN10865, 
                           CK => net325246, Q => toMemoryPortxDATAINxx28x(0), 
                           QN => n_2110);
   IF_ISAxtoMemoryPort_regxDATAINxx24x : DFF_X1 port map( D => IF_ISAxN10861, 
                           CK => net325246, Q => toMemoryPortxDATAINxx24x(0), 
                           QN => n_2111);
   IF_ISAxtoMemoryPort_regxDATAINxx16x : DFF_X1 port map( D => IF_ISAxN10853, 
                           CK => net325246, Q => toMemoryPortxDATAINxx16x(0), 
                           QN => n_2112);
   IF_ISAxtoMemoryPort_regxDATAINxx30x : DFF_X1 port map( D => IF_ISAxN10867, 
                           CK => net325246, Q => toMemoryPortxDATAINxx30x(0), 
                           QN => n_2113);
   IF_ISAxtoMemoryPort_regxDATAINxx29x : DFF_X1 port map( D => IF_ISAxN10866, 
                           CK => net325246, Q => toMemoryPortxDATAINxx29x(0), 
                           QN => n_2114);
   IF_ISAxtoMemoryPort_regxDATAINxx27x : DFF_X1 port map( D => IF_ISAxN10864, 
                           CK => net325246, Q => toMemoryPortxDATAINxx27x(0), 
                           QN => n_2115);
   IF_ISAxtoMemoryPort_regxDATAINxx23x : DFF_X1 port map( D => IF_ISAxN10860, 
                           CK => net325246, Q => toMemoryPortxDATAINxx23x(0), 
                           QN => n_2116);
   IF_ISAxtoMemoryPort_regxDATAINxx15x : DFF_X1 port map( D => IF_ISAxN10852, 
                           CK => net325246, Q => toMemoryPortxDATAINxx15x(0), 
                           QN => n_2117);
   IF_ISAxtoMemoryPort_regxDATAINxx31x : DFF_X1 port map( D => IF_ISAxN10868, 
                           CK => net325246, Q => toMemoryPortxDATAINxx31x(0), 
                           QN => n_2118);
   DP_OP_679J14_122_3096xU33 : FA_X1 port map( A => ashr_25xAx0x, B => n7551, 
                           CI => DP_OP_679J14_122_3096xn68, CO => 
                           DP_OP_679J14_122_3096xn32, S => 
                           DP_OP_679J14_122_3096xn69);
   DP_OP_679J14_122_3096xU32 : FA_X1 port map( A => DP_OP_679J14_122_3096xn67, 
                           B => ashr_25xAx1x, CI => DP_OP_679J14_122_3096xn32, 
                           CO => DP_OP_679J14_122_3096xn31, S => 
                           DP_OP_679J14_122_3096xn70);
   DP_OP_679J14_122_3096xU31 : FA_X1 port map( A => DP_OP_679J14_122_3096xn66, 
                           B => ashr_25xAx2x, CI => DP_OP_679J14_122_3096xn31, 
                           CO => DP_OP_679J14_122_3096xn30, S => 
                           DP_OP_679J14_122_3096xn71);
   DP_OP_679J14_122_3096xU30 : FA_X1 port map( A => DP_OP_679J14_122_3096xn65, 
                           B => ashr_25xAx3x, CI => DP_OP_679J14_122_3096xn30, 
                           CO => DP_OP_679J14_122_3096xn29, S => 
                           DP_OP_679J14_122_3096xn72);
   DP_OP_679J14_122_3096xU29 : FA_X1 port map( A => DP_OP_679J14_122_3096xn64, 
                           B => ashr_25xAx4x, CI => DP_OP_679J14_122_3096xn29, 
                           CO => DP_OP_679J14_122_3096xn28, S => 
                           DP_OP_679J14_122_3096xn73);
   DP_OP_679J14_122_3096xU28 : FA_X1 port map( A => DP_OP_679J14_122_3096xn63, 
                           B => ashr_25xAx5x, CI => DP_OP_679J14_122_3096xn28, 
                           CO => DP_OP_679J14_122_3096xn27, S => 
                           DP_OP_679J14_122_3096xn74);
   DP_OP_679J14_122_3096xU27 : FA_X1 port map( A => DP_OP_679J14_122_3096xn62, 
                           B => ashr_25xAx6x, CI => DP_OP_679J14_122_3096xn27, 
                           CO => DP_OP_679J14_122_3096xn26, S => 
                           DP_OP_679J14_122_3096xn75);
   DP_OP_679J14_122_3096xU26 : FA_X1 port map( A => DP_OP_679J14_122_3096xn61, 
                           B => ashr_25xAx7x, CI => DP_OP_679J14_122_3096xn26, 
                           CO => DP_OP_679J14_122_3096xn25, S => 
                           DP_OP_679J14_122_3096xn76);
   DP_OP_679J14_122_3096xU25 : FA_X1 port map( A => DP_OP_679J14_122_3096xn60, 
                           B => ashr_25xAx8x, CI => DP_OP_679J14_122_3096xn25, 
                           CO => DP_OP_679J14_122_3096xn24, S => 
                           DP_OP_679J14_122_3096xn77);
   DP_OP_679J14_122_3096xU24 : FA_X1 port map( A => DP_OP_679J14_122_3096xn59, 
                           B => ashr_25xAx9x, CI => DP_OP_679J14_122_3096xn24, 
                           CO => DP_OP_679J14_122_3096xn23, S => 
                           DP_OP_679J14_122_3096xn78);
   DP_OP_679J14_122_3096xU23 : FA_X1 port map( A => DP_OP_679J14_122_3096xn58, 
                           B => ashr_25xAx10x, CI => DP_OP_679J14_122_3096xn23,
                           CO => DP_OP_679J14_122_3096xn22, S => 
                           DP_OP_679J14_122_3096xn79);
   DP_OP_679J14_122_3096xU22 : FA_X1 port map( A => DP_OP_679J14_122_3096xn57, 
                           B => ashr_25xAx11x, CI => DP_OP_679J14_122_3096xn22,
                           CO => DP_OP_679J14_122_3096xn21, S => 
                           DP_OP_679J14_122_3096xn80);
   DP_OP_679J14_122_3096xU21 : FA_X1 port map( A => DP_OP_679J14_122_3096xn56, 
                           B => ashr_25xAx12x, CI => DP_OP_679J14_122_3096xn21,
                           CO => DP_OP_679J14_122_3096xn20, S => 
                           DP_OP_679J14_122_3096xn81);
   DP_OP_679J14_122_3096xU20 : FA_X1 port map( A => DP_OP_679J14_122_3096xn55, 
                           B => ashr_25xAx13x, CI => DP_OP_679J14_122_3096xn20,
                           CO => DP_OP_679J14_122_3096xn19, S => 
                           DP_OP_679J14_122_3096xn82);
   DP_OP_679J14_122_3096xU19 : FA_X1 port map( A => DP_OP_679J14_122_3096xn54, 
                           B => ashr_25xAx14x, CI => DP_OP_679J14_122_3096xn19,
                           CO => DP_OP_679J14_122_3096xn18, S => 
                           DP_OP_679J14_122_3096xn83);
   DP_OP_679J14_122_3096xU18 : FA_X1 port map( A => DP_OP_679J14_122_3096xn53, 
                           B => ashr_25xAx15x, CI => DP_OP_679J14_122_3096xn18,
                           CO => DP_OP_679J14_122_3096xn17, S => 
                           DP_OP_679J14_122_3096xn84);
   DP_OP_679J14_122_3096xU17 : FA_X1 port map( A => DP_OP_679J14_122_3096xn52, 
                           B => ashr_25xAx16x, CI => DP_OP_679J14_122_3096xn17,
                           CO => DP_OP_679J14_122_3096xn16, S => 
                           DP_OP_679J14_122_3096xn85);
   DP_OP_679J14_122_3096xU16 : FA_X1 port map( A => DP_OP_679J14_122_3096xn51, 
                           B => ashr_25xAx17x, CI => DP_OP_679J14_122_3096xn16,
                           CO => DP_OP_679J14_122_3096xn15, S => 
                           DP_OP_679J14_122_3096xn86);
   DP_OP_679J14_122_3096xU15 : FA_X1 port map( A => DP_OP_679J14_122_3096xn50, 
                           B => ashr_25xAx18x, CI => DP_OP_679J14_122_3096xn15,
                           CO => DP_OP_679J14_122_3096xn14, S => 
                           DP_OP_679J14_122_3096xn87);
   DP_OP_679J14_122_3096xU14 : FA_X1 port map( A => DP_OP_679J14_122_3096xn49, 
                           B => ashr_25xAx19x, CI => DP_OP_679J14_122_3096xn14,
                           CO => DP_OP_679J14_122_3096xn13, S => 
                           DP_OP_679J14_122_3096xn88);
   DP_OP_679J14_122_3096xU13 : FA_X1 port map( A => DP_OP_679J14_122_3096xn48, 
                           B => ashr_25xAx20x, CI => DP_OP_679J14_122_3096xn13,
                           CO => DP_OP_679J14_122_3096xn12, S => 
                           DP_OP_679J14_122_3096xn89);
   DP_OP_679J14_122_3096xU12 : FA_X1 port map( A => DP_OP_679J14_122_3096xn47, 
                           B => ashr_25xAx21x, CI => DP_OP_679J14_122_3096xn12,
                           CO => DP_OP_679J14_122_3096xn11, S => 
                           DP_OP_679J14_122_3096xn90);
   DP_OP_679J14_122_3096xU11 : FA_X1 port map( A => DP_OP_679J14_122_3096xn46, 
                           B => ashr_25xAx22x, CI => DP_OP_679J14_122_3096xn11,
                           CO => DP_OP_679J14_122_3096xn10, S => 
                           DP_OP_679J14_122_3096xn91);
   DP_OP_679J14_122_3096xU10 : FA_X1 port map( A => DP_OP_679J14_122_3096xn45, 
                           B => ashr_25xAx23x, CI => DP_OP_679J14_122_3096xn10,
                           CO => DP_OP_679J14_122_3096xn9, S => 
                           DP_OP_679J14_122_3096xn92);
   DP_OP_679J14_122_3096xU9 : FA_X1 port map( A => DP_OP_679J14_122_3096xn44, B
                           => ashr_25xAx24x, CI => DP_OP_679J14_122_3096xn9, CO
                           => DP_OP_679J14_122_3096xn8, S => 
                           DP_OP_679J14_122_3096xn93);
   DP_OP_679J14_122_3096xU8 : FA_X1 port map( A => DP_OP_679J14_122_3096xn43, B
                           => ashr_25xAx25x, CI => DP_OP_679J14_122_3096xn8, CO
                           => DP_OP_679J14_122_3096xn7, S => 
                           DP_OP_679J14_122_3096xn94);
   DP_OP_679J14_122_3096xU7 : FA_X1 port map( A => DP_OP_679J14_122_3096xn42, B
                           => ashr_25xAx26x, CI => DP_OP_679J14_122_3096xn7, CO
                           => DP_OP_679J14_122_3096xn6, S => 
                           DP_OP_679J14_122_3096xn95);
   DP_OP_679J14_122_3096xU6 : FA_X1 port map( A => DP_OP_679J14_122_3096xn41, B
                           => ashr_25xAx27x, CI => DP_OP_679J14_122_3096xn6, CO
                           => DP_OP_679J14_122_3096xn5, S => 
                           DP_OP_679J14_122_3096xn96);
   DP_OP_679J14_122_3096xU5 : FA_X1 port map( A => DP_OP_679J14_122_3096xn40, B
                           => ashr_25xAx28x, CI => DP_OP_679J14_122_3096xn5, CO
                           => DP_OP_679J14_122_3096xn4, S => 
                           DP_OP_679J14_122_3096xn97);
   DP_OP_679J14_122_3096xU4 : FA_X1 port map( A => DP_OP_679J14_122_3096xn39, B
                           => ashr_25xAx29x, CI => DP_OP_679J14_122_3096xn4, CO
                           => DP_OP_679J14_122_3096xn3, S => 
                           DP_OP_679J14_122_3096xn98);
   DP_OP_679J14_122_3096xU3 : FA_X1 port map( A => DP_OP_679J14_122_3096xn38, B
                           => ashr_25xAx30x, CI => DP_OP_679J14_122_3096xn3, CO
                           => DP_OP_679J14_122_3096xn2, S => 
                           DP_OP_679J14_122_3096xn99);
   DP_OP_719J14_125_1055xU33 : FA_X1 port map( A => DP_OP_719J14_125_1055xn134,
                           B => n7550, CI => DP_OP_719J14_125_1055xn68, CO => 
                           DP_OP_719J14_125_1055xn32, S => 
                           DP_OP_719J14_125_1055xn69);
   DP_OP_719J14_125_1055xU32 : FA_X1 port map( A => DP_OP_719J14_125_1055xn67, 
                           B => DP_OP_719J14_125_1055xn135, CI => 
                           DP_OP_719J14_125_1055xn32, CO => 
                           DP_OP_719J14_125_1055xn31, S => 
                           DP_OP_719J14_125_1055xn70);
   DP_OP_719J14_125_1055xU31 : FA_X1 port map( A => DP_OP_719J14_125_1055xn66, 
                           B => DP_OP_719J14_125_1055xn136, CI => 
                           DP_OP_719J14_125_1055xn31, CO => 
                           DP_OP_719J14_125_1055xn30, S => 
                           DP_OP_719J14_125_1055xn71);
   DP_OP_719J14_125_1055xU30 : FA_X1 port map( A => DP_OP_719J14_125_1055xn65, 
                           B => DP_OP_719J14_125_1055xn137, CI => 
                           DP_OP_719J14_125_1055xn30, CO => 
                           DP_OP_719J14_125_1055xn29, S => 
                           DP_OP_719J14_125_1055xn72);
   DP_OP_719J14_125_1055xU29 : FA_X1 port map( A => DP_OP_719J14_125_1055xn64, 
                           B => DP_OP_719J14_125_1055xn138, CI => 
                           DP_OP_719J14_125_1055xn29, CO => 
                           DP_OP_719J14_125_1055xn28, S => 
                           DP_OP_719J14_125_1055xn73);
   DP_OP_719J14_125_1055xU28 : FA_X1 port map( A => DP_OP_719J14_125_1055xn63, 
                           B => DP_OP_719J14_125_1055xn139, CI => 
                           DP_OP_719J14_125_1055xn28, CO => 
                           DP_OP_719J14_125_1055xn27, S => 
                           DP_OP_719J14_125_1055xn74);
   DP_OP_719J14_125_1055xU27 : FA_X1 port map( A => DP_OP_719J14_125_1055xn62, 
                           B => DP_OP_719J14_125_1055xn140, CI => 
                           DP_OP_719J14_125_1055xn27, CO => 
                           DP_OP_719J14_125_1055xn26, S => 
                           DP_OP_719J14_125_1055xn75);
   DP_OP_719J14_125_1055xU26 : FA_X1 port map( A => DP_OP_719J14_125_1055xn61, 
                           B => DP_OP_719J14_125_1055xn141, CI => 
                           DP_OP_719J14_125_1055xn26, CO => 
                           DP_OP_719J14_125_1055xn25, S => 
                           DP_OP_719J14_125_1055xn76);
   DP_OP_719J14_125_1055xU25 : FA_X1 port map( A => DP_OP_719J14_125_1055xn60, 
                           B => DP_OP_719J14_125_1055xn142, CI => 
                           DP_OP_719J14_125_1055xn25, CO => 
                           DP_OP_719J14_125_1055xn24, S => 
                           DP_OP_719J14_125_1055xn77);
   DP_OP_719J14_125_1055xU24 : FA_X1 port map( A => DP_OP_719J14_125_1055xn59, 
                           B => DP_OP_719J14_125_1055xn143, CI => 
                           DP_OP_719J14_125_1055xn24, CO => 
                           DP_OP_719J14_125_1055xn23, S => 
                           DP_OP_719J14_125_1055xn78);
   DP_OP_719J14_125_1055xU23 : FA_X1 port map( A => DP_OP_719J14_125_1055xn58, 
                           B => DP_OP_719J14_125_1055xn144, CI => 
                           DP_OP_719J14_125_1055xn23, CO => 
                           DP_OP_719J14_125_1055xn22, S => 
                           DP_OP_719J14_125_1055xn79);
   DP_OP_719J14_125_1055xU22 : FA_X1 port map( A => DP_OP_719J14_125_1055xn57, 
                           B => DP_OP_719J14_125_1055xn145, CI => 
                           DP_OP_719J14_125_1055xn22, CO => 
                           DP_OP_719J14_125_1055xn21, S => 
                           DP_OP_719J14_125_1055xn80);
   DP_OP_719J14_125_1055xU21 : FA_X1 port map( A => DP_OP_719J14_125_1055xn56, 
                           B => DP_OP_719J14_125_1055xn146, CI => 
                           DP_OP_719J14_125_1055xn21, CO => 
                           DP_OP_719J14_125_1055xn20, S => 
                           DP_OP_719J14_125_1055xn81);
   DP_OP_719J14_125_1055xU20 : FA_X1 port map( A => DP_OP_719J14_125_1055xn55, 
                           B => DP_OP_719J14_125_1055xn147, CI => 
                           DP_OP_719J14_125_1055xn20, CO => 
                           DP_OP_719J14_125_1055xn19, S => 
                           DP_OP_719J14_125_1055xn82);
   DP_OP_719J14_125_1055xU19 : FA_X1 port map( A => DP_OP_719J14_125_1055xn54, 
                           B => DP_OP_719J14_125_1055xn148, CI => 
                           DP_OP_719J14_125_1055xn19, CO => 
                           DP_OP_719J14_125_1055xn18, S => 
                           DP_OP_719J14_125_1055xn83);
   DP_OP_719J14_125_1055xU18 : FA_X1 port map( A => DP_OP_719J14_125_1055xn53, 
                           B => DP_OP_719J14_125_1055xn149, CI => 
                           DP_OP_719J14_125_1055xn18, CO => 
                           DP_OP_719J14_125_1055xn17, S => 
                           DP_OP_719J14_125_1055xn84);
   DP_OP_719J14_125_1055xU17 : FA_X1 port map( A => DP_OP_719J14_125_1055xn52, 
                           B => DP_OP_719J14_125_1055xn150, CI => 
                           DP_OP_719J14_125_1055xn17, CO => 
                           DP_OP_719J14_125_1055xn16, S => 
                           DP_OP_719J14_125_1055xn85);
   DP_OP_719J14_125_1055xU16 : FA_X1 port map( A => DP_OP_719J14_125_1055xn51, 
                           B => DP_OP_719J14_125_1055xn151, CI => 
                           DP_OP_719J14_125_1055xn16, CO => 
                           DP_OP_719J14_125_1055xn15, S => 
                           DP_OP_719J14_125_1055xn86);
   DP_OP_719J14_125_1055xU15 : FA_X1 port map( A => DP_OP_719J14_125_1055xn50, 
                           B => DP_OP_719J14_125_1055xn152, CI => 
                           DP_OP_719J14_125_1055xn15, CO => 
                           DP_OP_719J14_125_1055xn14, S => 
                           DP_OP_719J14_125_1055xn87);
   DP_OP_719J14_125_1055xU14 : FA_X1 port map( A => DP_OP_719J14_125_1055xn49, 
                           B => DP_OP_719J14_125_1055xn153, CI => 
                           DP_OP_719J14_125_1055xn14, CO => 
                           DP_OP_719J14_125_1055xn13, S => 
                           DP_OP_719J14_125_1055xn88);
   DP_OP_719J14_125_1055xU13 : FA_X1 port map( A => DP_OP_719J14_125_1055xn48, 
                           B => DP_OP_719J14_125_1055xn154, CI => 
                           DP_OP_719J14_125_1055xn13, CO => 
                           DP_OP_719J14_125_1055xn12, S => 
                           DP_OP_719J14_125_1055xn89);
   DP_OP_719J14_125_1055xU12 : FA_X1 port map( A => DP_OP_719J14_125_1055xn47, 
                           B => DP_OP_719J14_125_1055xn155, CI => 
                           DP_OP_719J14_125_1055xn12, CO => 
                           DP_OP_719J14_125_1055xn11, S => 
                           DP_OP_719J14_125_1055xn90);
   DP_OP_719J14_125_1055xU11 : FA_X1 port map( A => DP_OP_719J14_125_1055xn46, 
                           B => DP_OP_719J14_125_1055xn156, CI => 
                           DP_OP_719J14_125_1055xn11, CO => 
                           DP_OP_719J14_125_1055xn10, S => 
                           DP_OP_719J14_125_1055xn91);
   DP_OP_719J14_125_1055xU10 : FA_X1 port map( A => DP_OP_719J14_125_1055xn45, 
                           B => DP_OP_719J14_125_1055xn157, CI => 
                           DP_OP_719J14_125_1055xn10, CO => 
                           DP_OP_719J14_125_1055xn9, S => 
                           DP_OP_719J14_125_1055xn92);
   DP_OP_719J14_125_1055xU9 : FA_X1 port map( A => DP_OP_719J14_125_1055xn44, B
                           => DP_OP_719J14_125_1055xn158, CI => 
                           DP_OP_719J14_125_1055xn9, CO => 
                           DP_OP_719J14_125_1055xn8, S => 
                           DP_OP_719J14_125_1055xn93);
   DP_OP_719J14_125_1055xU8 : FA_X1 port map( A => DP_OP_719J14_125_1055xn43, B
                           => DP_OP_719J14_125_1055xn159, CI => 
                           DP_OP_719J14_125_1055xn8, CO => 
                           DP_OP_719J14_125_1055xn7, S => 
                           DP_OP_719J14_125_1055xn94);
   DP_OP_719J14_125_1055xU7 : FA_X1 port map( A => DP_OP_719J14_125_1055xn42, B
                           => DP_OP_719J14_125_1055xn160, CI => 
                           DP_OP_719J14_125_1055xn7, CO => 
                           DP_OP_719J14_125_1055xn6, S => 
                           DP_OP_719J14_125_1055xn95);
   DP_OP_719J14_125_1055xU6 : FA_X1 port map( A => DP_OP_719J14_125_1055xn41, B
                           => DP_OP_719J14_125_1055xn161, CI => 
                           DP_OP_719J14_125_1055xn6, CO => 
                           DP_OP_719J14_125_1055xn5, S => 
                           DP_OP_719J14_125_1055xn96);
   DP_OP_719J14_125_1055xU5 : FA_X1 port map( A => DP_OP_719J14_125_1055xn40, B
                           => DP_OP_719J14_125_1055xn162, CI => 
                           DP_OP_719J14_125_1055xn5, CO => 
                           DP_OP_719J14_125_1055xn4, S => 
                           DP_OP_719J14_125_1055xn97);
   DP_OP_719J14_125_1055xU4 : FA_X1 port map( A => DP_OP_719J14_125_1055xn39, B
                           => DP_OP_719J14_125_1055xn163, CI => 
                           DP_OP_719J14_125_1055xn4, CO => 
                           DP_OP_719J14_125_1055xn3, S => 
                           DP_OP_719J14_125_1055xn98);
   DP_OP_719J14_125_1055xU3 : FA_X1 port map( A => DP_OP_719J14_125_1055xn38, B
                           => DP_OP_719J14_125_1055xn164, CI => 
                           DP_OP_719J14_125_1055xn3, CO => 
                           DP_OP_719J14_125_1055xn2, S => 
                           DP_OP_719J14_125_1055xn99);
   intadd_25xU30 : FA_X1 port map( A => IF_ISAxpcReg_signal_2_port, B => 
                           intadd_25xBx0x, CI => intadd_25xCI, CO => 
                           intadd_25xn29, S => intadd_25xSUMx0x);
   intadd_25xU29 : FA_X1 port map( A => IF_ISAxpcReg_signal_3_port, B => 
                           ashr_25xSHx3x, CI => intadd_25xn29, CO => 
                           intadd_25xn28, S => intadd_25xSUMx1x);
   intadd_25xU28 : FA_X1 port map( A => IF_ISAxpcReg_signal_4_port, B => 
                           ashr_25xSHx4x, CI => intadd_25xn28, CO => 
                           intadd_25xn27, S => intadd_25xSUMx2x);
   intadd_25xU27 : FA_X1 port map( A => IF_ISAxpcReg_signal_5_port, B => 
                           add_x_26xBx5x, CI => intadd_25xn27, CO => 
                           intadd_25xn26, S => intadd_25xSUMx3x);
   intadd_25xU26 : FA_X1 port map( A => IF_ISAxpcReg_signal_6_port, B => 
                           add_x_26xBx6x, CI => intadd_25xn26, CO => 
                           intadd_25xn25, S => intadd_25xSUMx4x);
   intadd_25xU25 : FA_X1 port map( A => IF_ISAxpcReg_signal_7_port, B => 
                           add_x_26xBx7x, CI => intadd_25xn25, CO => 
                           intadd_25xn24, S => intadd_25xSUMx5x);
   intadd_25xU24 : FA_X1 port map( A => IF_ISAxpcReg_signal_8_port, B => 
                           add_x_26xBx8x, CI => intadd_25xn24, CO => 
                           intadd_25xn23, S => intadd_25xSUMx6x);
   intadd_25xU23 : FA_X1 port map( A => IF_ISAxpcReg_signal_9_port, B => 
                           add_x_26xBx9x, CI => intadd_25xn23, CO => 
                           intadd_25xn22, S => intadd_25xSUMx7x);
   intadd_25xU22 : FA_X1 port map( A => IF_ISAxpcReg_signal_10_port, B => 
                           add_x_26xBx10x, CI => intadd_25xn22, CO => 
                           intadd_25xn21, S => intadd_25xSUMx8x);
   intadd_25xU21 : FA_X1 port map( A => IF_ISAxpcReg_signal_11_port, B => 
                           add_x_26xBx11x, CI => intadd_25xn21, CO => 
                           intadd_25xn20, S => intadd_25xSUMx9x);
   intadd_25xU20 : FA_X1 port map( A => IF_ISAxpcReg_signal_12_port, B => 
                           add_x_26xBx12x, CI => intadd_25xn20, CO => 
                           intadd_25xn19, S => intadd_25xSUMx10x);
   intadd_25xU19 : FA_X1 port map( A => IF_ISAxpcReg_signal_13_port, B => 
                           add_x_26xBx13x, CI => intadd_25xn19, CO => 
                           intadd_25xn18, S => intadd_25xSUMx11x);
   intadd_25xU18 : FA_X1 port map( A => IF_ISAxpcReg_signal_14_port, B => 
                           add_x_26xBx14x, CI => intadd_25xn18, CO => 
                           intadd_25xn17, S => intadd_25xSUMx12x);
   intadd_25xU17 : FA_X1 port map( A => IF_ISAxpcReg_signal_15_port, B => 
                           add_x_26xBx15x, CI => intadd_25xn17, CO => 
                           intadd_25xn16, S => intadd_25xSUMx13x);
   intadd_25xU16 : FA_X1 port map( A => IF_ISAxpcReg_signal_16_port, B => 
                           add_x_26xBx16x, CI => intadd_25xn16, CO => 
                           intadd_25xn15, S => intadd_25xSUMx14x);
   intadd_25xU15 : FA_X1 port map( A => IF_ISAxpcReg_signal_17_port, B => 
                           add_x_26xBx17x, CI => intadd_25xn15, CO => 
                           intadd_25xn14, S => intadd_25xSUMx15x);
   intadd_25xU14 : FA_X1 port map( A => IF_ISAxpcReg_signal_18_port, B => 
                           add_x_26xBx18x, CI => intadd_25xn14, CO => 
                           intadd_25xn13, S => intadd_25xSUMx16x);
   intadd_25xU13 : FA_X1 port map( A => IF_ISAxpcReg_signal_19_port, B => 
                           add_x_26xBx19x, CI => intadd_25xn13, CO => 
                           intadd_25xn12, S => intadd_25xSUMx17x);
   intadd_25xU12 : FA_X1 port map( A => IF_ISAxpcReg_signal_20_port, B => 
                           add_x_26xBx20x, CI => intadd_25xn12, CO => 
                           intadd_25xn11, S => intadd_25xSUMx18x);
   intadd_25xU11 : FA_X1 port map( A => IF_ISAxpcReg_signal_21_port, B => 
                           add_x_26xBx21x, CI => intadd_25xn11, CO => 
                           intadd_25xn10, S => intadd_25xSUMx19x);
   intadd_25xU10 : FA_X1 port map( A => IF_ISAxpcReg_signal_22_port, B => 
                           add_x_26xBx22x, CI => intadd_25xn10, CO => 
                           intadd_25xn9, S => intadd_25xSUMx20x);
   intadd_25xU9 : FA_X1 port map( A => IF_ISAxpcReg_signal_23_port, B => 
                           add_x_26xBx23x, CI => intadd_25xn9, CO => 
                           intadd_25xn8, S => intadd_25xSUMx21x);
   intadd_25xU8 : FA_X1 port map( A => IF_ISAxpcReg_signal_24_port, B => 
                           add_x_26xBx24x, CI => intadd_25xn8, CO => 
                           intadd_25xn7, S => intadd_25xSUMx22x);
   intadd_25xU7 : FA_X1 port map( A => IF_ISAxpcReg_signal_25_port, B => 
                           add_x_26xBx25x, CI => intadd_25xn7, CO => 
                           intadd_25xn6, S => intadd_25xSUMx23x);
   intadd_25xU6 : FA_X1 port map( A => IF_ISAxpcReg_signal_26_port, B => 
                           add_x_26xBx26x, CI => intadd_25xn6, CO => 
                           intadd_25xn5, S => intadd_25xSUMx24x);
   intadd_25xU5 : FA_X1 port map( A => IF_ISAxpcReg_signal_27_port, B => 
                           add_x_26xBx27x, CI => intadd_25xn5, CO => 
                           intadd_25xn4, S => intadd_25xSUMx25x);
   intadd_25xU4 : FA_X1 port map( A => IF_ISAxpcReg_signal_28_port, B => 
                           add_x_26xBx28x, CI => intadd_25xn4, CO => 
                           intadd_25xn3, S => intadd_25xSUMx26x);
   intadd_25xU3 : FA_X1 port map( A => IF_ISAxpcReg_signal_29_port, B => 
                           add_x_26xBx29x, CI => intadd_25xn3, CO => 
                           intadd_25xn2, S => intadd_25xSUMx27x);
   intadd_25xU2 : FA_X1 port map( A => IF_ISAxpcReg_signal_30_port, B => 
                           add_x_26xBx30x, CI => intadd_25xn2, CO => 
                           intadd_25xn1, S => intadd_25xSUMx28x);
   intadd_26xU9 : FA_X1 port map( A => intadd_26xAx0x, B => intadd_26xBx0x, CI 
                           => intadd_26xCI, CO => intadd_26xn8, S => 
                           intadd_26xSUMx0x);
   intadd_26xU8 : FA_X1 port map( A => intadd_26xAx1x, B => intadd_26xBx1x, CI 
                           => intadd_26xn8, CO => intadd_26xn7, S => 
                           intadd_26xSUMx1x);
   intadd_26xU7 : FA_X1 port map( A => intadd_26xAx2x, B => intadd_26xBx2x, CI 
                           => intadd_26xn7, CO => intadd_26xn6, S => 
                           intadd_26xSUMx2x);
   intadd_26xU6 : FA_X1 port map( A => intadd_26xAx3x, B => intadd_26xBx3x, CI 
                           => intadd_26xn6, CO => intadd_26xn5, S => 
                           intadd_26xSUMx3x);
   intadd_26xU5 : FA_X1 port map( A => intadd_26xAx4x, B => intadd_26xBx4x, CI 
                           => intadd_26xn5, CO => intadd_26xn4, S => 
                           intadd_26xSUMx4x);
   intadd_26xU4 : FA_X1 port map( A => intadd_26xAx5x, B => intadd_26xBx5x, CI 
                           => intadd_26xn4, CO => intadd_26xn3, S => 
                           intadd_26xSUMx5x);
   intadd_26xU3 : FA_X1 port map( A => intadd_26xAx6x, B => intadd_26xBx6x, CI 
                           => intadd_26xn3, CO => intadd_26xn2, S => 
                           intadd_26xSUMx6x);
   intadd_26xU2 : FA_X1 port map( A => intadd_26xAx7x, B => intadd_26xBx7x, CI 
                           => intadd_26xn2, CO => intadd_26xn1, S => 
                           intadd_26xSUMx7x);
   intadd_27xU5 : FA_X1 port map( A => intadd_27xAx0x, B => intadd_27xBx0x, CI 
                           => intadd_27xCI, CO => intadd_27xn4, S => 
                           intadd_27xSUMx0x);
   intadd_27xU4 : FA_X1 port map( A => intadd_27xAx1x, B => intadd_27xBx1x, CI 
                           => intadd_27xn4, CO => intadd_27xn3, S => 
                           intadd_27xSUMx1x);
   intadd_27xU3 : FA_X1 port map( A => intadd_27xAx2x, B => intadd_27xBx2x, CI 
                           => intadd_27xn3, CO => intadd_27xn2, S => 
                           intadd_27xSUMx2x);
   intadd_27xU2 : FA_X1 port map( A => intadd_27xAx3x, B => intadd_27xBx3x, CI 
                           => intadd_27xn2, CO => intadd_27xn1, S => 
                           intadd_27xSUMx3x);
   intadd_28xU4 : FA_X1 port map( A => intadd_28xAx0x, B => intadd_28xBx0x, CI 
                           => intadd_28xCI, CO => intadd_28xn3, S => 
                           intadd_28xSUMx0x);
   intadd_28xU3 : FA_X1 port map( A => intadd_28xAx1x, B => intadd_28xBx1x, CI 
                           => intadd_28xn3, CO => intadd_28xn2, S => 
                           intadd_28xSUMx1x);
   intadd_28xU2 : FA_X1 port map( A => intadd_28xAx2x, B => intadd_28xBx2x, CI 
                           => intadd_28xn2, CO => intadd_28xn1, S => 
                           intadd_28xSUMx2x);
   intadd_29xU4 : FA_X1 port map( A => intadd_29xAx0x, B => intadd_29xBx0x, CI 
                           => intadd_29xCI, CO => intadd_29xn3, S => 
                           intadd_29xSUMx0x);
   intadd_29xU3 : FA_X1 port map( A => intadd_29xAx1x, B => intadd_29xBx1x, CI 
                           => intadd_29xn3, CO => intadd_29xn2, S => 
                           intadd_29xSUMx1x);
   intadd_29xU2 : FA_X1 port map( A => intadd_29xAx2x, B => intadd_29xBx2x, CI 
                           => intadd_29xn2, CO => intadd_29xn1, S => 
                           intadd_29xSUMx2x);
   U3775 : AOI21_X2 port map( B1 => n7435, B2 => n7349, A => n6386, ZN => n7353
                           );
   U3776 : NOR3_X4 port map( A1 => n5716, A2 => n5719, A3 => n5715, ZN => n7320
                           );
   U3777 : NAND2_X2 port map( A1 => n3564, A2 => n3563, ZN => ashr_25xSHx3x);
   U3778 : OR2_X1 port map( A1 => n3622, A2 => n3621, ZN => n3558);
   U3779 : INV_X1 port map( A => n5441, ZN => n5658);
   U3780 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(0), A2 => 
                           fromMemoryPortxLOADEDDATAx(1), ZN => n3559);
   U3781 : NOR4_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(2), A2 => 
                           fromMemoryPortxLOADEDDATAx(4), A3 => 
                           fromMemoryPortxLOADEDDATAx(3), A4 => n3559, ZN => 
                           n3561);
   U3782 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(5), A2 => n3561, 
                           ZN => n7446);
   U3783 : NAND2_X1 port map( A1 => n7446, A2 => fromMemoryPortxLOADEDDATAx(10)
                           , ZN => n3564);
   U3784 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(2), A2 => 
                           fromMemoryPortxLOADEDDATAx(6), ZN => n5748);
   U3785 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(4), ZN => n6270);
   U3786 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(5), A2 => n6270,
                           ZN => n5749);
   U3787 : NOR3_X1 port map( A1 => n5748, A2 => n3559, A3 => n5749, ZN => n7445
                           );
   U3788 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(5), ZN => n3560);
   U3789 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(6), ZN => n6361);
   U3790 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(3), ZN => n5739);
   U3791 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(4), A2 => n6361,
                           A3 => n5739, ZN => n5755);
   U3792 : NOR2_X2 port map( A1 => n3559, A2 => n5755, ZN => n7118);
   U3793 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(2), ZN => n6157);
   U3794 : NAND2_X1 port map( A1 => n7118, A2 => n6157, ZN => n5681);
   U3795 : INV_X1 port map( A => n5681, ZN => n3565);
   U3796 : NAND2_X1 port map( A1 => n3560, A2 => n3565, ZN => n5715);
   U3797 : NAND2_X1 port map( A1 => n3561, A2 => n6361, ZN => n7490);
   U3798 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(5), A2 => n7490, 
                           ZN => n7444);
   U3799 : INV_X1 port map( A => n7444, ZN => n7452);
   U3800 : NAND2_X1 port map( A1 => n5715, A2 => n7452, ZN => n3562);
   U3801 : OR2_X1 port map( A1 => n7445, A2 => n3562, ZN => n3723);
   U3802 : NAND2_X1 port map( A1 => n3723, A2 => fromMemoryPortxLOADEDDATAx(23)
                           , ZN => n3563);
   U3803 : INV_X1 port map( A => n7445, ZN => n3570);
   U3804 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(14), A2 => 
                           fromMemoryPortxLOADEDDATAx(12), ZN => n5954);
   U3805 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(13), A2 => n5954,
                           ZN => n3601);
   U3806 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(5), A2 => n3565, 
                           ZN => n6020);
   U3807 : NOR4_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(29), A2 => 
                           fromMemoryPortxLOADEDDATAx(25), A3 => 
                           fromMemoryPortxLOADEDDATAx(27), A4 => 
                           fromMemoryPortxLOADEDDATAx(26), ZN => n3566);
   U3808 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(28), ZN => n7249);
   U3809 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(31), ZN => n7440);
   U3810 : NAND3_X1 port map( A1 => n3566, A2 => n7249, A3 => n7440, ZN => 
                           n3597);
   U3811 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(30), ZN => n7362);
   U3812 : NOR2_X1 port map( A1 => n3597, A2 => n7362, ZN => n3589);
   U3813 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(13), ZN => n6670);
   U3814 : AND2_X1 port map( A1 => n3589, A2 => n6670, ZN => n3573);
   U3815 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(12), B2 => 
                           fromMemoryPortxLOADEDDATAx(14), A => n5954, ZN => 
                           n3590);
   U3816 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(14), ZN => n6716);
   U3817 : NAND2_X1 port map( A1 => n6670, A2 => n6716, ZN => n3586);
   U3818 : OAI21_X1 port map( B1 => n3573, B2 => n3590, A => n3586, ZN => n3567
                           );
   U3819 : AND2_X1 port map( A1 => n7446, A2 => fromMemoryPortxLOADEDDATAx(6), 
                           ZN => n4768);
   U3820 : INV_X1 port map( A => n4768, ZN => n7457);
   U3821 : OAI22_X1 port map( A1 => n5715, A2 => n3567, B1 => n7457, B2 => 
                           n3590, ZN => n3568);
   U3822 : AOI21_X1 port map( B1 => n3601, B2 => n6020, A => n3568, ZN => n3569
                           );
   U3823 : AND2_X1 port map( A1 => n7446, A2 => n6361, ZN => n7460);
   U3824 : INV_X1 port map( A => n7460, ZN => n5963);
   U3825 : NAND3_X1 port map( A1 => n3570, A2 => n3569, A3 => n5963, ZN => 
                           n5702);
   U3826 : INV_X1 port map( A => n5702, ZN => n3611);
   U3827 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(30), A2 => n3597,
                           ZN => n3591);
   U3828 : INV_X1 port map( A => n3586, ZN => n5955);
   U3829 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(12), ZN => n5741);
   U3830 : NAND2_X1 port map( A1 => n5955, A2 => n5741, ZN => n3598);
   U3831 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(14), A2 => n6670
                           , ZN => n3575);
   U3832 : OAI21_X1 port map( B1 => n3591, B2 => n3598, A => n3575, ZN => n3571
                           );
   U3833 : INV_X1 port map( A => n3571, ZN => n3574);
   U3834 : INV_X1 port map( A => n6020, ZN => n5710);
   U3835 : INV_X1 port map( A => n5715, ZN => n6022);
   U3836 : OAI21_X1 port map( B1 => n3586, B2 => fromMemoryPortxLOADEDDATAx(12)
                           , A => n6022, ZN => n3584);
   U3837 : NAND2_X1 port map( A1 => n6670, A2 => n5741, ZN => n3572);
   U3838 : OAI21_X1 port map( B1 => n6716, B2 => n3573, A => n3572, ZN => n3585
                           );
   U3839 : NAND2_X1 port map( A1 => n6670, A2 => n3585, ZN => n3577);
   U3840 : INV_X1 port map( A => n7446, ZN => n3595);
   U3841 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(13), A2 => n6716
                           , ZN => n5444);
   U3842 : OAI222_X1 port map( A1 => n3574, A2 => n5710, B1 => n3584, B2 => 
                           n3577, C1 => n3595, C2 => n5444, ZN => n3608);
   U3843 : AND2_X1 port map( A1 => n7118, A2 => fromMemoryPortxLOADEDDATAx(2), 
                           ZN => n5694);
   U3844 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(13), A2 => n5741
                           , B1 => fromMemoryPortxLOADEDDATAx(12), B2 => n6670,
                           ZN => n3579);
   U3845 : INV_X1 port map( A => n3575, ZN => n3592);
   U3846 : NAND2_X1 port map( A1 => n3592, A2 => n3597, ZN => n3576);
   U3847 : AOI22_X1 port map( A1 => n6022, A2 => n3577, B1 => n6020, B2 => 
                           n3576, ZN => n3578);
   U3848 : AOI21_X1 port map( B1 => n3579, B2 => n5444, A => n3578, ZN => n3580
                           );
   U3849 : AOI211_X1 port map( C1 => fromMemoryPortxLOADEDDATAx(5), C2 => n5694
                           , A => n7460, B => n3580, ZN => n3607);
   U3850 : INV_X1 port map( A => n3607, ZN => n3613);
   U3851 : OR2_X1 port map( A1 => n3608, A2 => n3613, ZN => n3603);
   U3852 : NOR2_X1 port map( A1 => n3611, A2 => n3603, ZN => n5637);
   U3853 : AOI21_X1 port map( B1 => n4768, B2 => n3590, A => n7445, ZN => n3583
                           );
   U3854 : INV_X1 port map( A => n5444, ZN => n3581);
   U3855 : OAI221_X1 port map( B1 => n3581, B2 => n3592, C1 => n3581, C2 => 
                           fromMemoryPortxLOADEDDATAx(12), A => n6020, ZN => 
                           n3582);
   U3856 : OAI211_X1 port map( C1 => n3585, C2 => n3584, A => n3583, B => n3582
                           , ZN => n3621);
   U3857 : OAI21_X1 port map( B1 => n6670, B2 => n5954, A => n3586, ZN => n3587
                           );
   U3858 : INV_X1 port map( A => n3587, ZN => n3588);
   U3859 : AOI221_X1 port map( B1 => n3589, B2 => n3588, C1 => n5741, C2 => 
                           n3588, A => n5710, ZN => n3599);
   U3860 : AOI211_X1 port map( C1 => n3592, C2 => n3591, A => n5715, B => n3590
                           , ZN => n3593);
   U3861 : INV_X1 port map( A => n3593, ZN => n3594);
   U3862 : OAI21_X1 port map( B1 => n3595, B2 => n5741, A => n3594, ZN => n3596
                           );
   U3863 : AOI222_X1 port map( A1 => n3599, A2 => n3598, B1 => n3599, B2 => 
                           n3597, C1 => n3598, C2 => n3596, ZN => n3600);
   U3864 : INV_X1 port map( A => n3600, ZN => n3633);
   U3865 : NOR2_X1 port map( A1 => n3621, A2 => n3633, ZN => n3609);
   U3866 : OAI21_X1 port map( B1 => n3601, B2 => n7457, A => n5710, ZN => n3602
                           );
   U3867 : NOR2_X1 port map( A1 => n7460, A2 => n3602, ZN => n3610);
   U3868 : NOR2_X1 port map( A1 => n5702, A2 => n3603, ZN => n3612);
   U3869 : NAND2_X1 port map( A1 => n3612, A2 => n3621, ZN => n5639);
   U3870 : INV_X1 port map( A => n5637, ZN => n3604);
   U3871 : INV_X1 port map( A => n3621, ZN => n5636);
   U3872 : NAND2_X1 port map( A1 => n3633, A2 => n5636, ZN => n3616);
   U3873 : NOR2_X1 port map( A1 => n3604, A2 => n3616, ZN => n3635);
   U3874 : INV_X1 port map( A => n3635, ZN => n3605);
   U3875 : NAND2_X1 port map( A1 => n5639, A2 => n3605, ZN => n3606);
   U3876 : AOI22_X1 port map( A1 => n5637, A2 => n3609, B1 => n3610, B2 => 
                           n3606, ZN => n3630);
   U3877 : NAND2_X1 port map( A1 => n3600, A2 => n3610, ZN => n3615);
   U3878 : NOR2_X1 port map( A1 => n3600, A2 => n3610, ZN => n3620);
   U3879 : INV_X1 port map( A => n3620, ZN => n3625);
   U3880 : NAND2_X1 port map( A1 => n3615, A2 => n3625, ZN => n3623);
   U3881 : INV_X1 port map( A => n3623, ZN => n3619);
   U3882 : NOR2_X1 port map( A1 => n5636, A2 => n3607, ZN => n3637);
   U3883 : NAND2_X1 port map( A1 => n3609, A2 => n3608, ZN => n3626);
   U3884 : AOI21_X1 port map( B1 => n3611, B2 => n3610, A => n3626, ZN => n3618
                           );
   U3885 : INV_X1 port map( A => n3612, ZN => n3622);
   U3886 : NOR2_X1 port map( A1 => n3620, A2 => n5702, ZN => n3614);
   U3887 : NAND2_X1 port map( A1 => n5636, A2 => n3613, ZN => n5701);
   U3888 : OR2_X1 port map( A1 => n3614, A2 => n5701, ZN => n3624);
   U3889 : AOI21_X2 port map( B1 => n5702, B2 => n3615, A => n3624, ZN => n7251
                           );
   U3890 : INV_X1 port map( A => n7251, ZN => n7387);
   U3891 : OAI21_X1 port map( B1 => n3616, B2 => n3622, A => n7387, ZN => n3617
                           );
   U3892 : AOI211_X1 port map( C1 => n3619, C2 => n3637, A => n3618, B => n3617
                           , ZN => n5699);
   U3893 : NAND2_X1 port map( A1 => n3630, A2 => n5699, ZN => n5630);
   U3894 : NAND2_X1 port map( A1 => n3620, A2 => n5702, ZN => n3636);
   U3895 : NOR2_X1 port map( A1 => n5701, A2 => n3636, ZN => n3631);
   U3896 : OAI21_X1 port map( B1 => n3624, B2 => n3623, A => n3558, ZN => n3638
                           );
   U3897 : INV_X1 port map( A => n3637, ZN => n3628);
   U3898 : XNOR2_X1 port map( A => n5702, B => n3625, ZN => n3627);
   U3899 : OAI22_X1 port map( A1 => n3628, A2 => n3627, B1 => n5702, B2 => 
                           n3626, ZN => n3629);
   U3900 : NOR3_X1 port map( A1 => n3631, A2 => n3638, A3 => n3629, ZN => n5632
                           );
   U3901 : NAND2_X1 port map( A1 => n3630, A2 => n5632, ZN => n5698);
   U3902 : NAND2_X1 port map( A1 => n5630, A2 => n5698, ZN => n5719);
   U3903 : INV_X1 port map( A => n3631, ZN => n3632);
   U3904 : OAI21_X1 port map( B1 => n3633, B2 => n5639, A => n3632, ZN => n3634
                           );
   U3905 : AOI211_X1 port map( C1 => n3637, C2 => n3636, A => n3635, B => n3634
                           , ZN => n5692);
   U3906 : NOR2_X1 port map( A1 => n3638, A2 => n7251, ZN => n5716);
   U3907 : AND2_X1 port map( A1 => n5692, A2 => n5716, ZN => n5690);
   U3908 : INV_X1 port map( A => n5690, ZN => n5697);
   U3909 : NOR2_X1 port map( A1 => n5719, A2 => n5697, ZN => n5680);
   U3910 : INV_X1 port map( A => n5680, ZN => n3639);
   U3911 : NOR2_X1 port map( A1 => n3639, A2 => n5710, ZN => n4242);
   U3912 : CLKBUF_X1 port map( A => n4242, Z => n7550);
   U3913 : NAND2_X1 port map( A1 => n7446, A2 => fromMemoryPortxLOADEDDATAx(9),
                           ZN => n3641);
   U3914 : NAND2_X1 port map( A1 => n3723, A2 => fromMemoryPortxLOADEDDATAx(22)
                           , ZN => n3640);
   U3915 : NAND2_X1 port map( A1 => n3641, A2 => n3640, ZN => n6456);
   U3916 : CLKBUF_X1 port map( A => n6456, Z => intadd_25xBx0x);
   U3917 : NAND2_X1 port map( A1 => n7446, A2 => fromMemoryPortxLOADEDDATAx(8),
                           ZN => n3643);
   U3918 : NAND2_X1 port map( A1 => n3723, A2 => fromMemoryPortxLOADEDDATAx(21)
                           , ZN => n3642);
   U3919 : NAND2_X1 port map( A1 => n3643, A2 => n3642, ZN => n7259);
   U3920 : CLKBUF_X1 port map( A => n7259, Z => n7416);
   U3921 : INV_X1 port map( A => n7416, ZN => intadd_29xBx0x);
   U3922 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(13), A2 => n5741,
                           ZN => n3645);
   U3923 : NAND2_X1 port map( A1 => n7445, A2 => n5739, ZN => n5110);
   U3924 : AND2_X1 port map( A1 => n7490, A2 => n5110, ZN => n3644);
   U3925 : OAI21_X1 port map( B1 => n5715, B2 => n3645, A => n3644, ZN => n4533
                           );
   U3926 : OR3_X1 port map( A1 => n4768, A2 => n7445, A3 => n4533, ZN => n4944)
                           ;
   U3927 : NAND2_X1 port map( A1 => n4944, A2 => fromMemoryPortxLOADEDDATAx(31)
                           , ZN => n4504);
   U3928 : INV_X1 port map( A => n5694, ZN => n4534);
   U3929 : NAND2_X1 port map( A1 => n4504, A2 => n4534, ZN => n4445);
   U3930 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(27), ZN => n3646);
   U3931 : NAND2_X1 port map( A1 => n4504, A2 => n3646, ZN => n3647);
   U3932 : AND2_X1 port map( A1 => n4445, A2 => n3647, ZN => add_x_26xBx27x);
   U3933 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(27), A2 => n4944,
                           ZN => add_x_26xBx7x);
   U3934 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(28), A2 => n4944,
                           ZN => add_x_26xBx8x);
   U3935 : INV_X1 port map( A => rst, ZN => n7523);
   U3936 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx26x, A2 => n7523, ZN => 
                           IF_RegsxN686);
   U3937 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx10x, A2 => n7523, ZN => 
                           IF_RegsxN670);
   U3938 : CLKBUF_X1 port map( A => n7523, Z => n7520);
   U3939 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx28x, A2 => n7520, ZN => 
                           IF_RegsxN688);
   U3940 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx12x, A2 => n7523, ZN => 
                           IF_RegsxN672);
   U3941 : CLKBUF_X1 port map( A => n7523, Z => n7509);
   U3942 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx11x, A2 => n7509, ZN => 
                           IF_RegsxN671);
   U3943 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx8x, A2 => n7509, ZN => 
                           IF_RegsxN668);
   U3944 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx22x, A2 => n7523, ZN => 
                           IF_RegsxN682);
   U3945 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx20x, A2 => n7523, ZN => 
                           IF_RegsxN680);
   U3946 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx27x, A2 => n7509, ZN => 
                           IF_RegsxN687);
   U3947 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx23x, A2 => n7509, ZN => 
                           IF_RegsxN683);
   U3948 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx15x, A2 => n7509, ZN => 
                           IF_RegsxN675);
   U3949 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx31x, A2 => n7523, ZN => 
                           IF_RegsxN691);
   U3950 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx24x, A2 => n7523, ZN => 
                           IF_RegsxN684);
   U3951 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx16x, A2 => n7523, ZN => 
                           IF_RegsxN676);
   U3952 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx30x, A2 => n7523, ZN => 
                           IF_RegsxN690);
   U3953 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx29x, A2 => n7523, ZN => 
                           IF_RegsxN689);
   U3954 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx3x, A2 => n7523, ZN => 
                           IF_RegsxN663);
   U3955 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx2x, A2 => n7509, ZN => 
                           IF_RegsxN662);
   U3956 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx7x, A2 => n7523, ZN => 
                           IF_RegsxN667);
   U3957 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx1x, A2 => n7509, ZN => 
                           IF_RegsxN661);
   U3958 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx9x, A2 => n7520, ZN => 
                           IF_RegsxN669);
   U3959 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx5x, A2 => n7523, ZN => 
                           IF_RegsxN665);
   U3960 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx21x, A2 => n7509, ZN => 
                           IF_RegsxN681);
   U3961 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx0x, A2 => n7509, ZN => 
                           IF_RegsxN660);
   U3962 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx17x, A2 => n7509, ZN => 
                           IF_RegsxN677);
   U3963 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx4x, A2 => n7509, ZN => 
                           IF_RegsxN664);
   U3964 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx14x, A2 => n7523, ZN => 
                           IF_RegsxN674);
   U3965 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx13x, A2 => n7509, ZN => 
                           IF_RegsxN673);
   U3966 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx19x, A2 => n7509, ZN => 
                           IF_RegsxN679);
   U3967 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx18x, A2 => n7523, ZN => 
                           IF_RegsxN678);
   U3968 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx6x, A2 => n7509, ZN => 
                           IF_RegsxN666);
   U3969 : AND2_X1 port map( A1 => toRegsPortxDSTDATAxx25x, A2 => n7509, ZN => 
                           IF_RegsxN685);
   U3970 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(26), A2 => n4944,
                           ZN => add_x_26xBx6x);
   U3971 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(16), A2 => 
                           fromMemoryPortxLOADEDDATAx(15), ZN => n3652);
   U3972 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(17), ZN => n6839);
   U3973 : NAND2_X1 port map( A1 => n3652, A2 => n6839, ZN => n3665);
   U3974 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(18), ZN => n6877);
   U3975 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(19), A2 => n6877
                           , ZN => n3658);
   U3976 : NOR2_X1 port map( A1 => n3665, A2 => n3658, ZN => n3959);
   U3977 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(15), ZN => n6759);
   U3978 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(16), A2 => n6839
                           , A3 => n6759, ZN => n3671);
   U3979 : NOR2_X1 port map( A1 => n3658, A2 => n3671, ZN => n5166);
   U3980 : AOI22_X1 port map( A1 => n3959, A2 => fromRegsPortxREG_FILE_16xx12x,
                           B1 => n5166, B2 => fromRegsPortxREG_FILE_18xx12x, ZN
                           => n3651);
   U3981 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(18), A2 => 
                           fromMemoryPortxLOADEDDATAx(19), ZN => n3672);
   U3982 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(17), A2 => 
                           fromMemoryPortxLOADEDDATAx(16), A3 => 
                           fromMemoryPortxLOADEDDATAx(15), ZN => n3668);
   U3983 : NOR2_X1 port map( A1 => n3672, A2 => n3668, ZN => n5158);
   U3984 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(19), ZN => n6916);
   U3985 : NAND2_X1 port map( A1 => n6877, A2 => n6916, ZN => n3669);
   U3986 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(16), A2 => 
                           fromMemoryPortxLOADEDDATAx(15), A3 => n6839, ZN => 
                           n3670);
   U3987 : NOR2_X1 port map( A1 => n3669, A2 => n3670, ZN => n5176);
   U3988 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_31xx12x,
                           B1 => n5176, B2 => fromRegsPortxREG_FILE_03xx12x, ZN
                           => n3650);
   U3989 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(16), A2 => 
                           fromMemoryPortxLOADEDDATAx(17), A3 => n6759, ZN => 
                           n3667);
   U3990 : NOR2_X1 port map( A1 => n3669, A2 => n3667, ZN => n5197);
   U3991 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(18), A2 => n6916
                           , ZN => n3659);
   U3992 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(16), ZN => n6800);
   U3993 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(17), A2 => 
                           fromMemoryPortxLOADEDDATAx(15), A3 => n6800, ZN => 
                           n3664);
   U3994 : NOR2_X1 port map( A1 => n3659, A2 => n3664, ZN => n5246);
   U3995 : AOI22_X1 port map( A1 => n5197, A2 => fromRegsPortxREG_FILE_06xx12x,
                           B1 => n5246, B2 => fromRegsPortxREG_FILE_13xx12x, ZN
                           => n3649);
   U3996 : NOR2_X1 port map( A1 => n3658, A2 => n3668, ZN => n5211);
   U3997 : NOR2_X1 port map( A1 => n3659, A2 => n3671, ZN => n5167);
   U3998 : AOI22_X1 port map( A1 => n5211, A2 => fromRegsPortxREG_FILE_23xx12x,
                           B1 => n5167, B2 => fromRegsPortxREG_FILE_10xx12x, ZN
                           => n3648);
   U3999 : AND4_X1 port map( A1 => n3651, A2 => n3650, A3 => n3649, A4 => n3648
                           , ZN => n3680);
   U4000 : NOR2_X1 port map( A1 => n3659, A2 => n3668, ZN => n5160);
   U4001 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(17), A2 => n3652
                           , ZN => n3657);
   U4002 : NOR2_X1 port map( A1 => n3659, A2 => n3657, ZN => n5202);
   U4003 : AOI22_X1 port map( A1 => n5160, A2 => fromRegsPortxREG_FILE_15xx12x,
                           B1 => n5202, B2 => fromRegsPortxREG_FILE_12xx12x, ZN
                           => n3656);
   U4004 : NOR2_X1 port map( A1 => n3672, A2 => n3664, ZN => n5153);
   U4005 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(15), A2 => n6839
                           , A3 => n6800, ZN => n3666);
   U4006 : NOR2_X1 port map( A1 => n3666, A2 => n3658, ZN => n5251);
   U4007 : AOI22_X1 port map( A1 => n5153, A2 => fromRegsPortxREG_FILE_29xx12x,
                           B1 => n5251, B2 => fromRegsPortxREG_FILE_17xx12x, ZN
                           => n3655);
   U4008 : NOR2_X1 port map( A1 => n3659, A2 => n3665, ZN => n5147);
   U4009 : NOR2_X1 port map( A1 => n3672, A2 => n3657, ZN => n5159);
   U4010 : AOI22_X1 port map( A1 => n5147, A2 => fromRegsPortxREG_FILE_08xx12x,
                           B1 => n5159, B2 => fromRegsPortxREG_FILE_28xx12x, ZN
                           => n3654);
   U4011 : NOR2_X1 port map( A1 => n3666, A2 => n3672, ZN => n5267);
   U4012 : NOR2_X1 port map( A1 => n3669, A2 => n3657, ZN => n5252);
   U4013 : CLKBUF_X1 port map( A => n5252, Z => n5357);
   U4014 : AOI22_X1 port map( A1 => n5267, A2 => fromRegsPortxREG_FILE_25xx12x,
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx12x, ZN
                           => n3653);
   U4015 : AND4_X1 port map( A1 => n3656, A2 => n3655, A3 => n3654, A4 => n3653
                           , ZN => n3679);
   U4016 : NOR2_X1 port map( A1 => n3659, A2 => n3670, ZN => n5258);
   U4017 : CLKBUF_X1 port map( A => n5258, Z => n5341);
   U4018 : NOR2_X1 port map( A1 => n3659, A2 => n3666, ZN => n5235);
   U4019 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_11xx12x,
                           B1 => n5235, B2 => fromRegsPortxREG_FILE_09xx12x, ZN
                           => n3663);
   U4020 : NOR2_X1 port map( A1 => n3658, A2 => n3657, ZN => n5165);
   U4021 : NOR2_X1 port map( A1 => n3667, A2 => n3658, ZN => n5225);
   U4022 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_20xx12x,
                           B1 => n5225, B2 => fromRegsPortxREG_FILE_22xx12x, ZN
                           => n3662);
   U4023 : NOR2_X1 port map( A1 => n3669, A2 => n3671, ZN => n5260);
   U4024 : NOR2_X1 port map( A1 => n3664, A2 => n3658, ZN => n5342);
   U4025 : AOI22_X1 port map( A1 => n5260, A2 => fromRegsPortxREG_FILE_02xx12x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_21xx12x, ZN
                           => n3661);
   U4026 : NOR2_X1 port map( A1 => n3658, A2 => n3670, ZN => n5244);
   U4027 : CLKBUF_X1 port map( A => n5244, Z => n5367);
   U4028 : NOR2_X1 port map( A1 => n3659, A2 => n3667, ZN => n5152);
   U4029 : AOI22_X1 port map( A1 => n5367, A2 => fromRegsPortxREG_FILE_19xx12x,
                           B1 => n5152, B2 => fromRegsPortxREG_FILE_14xx12x, ZN
                           => n3660);
   U4030 : AND4_X1 port map( A1 => n3663, A2 => n3662, A3 => n3661, A4 => n3660
                           , ZN => n3678);
   U4031 : NOR2_X1 port map( A1 => n3669, A2 => n3664, ZN => n5220);
   U4032 : NOR2_X1 port map( A1 => n3665, A2 => n3672, ZN => n5266);
   U4033 : AOI22_X1 port map( A1 => n5220, A2 => fromRegsPortxREG_FILE_05xx12x,
                           B1 => n5266, B2 => fromRegsPortxREG_FILE_24xx12x, ZN
                           => n3676);
   U4034 : NOR2_X1 port map( A1 => n3666, A2 => n3669, ZN => n5253);
   U4035 : CLKBUF_X1 port map( A => n5253, Z => n5380);
   U4036 : NOR2_X1 port map( A1 => n3672, A2 => n3667, ZN => n5268);
   U4037 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx12x,
                           B1 => n5268, B2 => fromRegsPortxREG_FILE_30xx12x, ZN
                           => n3675);
   U4038 : NOR2_X1 port map( A1 => n3669, A2 => n3668, ZN => n5230);
   U4039 : CLKBUF_X1 port map( A => n5230, Z => n5343);
   U4040 : NAND2_X1 port map( A1 => n5343, A2 => fromRegsPortxREG_FILE_07xx12x,
                           ZN => n3674);
   U4041 : NOR2_X1 port map( A1 => n3672, A2 => n3670, ZN => n5261);
   U4042 : NOR2_X1 port map( A1 => n3672, A2 => n3671, ZN => n5245);
   U4043 : AOI22_X1 port map( A1 => n5261, A2 => fromRegsPortxREG_FILE_27xx12x,
                           B1 => n5245, B2 => fromRegsPortxREG_FILE_26xx12x, ZN
                           => n3673);
   U4044 : AND4_X1 port map( A1 => n3676, A2 => n3675, A3 => n3674, A4 => n3673
                           , ZN => n3677);
   U4045 : NAND4_X1 port map( A1 => n3680, A2 => n3679, A3 => n3678, A4 => 
                           n3677, ZN => ashr_25xAx12x);
   U4046 : INV_X1 port map( A => ashr_25xAx12x, ZN => intadd_27xAx1x);
   U4047 : CLKBUF_X1 port map( A => n5220, Z => n5374);
   U4048 : CLKBUF_X1 port map( A => n5167, Z => n5369);
   U4049 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx2x, 
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx2x, ZN 
                           => n3684);
   U4050 : CLKBUF_X1 port map( A => n5165, Z => n5354);
   U4051 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx2x, 
                           B1 => n5244, B2 => fromRegsPortxREG_FILE_19xx2x, ZN 
                           => n3683);
   U4052 : CLKBUF_X1 port map( A => n5235, Z => n5340);
   U4053 : AOI22_X1 port map( A1 => n3959, A2 => fromRegsPortxREG_FILE_16xx2x, 
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx2x, ZN 
                           => n3682);
   U4054 : CLKBUF_X1 port map( A => n5147, Z => n5378);
   U4055 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx2x, 
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_01xx2x, ZN 
                           => n3681);
   U4056 : AND4_X1 port map( A1 => n3684, A2 => n3683, A3 => n3682, A4 => n3681
                           , ZN => n3700);
   U4057 : CLKBUF_X1 port map( A => n5159, Z => n5377);
   U4058 : CLKBUF_X1 port map( A => n5342, Z => n5259);
   U4059 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_28xx2x, 
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx2x, ZN 
                           => n3688);
   U4060 : CLKBUF_X1 port map( A => n5197, Z => n5362);
   U4061 : CLKBUF_X1 port map( A => n5202, Z => n5356);
   U4062 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx2x, 
                           B1 => n5356, B2 => fromRegsPortxREG_FILE_12xx2x, ZN 
                           => n3687);
   U4063 : CLKBUF_X1 port map( A => n5225, Z => n5352);
   U4064 : AOI22_X1 port map( A1 => n5260, A2 => fromRegsPortxREG_FILE_02xx2x, 
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx2x, ZN 
                           => n3686);
   U4065 : CLKBUF_X1 port map( A => n5211, Z => n5338);
   U4066 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx2x, 
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_11xx2x, ZN 
                           => n3685);
   U4067 : AND4_X1 port map( A1 => n3688, A2 => n3687, A3 => n3686, A4 => n3685
                           , ZN => n3699);
   U4068 : CLKBUF_X1 port map( A => n5153, Z => n5351);
   U4069 : CLKBUF_X1 port map( A => n5166, Z => n5364);
   U4070 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx2x, 
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx2x, ZN 
                           => n3692);
   U4071 : CLKBUF_X1 port map( A => n5176, Z => n5355);
   U4072 : CLKBUF_X1 port map( A => n5152, Z => n5368);
   U4073 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx2x, 
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx2x, ZN 
                           => n3691);
   U4074 : CLKBUF_X1 port map( A => n5268, Z => n5339);
   U4075 : CLKBUF_X1 port map( A => n5246, Z => n5366);
   U4076 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx2x, 
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx2x, ZN 
                           => n3690);
   U4077 : CLKBUF_X1 port map( A => n5160, Z => n5344);
   U4078 : CLKBUF_X1 port map( A => n5266, Z => n5376);
   U4079 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx2x, 
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_24xx2x, ZN 
                           => n3689);
   U4080 : AND4_X1 port map( A1 => n3692, A2 => n3691, A3 => n3690, A4 => n3689
                           , ZN => n3698);
   U4081 : CLKBUF_X1 port map( A => n5251, Z => n5350);
   U4082 : CLKBUF_X1 port map( A => n5158, Z => n5379);
   U4083 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx2x, 
                           B1 => n5379, B2 => fromRegsPortxREG_FILE_31xx2x, ZN 
                           => n3696);
   U4084 : CLKBUF_X1 port map( A => n5261, Z => n5353);
   U4085 : AOI22_X1 port map( A1 => n5343, A2 => fromRegsPortxREG_FILE_07xx2x, 
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx2x, ZN 
                           => n3695);
   U4086 : CLKBUF_X1 port map( A => n5267, Z => n5363);
   U4087 : CLKBUF_X1 port map( A => n5245, Z => n5365);
   U4088 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx2x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx2x, ZN 
                           => n3694);
   U4089 : NAND2_X1 port map( A1 => n5357, A2 => fromRegsPortxREG_FILE_04xx2x, 
                           ZN => n3693);
   U4090 : AND4_X1 port map( A1 => n3696, A2 => n3695, A3 => n3694, A4 => n3693
                           , ZN => n3697);
   U4091 : NAND4_X1 port map( A1 => n3700, A2 => n3699, A3 => n3698, A4 => 
                           n3697, ZN => ashr_25xAx2x);
   U4092 : INV_X1 port map( A => ashr_25xAx2x, ZN => intadd_29xAx1x);
   U4093 : AOI22_X1 port map( A1 => n5356, A2 => fromRegsPortxREG_FILE_12xx3x, 
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx3x, ZN 
                           => n3704);
   U4094 : CLKBUF_X1 port map( A => n5260, Z => n5375);
   U4095 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx3x, 
                           B1 => n5375, B2 => fromRegsPortxREG_FILE_02xx3x, ZN 
                           => n3703);
   U4096 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx3x, 
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx3x, ZN 
                           => n3702);
   U4097 : AOI22_X1 port map( A1 => n5367, A2 => fromRegsPortxREG_FILE_19xx3x, 
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx3x, ZN 
                           => n3701);
   U4098 : AND4_X1 port map( A1 => n3704, A2 => n3703, A3 => n3702, A4 => n3701
                           , ZN => n3722);
   U4099 : AOI22_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_27xx3x, 
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx3x, ZN 
                           => n3706);
   U4100 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx3x, 
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx3x, ZN 
                           => n3705);
   U4101 : NAND2_X1 port map( A1 => n3706, A2 => n3705, ZN => n3711);
   U4102 : AOI22_X1 port map( A1 => n3959, A2 => fromRegsPortxREG_FILE_16xx3x, 
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx3x, ZN 
                           => n3709);
   U4103 : NAND2_X1 port map( A1 => n5343, A2 => fromRegsPortxREG_FILE_07xx3x, 
                           ZN => n3708);
   U4104 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx3x, 
                           B1 => n5379, B2 => fromRegsPortxREG_FILE_31xx3x, ZN 
                           => n3707);
   U4105 : NAND3_X1 port map( A1 => n3709, A2 => n3708, A3 => n3707, ZN => 
                           n3710);
   U4106 : NOR2_X1 port map( A1 => n3711, A2 => n3710, ZN => n3721);
   U4107 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx3x, 
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx3x, ZN 
                           => n3715);
   U4108 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx3x, 
                           B1 => n5167, B2 => fromRegsPortxREG_FILE_10xx3x, ZN 
                           => n3714);
   U4109 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx3x, 
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_01xx3x, ZN 
                           => n3713);
   U4110 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx3x, 
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_11xx3x, ZN 
                           => n3712);
   U4111 : AND4_X1 port map( A1 => n3715, A2 => n3714, A3 => n3713, A4 => n3712
                           , ZN => n3720);
   U4112 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_20xx3x, 
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_28xx3x, ZN 
                           => n3718);
   U4113 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx3x, 
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_05xx3x, ZN 
                           => n3717);
   U4114 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_24xx3x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx3x, ZN 
                           => n3716);
   U4115 : AND3_X1 port map( A1 => n3718, A2 => n3717, A3 => n3716, ZN => n3719
                           );
   U4116 : NAND4_X1 port map( A1 => n3722, A2 => n3721, A3 => n3720, A4 => 
                           n3719, ZN => ashr_25xAx3x);
   U4117 : INV_X1 port map( A => ashr_25xAx3x, ZN => intadd_29xAx2x);
   U4118 : CLKBUF_X1 port map( A => n6456, Z => n6811);
   U4119 : INV_X2 port map( A => n6811, ZN => intadd_29xBx1x);
   U4120 : INV_X1 port map( A => ashr_25xSHx3x, ZN => n7236);
   U4121 : CLKBUF_X2 port map( A => n7236, Z => intadd_29xBx2x);
   U4122 : CLKBUF_X2 port map( A => n5680, Z => n7551);
   U4123 : NAND2_X1 port map( A1 => n7446, A2 => fromMemoryPortxLOADEDDATAx(11)
                           , ZN => n3725);
   U4124 : NAND2_X1 port map( A1 => n3723, A2 => fromMemoryPortxLOADEDDATAx(24)
                           , ZN => n3724);
   U4125 : NAND2_X1 port map( A1 => n3725, A2 => n3724, ZN => ashr_25xSHx4x);
   U4126 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_28xx26x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx26x, ZN
                           => n3729);
   U4127 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx26x,
                           B1 => n5351, B2 => fromRegsPortxREG_FILE_29xx26x, ZN
                           => n3728);
   U4128 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx26x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx26x, ZN
                           => n3727);
   U4129 : NAND2_X1 port map( A1 => n5357, A2 => fromRegsPortxREG_FILE_04xx26x,
                           ZN => n3726);
   U4130 : AND4_X1 port map( A1 => n3729, A2 => n3728, A3 => n3727, A4 => n3726
                           , ZN => n3745);
   U4131 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_24xx26x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_21xx26x, ZN
                           => n3733);
   U4132 : AOI22_X1 port map( A1 => n5340, A2 => fromRegsPortxREG_FILE_09xx26x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx26x, ZN
                           => n3732);
   U4133 : CLKBUF_X1 port map( A => n3959, Z => n5345);
   U4134 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx26x,
                           B1 => n5345, B2 => fromRegsPortxREG_FILE_16xx26x, ZN
                           => n3731);
   U4135 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx26x,
                           B1 => n5356, B2 => fromRegsPortxREG_FILE_12xx26x, ZN
                           => n3730);
   U4136 : AND4_X1 port map( A1 => n3733, A2 => n3732, A3 => n3731, A4 => n3730
                           , ZN => n3744);
   U4137 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx26x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx26x, ZN
                           => n3737);
   U4138 : AOI22_X1 port map( A1 => n5367, A2 => fromRegsPortxREG_FILE_19xx26x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx26x, ZN
                           => n3736);
   U4139 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx26x,
                           B1 => n5341, B2 => fromRegsPortxREG_FILE_11xx26x, ZN
                           => n3735);
   U4140 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx26x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx26x, ZN
                           => n3734);
   U4141 : AND4_X1 port map( A1 => n3737, A2 => n3736, A3 => n3735, A4 => n3734
                           , ZN => n3743);
   U4142 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx26x,
                           B1 => n5375, B2 => fromRegsPortxREG_FILE_02xx26x, ZN
                           => n3741);
   U4143 : AOI22_X1 port map( A1 => n5379, A2 => fromRegsPortxREG_FILE_31xx26x,
                           B1 => n5355, B2 => fromRegsPortxREG_FILE_03xx26x, ZN
                           => n3740);
   U4144 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx26x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx26x, ZN
                           => n3739);
   U4145 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx26x,
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx26x, ZN
                           => n3738);
   U4146 : AND4_X1 port map( A1 => n3741, A2 => n3740, A3 => n3739, A4 => n3738
                           , ZN => n3742);
   U4147 : NAND4_X1 port map( A1 => n3745, A2 => n3744, A3 => n3743, A4 => 
                           n3742, ZN => ashr_25xAx26x);
   U4148 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_31xx11x,
                           B1 => n5176, B2 => fromRegsPortxREG_FILE_03xx11x, ZN
                           => n3749);
   U4149 : AOI22_X1 port map( A1 => n5268, A2 => fromRegsPortxREG_FILE_30xx11x,
                           B1 => n5166, B2 => fromRegsPortxREG_FILE_18xx11x, ZN
                           => n3748);
   U4150 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx11x,
                           B1 => n5167, B2 => fromRegsPortxREG_FILE_10xx11x, ZN
                           => n3747);
   U4151 : AOI22_X1 port map( A1 => n5153, A2 => fromRegsPortxREG_FILE_29xx11x,
                           B1 => n5244, B2 => fromRegsPortxREG_FILE_19xx11x, ZN
                           => n3746);
   U4152 : AND4_X1 port map( A1 => n3749, A2 => n3748, A3 => n3747, A4 => n3746
                           , ZN => n3765);
   U4153 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_20xx11x,
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx11x, ZN
                           => n3753);
   U4154 : AOI22_X1 port map( A1 => n5260, A2 => fromRegsPortxREG_FILE_02xx11x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx11x, ZN
                           => n3752);
   U4155 : AOI22_X1 port map( A1 => n5147, A2 => fromRegsPortxREG_FILE_08xx11x,
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx11x, ZN
                           => n3751);
   U4156 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx11x,
                           B1 => n5251, B2 => fromRegsPortxREG_FILE_17xx11x, ZN
                           => n3750);
   U4157 : AND4_X1 port map( A1 => n3753, A2 => n3752, A3 => n3751, A4 => n3750
                           , ZN => n3764);
   U4158 : AOI22_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_01xx11x,
                           B1 => n5211, B2 => fromRegsPortxREG_FILE_23xx11x, ZN
                           => n3757);
   U4159 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_11xx11x,
                           B1 => n5152, B2 => fromRegsPortxREG_FILE_14xx11x, ZN
                           => n3756);
   U4160 : AOI22_X1 port map( A1 => n3959, A2 => fromRegsPortxREG_FILE_16xx11x,
                           B1 => n5160, B2 => fromRegsPortxREG_FILE_15xx11x, ZN
                           => n3755);
   U4161 : AOI22_X1 port map( A1 => n5230, A2 => fromRegsPortxREG_FILE_07xx11x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx11x, ZN
                           => n3754);
   U4162 : AND4_X1 port map( A1 => n3757, A2 => n3756, A3 => n3755, A4 => n3754
                           , ZN => n3763);
   U4163 : AOI22_X1 port map( A1 => n5159, A2 => fromRegsPortxREG_FILE_28xx11x,
                           B1 => n5266, B2 => fromRegsPortxREG_FILE_24xx11x, ZN
                           => n3761);
   U4164 : AOI22_X1 port map( A1 => n5356, A2 => fromRegsPortxREG_FILE_12xx11x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx11x, ZN
                           => n3760);
   U4165 : AOI22_X1 port map( A1 => n5197, A2 => fromRegsPortxREG_FILE_06xx11x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx11x, ZN
                           => n3759);
   U4166 : NAND2_X1 port map( A1 => n5246, A2 => fromRegsPortxREG_FILE_13xx11x,
                           ZN => n3758);
   U4167 : AND4_X1 port map( A1 => n3761, A2 => n3760, A3 => n3759, A4 => n3758
                           , ZN => n3762);
   U4168 : NAND4_X1 port map( A1 => n3765, A2 => n3764, A3 => n3763, A4 => 
                           n3762, ZN => ashr_25xAx11x);
   U4169 : INV_X1 port map( A => ashr_25xAx11x, ZN => intadd_27xAx0x);
   U4170 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx0x, 
                           B1 => n5354, B2 => fromRegsPortxREG_FILE_20xx0x, ZN 
                           => n3768);
   U4171 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx0x, 
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx0x, ZN 
                           => n3767);
   U4172 : AOI22_X1 port map( A1 => n5367, A2 => fromRegsPortxREG_FILE_19xx0x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx0x, ZN 
                           => n3766);
   U4173 : AND3_X1 port map( A1 => n3768, A2 => n3767, A3 => n3766, ZN => n3787
                           );
   U4174 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx0x, 
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_28xx0x, ZN 
                           => n3770);
   U4175 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx0x, 
                           B1 => n5345, B2 => fromRegsPortxREG_FILE_16xx0x, ZN 
                           => n3769);
   U4176 : NAND2_X1 port map( A1 => n3770, A2 => n3769, ZN => n3775);
   U4177 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_24xx0x, 
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx0x, ZN 
                           => n3773);
   U4178 : NAND2_X1 port map( A1 => n5357, A2 => fromRegsPortxREG_FILE_04xx0x, 
                           ZN => n3772);
   U4179 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx0x, 
                           B1 => n5379, B2 => fromRegsPortxREG_FILE_31xx0x, ZN 
                           => n3771);
   U4180 : NAND3_X1 port map( A1 => n3773, A2 => n3772, A3 => n3771, ZN => 
                           n3774);
   U4181 : NOR2_X1 port map( A1 => n3775, A2 => n3774, ZN => n3786);
   U4182 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx0x, 
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx0x, ZN 
                           => n3779);
   U4183 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_11xx0x, 
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx0x, ZN 
                           => n3778);
   U4184 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx0x, 
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx0x, ZN 
                           => n3777);
   U4185 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx0x, 
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx0x, ZN 
                           => n3776);
   U4186 : AND4_X1 port map( A1 => n3779, A2 => n3778, A3 => n3777, A4 => n3776
                           , ZN => n3785);
   U4187 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx0x, 
                           B1 => n5375, B2 => fromRegsPortxREG_FILE_02xx0x, ZN 
                           => n3783);
   U4188 : AOI22_X1 port map( A1 => n5356, A2 => fromRegsPortxREG_FILE_12xx0x, 
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx0x, ZN 
                           => n3782);
   U4189 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx0x, 
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx0x, ZN 
                           => n3781);
   U4190 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx0x, 
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx0x, ZN 
                           => n3780);
   U4191 : AND4_X1 port map( A1 => n3783, A2 => n3782, A3 => n3781, A4 => n3780
                           , ZN => n3784);
   U4192 : NAND4_X1 port map( A1 => n3787, A2 => n3786, A3 => n3785, A4 => 
                           n3784, ZN => ashr_25xAx0x);
   U4193 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx1x, 
                           B1 => n5379, B2 => fromRegsPortxREG_FILE_31xx1x, ZN 
                           => n3791);
   U4194 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx1x, 
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx1x, ZN 
                           => n3790);
   U4195 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_24xx1x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx1x, ZN 
                           => n3789);
   U4196 : NAND2_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_28xx1x, 
                           ZN => n3788);
   U4197 : AND4_X1 port map( A1 => n3791, A2 => n3790, A3 => n3789, A4 => n3788
                           , ZN => n3807);
   U4198 : AOI22_X1 port map( A1 => n5340, A2 => fromRegsPortxREG_FILE_09xx1x, 
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx1x, ZN 
                           => n3795);
   U4199 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx1x, 
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx1x, ZN 
                           => n3794);
   U4200 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx1x, 
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_23xx1x, ZN 
                           => n3793);
   U4201 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx1x, 
                           B1 => n5341, B2 => fromRegsPortxREG_FILE_11xx1x, ZN 
                           => n3792);
   U4202 : AND4_X1 port map( A1 => n3795, A2 => n3794, A3 => n3793, A4 => n3792
                           , ZN => n3806);
   U4203 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx1x, 
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx1x, ZN 
                           => n3799);
   U4204 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx1x, 
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx1x, ZN 
                           => n3798);
   U4205 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_02xx1x, 
                           B1 => n5252, B2 => fromRegsPortxREG_FILE_04xx1x, ZN 
                           => n3797);
   U4206 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx1x, 
                           B1 => n5344, B2 => fromRegsPortxREG_FILE_15xx1x, ZN 
                           => n3796);
   U4207 : AND4_X1 port map( A1 => n3799, A2 => n3798, A3 => n3797, A4 => n3796
                           , ZN => n3805);
   U4208 : AOI22_X1 port map( A1 => n5356, A2 => fromRegsPortxREG_FILE_12xx1x, 
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx1x, ZN 
                           => n3803);
   U4209 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx1x, 
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx1x, ZN 
                           => n3802);
   U4210 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx1x, 
                           B1 => n5367, B2 => fromRegsPortxREG_FILE_19xx1x, ZN 
                           => n3801);
   U4211 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx1x, 
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx1x, ZN 
                           => n3800);
   U4212 : AND4_X1 port map( A1 => n3803, A2 => n3802, A3 => n3801, A4 => n3800
                           , ZN => n3804);
   U4213 : NAND4_X1 port map( A1 => n3807, A2 => n3806, A3 => n3805, A4 => 
                           n3804, ZN => ashr_25xAx1x);
   U4214 : AOI22_X1 port map( A1 => n5379, A2 => fromRegsPortxREG_FILE_31xx4x, 
                           B1 => n5220, B2 => fromRegsPortxREG_FILE_05xx4x, ZN 
                           => n3811);
   U4215 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx4x, 
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_06xx4x, ZN 
                           => n3810);
   U4216 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_22xx4x, 
                           B1 => n5244, B2 => fromRegsPortxREG_FILE_19xx4x, ZN 
                           => n3809);
   U4217 : AOI22_X1 port map( A1 => n5261, A2 => fromRegsPortxREG_FILE_27xx4x, 
                           B1 => n5166, B2 => fromRegsPortxREG_FILE_18xx4x, ZN 
                           => n3808);
   U4218 : AND4_X1 port map( A1 => n3811, A2 => n3810, A3 => n3809, A4 => n3808
                           , ZN => n3827);
   U4219 : AOI22_X1 port map( A1 => n5235, A2 => fromRegsPortxREG_FILE_09xx4x, 
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx4x, ZN 
                           => n3815);
   U4220 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx4x, 
                           B1 => n5202, B2 => fromRegsPortxREG_FILE_12xx4x, ZN 
                           => n3814);
   U4221 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx4x, 
                           B1 => n5165, B2 => fromRegsPortxREG_FILE_20xx4x, ZN 
                           => n3813);
   U4222 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx4x, 
                           B1 => n5159, B2 => fromRegsPortxREG_FILE_28xx4x, ZN 
                           => n3812);
   U4223 : AND4_X1 port map( A1 => n3815, A2 => n3814, A3 => n3813, A4 => n3812
                           , ZN => n3826);
   U4224 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_11xx4x, 
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx4x, ZN 
                           => n3819);
   U4225 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx4x, 
                           B1 => n5167, B2 => fromRegsPortxREG_FILE_10xx4x, ZN 
                           => n3818);
   U4226 : AOI22_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_01xx4x, 
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx4x, ZN 
                           => n3817);
   U4227 : AOI22_X1 port map( A1 => n3959, A2 => fromRegsPortxREG_FILE_16xx4x, 
                           B1 => n5160, B2 => fromRegsPortxREG_FILE_15xx4x, ZN 
                           => n3816);
   U4228 : AND4_X1 port map( A1 => n3819, A2 => n3818, A3 => n3817, A4 => n3816
                           , ZN => n3825);
   U4229 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_24xx4x, 
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx4x, ZN 
                           => n3823);
   U4230 : NAND2_X1 port map( A1 => n5260, A2 => fromRegsPortxREG_FILE_02xx4x, 
                           ZN => n3822);
   U4231 : AOI22_X1 port map( A1 => n5366, A2 => fromRegsPortxREG_FILE_13xx4x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx4x, ZN 
                           => n3821);
   U4232 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx4x, 
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_30xx4x, ZN 
                           => n3820);
   U4233 : AND4_X1 port map( A1 => n3823, A2 => n3822, A3 => n3821, A4 => n3820
                           , ZN => n3824);
   U4234 : NAND4_X1 port map( A1 => n3827, A2 => n3826, A3 => n3825, A4 => 
                           n3824, ZN => ashr_25xAx4x);
   U4235 : AOI22_X1 port map( A1 => n5252, A2 => fromRegsPortxREG_FILE_04xx5x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx5x, ZN 
                           => n3831);
   U4236 : AOI22_X1 port map( A1 => n5153, A2 => fromRegsPortxREG_FILE_29xx5x, 
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx5x, ZN 
                           => n3830);
   U4237 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx5x, 
                           B1 => n5268, B2 => fromRegsPortxREG_FILE_30xx5x, ZN 
                           => n3829);
   U4238 : NAND2_X1 port map( A1 => n5266, A2 => fromRegsPortxREG_FILE_24xx5x, 
                           ZN => n3828);
   U4239 : AND4_X1 port map( A1 => n3831, A2 => n3830, A3 => n3829, A4 => n3828
                           , ZN => n3847);
   U4240 : AOI22_X1 port map( A1 => n5197, A2 => fromRegsPortxREG_FILE_06xx5x, 
                           B1 => n5345, B2 => fromRegsPortxREG_FILE_16xx5x, ZN 
                           => n3835);
   U4241 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_31xx5x, 
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx5x, ZN 
                           => n3834);
   U4242 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx5x, 
                           B1 => n5159, B2 => fromRegsPortxREG_FILE_28xx5x, ZN 
                           => n3833);
   U4243 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx5x, 
                           B1 => n5202, B2 => fromRegsPortxREG_FILE_12xx5x, ZN 
                           => n3832);
   U4244 : AND4_X1 port map( A1 => n3835, A2 => n3834, A3 => n3833, A4 => n3832
                           , ZN => n3846);
   U4245 : AOI22_X1 port map( A1 => n5367, A2 => fromRegsPortxREG_FILE_19xx5x, 
                           B1 => n5167, B2 => fromRegsPortxREG_FILE_10xx5x, ZN 
                           => n3839);
   U4246 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_20xx5x, 
                           B1 => n5152, B2 => fromRegsPortxREG_FILE_14xx5x, ZN 
                           => n3838);
   U4247 : AOI22_X1 port map( A1 => n5225, A2 => fromRegsPortxREG_FILE_22xx5x, 
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx5x, ZN 
                           => n3837);
   U4248 : AOI22_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_01xx5x, 
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_11xx5x, ZN 
                           => n3836);
   U4249 : AND4_X1 port map( A1 => n3839, A2 => n3838, A3 => n3837, A4 => n3836
                           , ZN => n3845);
   U4250 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx5x, 
                           B1 => n5375, B2 => fromRegsPortxREG_FILE_02xx5x, ZN 
                           => n3843);
   U4251 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx5x, 
                           B1 => n5220, B2 => fromRegsPortxREG_FILE_05xx5x, ZN 
                           => n3842);
   U4252 : AOI22_X1 port map( A1 => n5235, A2 => fromRegsPortxREG_FILE_09xx5x, 
                           B1 => n5166, B2 => fromRegsPortxREG_FILE_18xx5x, ZN 
                           => n3841);
   U4253 : AOI22_X1 port map( A1 => n5147, A2 => fromRegsPortxREG_FILE_08xx5x, 
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx5x, ZN 
                           => n3840);
   U4254 : AND4_X1 port map( A1 => n3843, A2 => n3842, A3 => n3841, A4 => n3840
                           , ZN => n3844);
   U4255 : NAND4_X1 port map( A1 => n3847, A2 => n3846, A3 => n3845, A4 => 
                           n3844, ZN => ashr_25xAx5x);
   U4256 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_28xx6x, 
                           B1 => n5244, B2 => fromRegsPortxREG_FILE_19xx6x, ZN 
                           => n3851);
   U4257 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx6x, 
                           B1 => n5166, B2 => fromRegsPortxREG_FILE_18xx6x, ZN 
                           => n3850);
   U4258 : AOI22_X1 port map( A1 => n5365, A2 => fromRegsPortxREG_FILE_26xx6x, 
                           B1 => n5167, B2 => fromRegsPortxREG_FILE_10xx6x, ZN 
                           => n3849);
   U4259 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx6x, 
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx6x, ZN 
                           => n3848);
   U4260 : AND4_X1 port map( A1 => n3851, A2 => n3850, A3 => n3849, A4 => n3848
                           , ZN => n3867);
   U4261 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx6x, 
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx6x, ZN 
                           => n3855);
   U4262 : AOI22_X1 port map( A1 => n5147, A2 => fromRegsPortxREG_FILE_08xx6x, 
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx6x, ZN 
                           => n3854);
   U4263 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx6x, 
                           B1 => n5354, B2 => fromRegsPortxREG_FILE_20xx6x, ZN 
                           => n3853);
   U4264 : AOI22_X1 port map( A1 => n5230, A2 => fromRegsPortxREG_FILE_07xx6x, 
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx6x, ZN 
                           => n3852);
   U4265 : AND4_X1 port map( A1 => n3855, A2 => n3854, A3 => n3853, A4 => n3852
                           , ZN => n3866);
   U4266 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx6x, 
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx6x, ZN 
                           => n3859);
   U4267 : AOI22_X1 port map( A1 => n5356, A2 => fromRegsPortxREG_FILE_12xx6x, 
                           B1 => n5152, B2 => fromRegsPortxREG_FILE_14xx6x, ZN 
                           => n3858);
   U4268 : AOI22_X1 port map( A1 => n3959, A2 => fromRegsPortxREG_FILE_16xx6x, 
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_01xx6x, ZN 
                           => n3857);
   U4269 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_24xx6x, 
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_11xx6x, ZN 
                           => n3856);
   U4270 : AND4_X1 port map( A1 => n3859, A2 => n3858, A3 => n3857, A4 => n3856
                           , ZN => n3865);
   U4271 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_31xx6x, 
                           B1 => n5220, B2 => fromRegsPortxREG_FILE_05xx6x, ZN 
                           => n3863);
   U4272 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx6x, 
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx6x, ZN 
                           => n3862);
   U4273 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx6x, 
                           B1 => n5268, B2 => fromRegsPortxREG_FILE_30xx6x, ZN 
                           => n3861);
   U4274 : NAND2_X1 port map( A1 => n5260, A2 => fromRegsPortxREG_FILE_02xx6x, 
                           ZN => n3860);
   U4275 : AND4_X1 port map( A1 => n3863, A2 => n3862, A3 => n3861, A4 => n3860
                           , ZN => n3864);
   U4276 : NAND4_X1 port map( A1 => n3867, A2 => n3866, A3 => n3865, A4 => 
                           n3864, ZN => ashr_25xAx6x);
   U4277 : AOI22_X1 port map( A1 => n5147, A2 => fromRegsPortxREG_FILE_08xx7x, 
                           B1 => n5176, B2 => fromRegsPortxREG_FILE_03xx7x, ZN 
                           => n3871);
   U4278 : AOI22_X1 port map( A1 => n5246, A2 => fromRegsPortxREG_FILE_13xx7x, 
                           B1 => n5166, B2 => fromRegsPortxREG_FILE_18xx7x, ZN 
                           => n3870);
   U4279 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_24xx7x, 
                           B1 => n5152, B2 => fromRegsPortxREG_FILE_14xx7x, ZN 
                           => n3869);
   U4280 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_22xx7x, 
                           B1 => n5167, B2 => fromRegsPortxREG_FILE_10xx7x, ZN 
                           => n3868);
   U4281 : AND4_X1 port map( A1 => n3871, A2 => n3870, A3 => n3869, A4 => n3868
                           , ZN => n3887);
   U4282 : AOI22_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_01xx7x, 
                           B1 => n5202, B2 => fromRegsPortxREG_FILE_12xx7x, ZN 
                           => n3875);
   U4283 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx7x, 
                           B1 => n5159, B2 => fromRegsPortxREG_FILE_28xx7x, ZN 
                           => n3874);
   U4284 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx7x, 
                           B1 => n5354, B2 => fromRegsPortxREG_FILE_20xx7x, ZN 
                           => n3873);
   U4285 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx7x, 
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx7x, ZN 
                           => n3872);
   U4286 : AND4_X1 port map( A1 => n3875, A2 => n3874, A3 => n3873, A4 => n3872
                           , ZN => n3886);
   U4287 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx7x, 
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_11xx7x, ZN 
                           => n3879);
   U4288 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_31xx7x, 
                           B1 => n5244, B2 => fromRegsPortxREG_FILE_19xx7x, ZN 
                           => n3878);
   U4289 : AOI22_X1 port map( A1 => n3959, A2 => fromRegsPortxREG_FILE_16xx7x, 
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx7x, ZN 
                           => n3877);
   U4290 : AOI22_X1 port map( A1 => n5153, A2 => fromRegsPortxREG_FILE_29xx7x, 
                           B1 => n5160, B2 => fromRegsPortxREG_FILE_15xx7x, ZN 
                           => n3876);
   U4291 : AND4_X1 port map( A1 => n3879, A2 => n3878, A3 => n3877, A4 => n3876
                           , ZN => n3885);
   U4292 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx7x, 
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx7x, ZN 
                           => n3883);
   U4293 : AOI22_X1 port map( A1 => n5260, A2 => fromRegsPortxREG_FILE_02xx7x, 
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx7x, ZN 
                           => n3882);
   U4294 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx7x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx7x, ZN 
                           => n3881);
   U4295 : NAND2_X1 port map( A1 => n5235, A2 => fromRegsPortxREG_FILE_09xx7x, 
                           ZN => n3880);
   U4296 : AND4_X1 port map( A1 => n3883, A2 => n3882, A3 => n3881, A4 => n3880
                           , ZN => n3884);
   U4297 : NAND4_X1 port map( A1 => n3887, A2 => n3886, A3 => n3885, A4 => 
                           n3884, ZN => ashr_25xAx7x);
   U4298 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx8x, 
                           B1 => n5176, B2 => fromRegsPortxREG_FILE_03xx8x, ZN 
                           => n3891);
   U4299 : AOI22_X1 port map( A1 => n5268, A2 => fromRegsPortxREG_FILE_30xx8x, 
                           B1 => n5375, B2 => fromRegsPortxREG_FILE_02xx8x, ZN 
                           => n3890);
   U4300 : AOI22_X1 port map( A1 => n5211, A2 => fromRegsPortxREG_FILE_23xx8x, 
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx8x, ZN 
                           => n3889);
   U4301 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_24xx8x, 
                           B1 => n5166, B2 => fromRegsPortxREG_FILE_18xx8x, ZN 
                           => n3888);
   U4302 : AND4_X1 port map( A1 => n3891, A2 => n3890, A3 => n3889, A4 => n3888
                           , ZN => n3907);
   U4303 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_20xx8x, 
                           B1 => n5202, B2 => fromRegsPortxREG_FILE_12xx8x, ZN 
                           => n3895);
   U4304 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx8x, 
                           B1 => n5225, B2 => fromRegsPortxREG_FILE_22xx8x, ZN 
                           => n3894);
   U4305 : AOI22_X1 port map( A1 => n5197, A2 => fromRegsPortxREG_FILE_06xx8x, 
                           B1 => n5159, B2 => fromRegsPortxREG_FILE_28xx8x, ZN 
                           => n3893);
   U4306 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx8x, 
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx8x, ZN 
                           => n3892);
   U4307 : AND4_X1 port map( A1 => n3895, A2 => n3894, A3 => n3893, A4 => n3892
                           , ZN => n3906);
   U4308 : AOI22_X1 port map( A1 => n5230, A2 => fromRegsPortxREG_FILE_07xx8x, 
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_11xx8x, ZN 
                           => n3899);
   U4309 : AOI22_X1 port map( A1 => n5369, A2 => fromRegsPortxREG_FILE_10xx8x, 
                           B1 => n5152, B2 => fromRegsPortxREG_FILE_14xx8x, ZN 
                           => n3898);
   U4310 : AOI22_X1 port map( A1 => n3959, A2 => fromRegsPortxREG_FILE_16xx8x, 
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx8x, ZN 
                           => n3897);
   U4311 : AOI22_X1 port map( A1 => n5251, A2 => fromRegsPortxREG_FILE_17xx8x, 
                           B1 => n5160, B2 => fromRegsPortxREG_FILE_15xx8x, ZN 
                           => n3896);
   U4312 : AND4_X1 port map( A1 => n3899, A2 => n3898, A3 => n3897, A4 => n3896
                           , ZN => n3905);
   U4313 : AOI22_X1 port map( A1 => n5235, A2 => fromRegsPortxREG_FILE_09xx8x, 
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx8x, ZN 
                           => n3903);
   U4314 : AOI22_X1 port map( A1 => n5147, A2 => fromRegsPortxREG_FILE_08xx8x, 
                           B1 => n5153, B2 => fromRegsPortxREG_FILE_29xx8x, ZN 
                           => n3902);
   U4315 : NAND2_X1 port map( A1 => n5367, A2 => fromRegsPortxREG_FILE_19xx8x, 
                           ZN => n3901);
   U4316 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_31xx8x, 
                           B1 => n5261, B2 => fromRegsPortxREG_FILE_27xx8x, ZN 
                           => n3900);
   U4317 : AND4_X1 port map( A1 => n3903, A2 => n3902, A3 => n3901, A4 => n3900
                           , ZN => n3904);
   U4318 : NAND4_X1 port map( A1 => n3907, A2 => n3906, A3 => n3905, A4 => 
                           n3904, ZN => ashr_25xAx8x);
   U4319 : AOI22_X1 port map( A1 => n3959, A2 => fromRegsPortxREG_FILE_16xx9x, 
                           B1 => n5166, B2 => fromRegsPortxREG_FILE_18xx9x, ZN 
                           => n3911);
   U4320 : AOI22_X1 port map( A1 => n5160, A2 => fromRegsPortxREG_FILE_15xx9x, 
                           B1 => n5375, B2 => fromRegsPortxREG_FILE_02xx9x, ZN 
                           => n3910);
   U4321 : AOI22_X1 port map( A1 => n5211, A2 => fromRegsPortxREG_FILE_23xx9x, 
                           B1 => n5246, B2 => fromRegsPortxREG_FILE_13xx9x, ZN 
                           => n3909);
   U4322 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_20xx9x, 
                           B1 => n5152, B2 => fromRegsPortxREG_FILE_14xx9x, ZN 
                           => n3908);
   U4323 : AND4_X1 port map( A1 => n3911, A2 => n3910, A3 => n3909, A4 => n3908
                           , ZN => n3927);
   U4324 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx9x, 
                           B1 => n5251, B2 => fromRegsPortxREG_FILE_17xx9x, ZN 
                           => n3915);
   U4325 : AOI22_X1 port map( A1 => n5176, A2 => fromRegsPortxREG_FILE_03xx9x, 
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx9x, ZN 
                           => n3914);
   U4326 : AOI22_X1 port map( A1 => n5252, A2 => fromRegsPortxREG_FILE_04xx9x, 
                           B1 => n5202, B2 => fromRegsPortxREG_FILE_12xx9x, ZN 
                           => n3913);
   U4327 : AOI22_X1 port map( A1 => n5153, A2 => fromRegsPortxREG_FILE_29xx9x, 
                           B1 => n5159, B2 => fromRegsPortxREG_FILE_28xx9x, ZN 
                           => n3912);
   U4328 : AND4_X1 port map( A1 => n3915, A2 => n3914, A3 => n3913, A4 => n3912
                           , ZN => n3926);
   U4329 : AOI22_X1 port map( A1 => n5261, A2 => fromRegsPortxREG_FILE_27xx9x, 
                           B1 => n5167, B2 => fromRegsPortxREG_FILE_10xx9x, ZN 
                           => n3919);
   U4330 : AOI22_X1 port map( A1 => n5259, A2 => fromRegsPortxREG_FILE_21xx9x, 
                           B1 => n5244, B2 => fromRegsPortxREG_FILE_19xx9x, ZN 
                           => n3918);
   U4331 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_31xx9x, 
                           B1 => n5235, B2 => fromRegsPortxREG_FILE_09xx9x, ZN 
                           => n3917);
   U4332 : AOI22_X1 port map( A1 => n5220, A2 => fromRegsPortxREG_FILE_05xx9x, 
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_11xx9x, ZN 
                           => n3916);
   U4333 : AND4_X1 port map( A1 => n3919, A2 => n3918, A3 => n3917, A4 => n3916
                           , ZN => n3925);
   U4334 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx9x, 
                           B1 => n5230, B2 => fromRegsPortxREG_FILE_07xx9x, ZN 
                           => n3923);
   U4335 : AOI22_X1 port map( A1 => n5197, A2 => fromRegsPortxREG_FILE_06xx9x, 
                           B1 => n5266, B2 => fromRegsPortxREG_FILE_24xx9x, ZN 
                           => n3922);
   U4336 : AOI22_X1 port map( A1 => n5147, A2 => fromRegsPortxREG_FILE_08xx9x, 
                           B1 => n5268, B2 => fromRegsPortxREG_FILE_30xx9x, ZN 
                           => n3921);
   U4337 : NAND2_X1 port map( A1 => n5245, A2 => fromRegsPortxREG_FILE_26xx9x, 
                           ZN => n3920);
   U4338 : AND4_X1 port map( A1 => n3923, A2 => n3922, A3 => n3921, A4 => n3920
                           , ZN => n3924);
   U4339 : NAND4_X1 port map( A1 => n3927, A2 => n3926, A3 => n3925, A4 => 
                           n3924, ZN => ashr_25xAx9x);
   U4340 : AOI22_X1 port map( A1 => n5147, A2 => fromRegsPortxREG_FILE_08xx10x,
                           B1 => n5197, B2 => fromRegsPortxREG_FILE_06xx10x, ZN
                           => n3931);
   U4341 : AOI22_X1 port map( A1 => n5153, A2 => fromRegsPortxREG_FILE_29xx10x,
                           B1 => n5176, B2 => fromRegsPortxREG_FILE_03xx10x, ZN
                           => n3930);
   U4342 : AOI22_X1 port map( A1 => n5356, A2 => fromRegsPortxREG_FILE_12xx10x,
                           B1 => n5244, B2 => fromRegsPortxREG_FILE_19xx10x, ZN
                           => n3929);
   U4343 : AOI22_X1 port map( A1 => n5245, A2 => fromRegsPortxREG_FILE_26xx10x,
                           B1 => n5166, B2 => fromRegsPortxREG_FILE_18xx10x, ZN
                           => n3928);
   U4344 : AND4_X1 port map( A1 => n3931, A2 => n3930, A3 => n3929, A4 => n3928
                           , ZN => n3947);
   U4345 : AOI22_X1 port map( A1 => n5252, A2 => fromRegsPortxREG_FILE_04xx10x,
                           B1 => n5167, B2 => fromRegsPortxREG_FILE_10xx10x, ZN
                           => n3935);
   U4346 : AOI22_X1 port map( A1 => n5260, A2 => fromRegsPortxREG_FILE_02xx10x,
                           B1 => n5152, B2 => fromRegsPortxREG_FILE_14xx10x, ZN
                           => n3934);
   U4347 : AOI22_X1 port map( A1 => n5251, A2 => fromRegsPortxREG_FILE_17xx10x,
                           B1 => n5211, B2 => fromRegsPortxREG_FILE_23xx10x, ZN
                           => n3933);
   U4348 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx10x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx10x, ZN
                           => n3932);
   U4349 : AND4_X1 port map( A1 => n3935, A2 => n3934, A3 => n3933, A4 => n3932
                           , ZN => n3946);
   U4350 : AOI22_X1 port map( A1 => n3959, A2 => fromRegsPortxREG_FILE_16xx10x,
                           B1 => n5160, B2 => fromRegsPortxREG_FILE_15xx10x, ZN
                           => n3939);
   U4351 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_31xx10x,
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx10x, ZN
                           => n3938);
   U4352 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_28xx10x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx10x, ZN
                           => n3937);
   U4353 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_20xx10x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx10x, ZN
                           => n3936);
   U4354 : AND4_X1 port map( A1 => n3939, A2 => n3938, A3 => n3937, A4 => n3936
                           , ZN => n3945);
   U4355 : AOI22_X1 port map( A1 => n5268, A2 => fromRegsPortxREG_FILE_30xx10x,
                           B1 => n5230, B2 => fromRegsPortxREG_FILE_07xx10x, ZN
                           => n3943);
   U4356 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx10x,
                           B1 => n5266, B2 => fromRegsPortxREG_FILE_24xx10x, ZN
                           => n3942);
   U4357 : NAND2_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_01xx10x,
                           ZN => n3941);
   U4358 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_11xx10x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx10x, ZN
                           => n3940);
   U4359 : AND4_X1 port map( A1 => n3943, A2 => n3942, A3 => n3941, A4 => n3940
                           , ZN => n3944);
   U4360 : NAND4_X1 port map( A1 => n3947, A2 => n3946, A3 => n3945, A4 => 
                           n3944, ZN => ashr_25xAx10x);
   U4361 : AOI22_X1 port map( A1 => n5153, A2 => fromRegsPortxREG_FILE_29xx13x,
                           B1 => n5166, B2 => fromRegsPortxREG_FILE_18xx13x, ZN
                           => n3951);
   U4362 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx13x,
                           B1 => n5375, B2 => fromRegsPortxREG_FILE_02xx13x, ZN
                           => n3950);
   U4363 : AOI22_X1 port map( A1 => n5197, A2 => fromRegsPortxREG_FILE_06xx13x,
                           B1 => n5244, B2 => fromRegsPortxREG_FILE_19xx13x, ZN
                           => n3949);
   U4364 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx13x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx13x, ZN
                           => n3948);
   U4365 : AND4_X1 port map( A1 => n3951, A2 => n3950, A3 => n3949, A4 => n3948
                           , ZN => n3970);
   U4366 : AOI22_X1 port map( A1 => n5252, A2 => fromRegsPortxREG_FILE_04xx13x,
                           B1 => n5225, B2 => fromRegsPortxREG_FILE_22xx13x, ZN
                           => n3953);
   U4367 : AOI22_X1 port map( A1 => n5159, A2 => fromRegsPortxREG_FILE_28xx13x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_21xx13x, ZN
                           => n3952);
   U4368 : NAND2_X1 port map( A1 => n3953, A2 => n3952, ZN => n3958);
   U4369 : AOI22_X1 port map( A1 => n5147, A2 => fromRegsPortxREG_FILE_08xx13x,
                           B1 => n5202, B2 => fromRegsPortxREG_FILE_12xx13x, ZN
                           => n3956);
   U4370 : NAND2_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_11xx13x,
                           ZN => n3955);
   U4371 : AOI22_X1 port map( A1 => n5261, A2 => fromRegsPortxREG_FILE_27xx13x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx13x, ZN
                           => n3954);
   U4372 : NAND3_X1 port map( A1 => n3956, A2 => n3955, A3 => n3954, ZN => 
                           n3957);
   U4373 : NOR2_X1 port map( A1 => n3958, A2 => n3957, ZN => n3969);
   U4374 : AOI22_X1 port map( A1 => n3959, A2 => fromRegsPortxREG_FILE_16xx13x,
                           B1 => n5152, B2 => fromRegsPortxREG_FILE_14xx13x, ZN
                           => n3963);
   U4375 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_31xx13x,
                           B1 => n5167, B2 => fromRegsPortxREG_FILE_10xx13x, ZN
                           => n3962);
   U4376 : AOI22_X1 port map( A1 => n5251, A2 => fromRegsPortxREG_FILE_17xx13x,
                           B1 => n5211, B2 => fromRegsPortxREG_FILE_23xx13x, ZN
                           => n3961);
   U4377 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_24xx13x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx13x, ZN
                           => n3960);
   U4378 : AND4_X1 port map( A1 => n3963, A2 => n3962, A3 => n3961, A4 => n3960
                           , ZN => n3968);
   U4379 : AOI22_X1 port map( A1 => n5176, A2 => fromRegsPortxREG_FILE_03xx13x,
                           B1 => n5165, B2 => fromRegsPortxREG_FILE_20xx13x, ZN
                           => n3966);
   U4380 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx13x,
                           B1 => n5230, B2 => fromRegsPortxREG_FILE_07xx13x, ZN
                           => n3965);
   U4381 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx13x,
                           B1 => n5220, B2 => fromRegsPortxREG_FILE_05xx13x, ZN
                           => n3964);
   U4382 : AND3_X1 port map( A1 => n3966, A2 => n3965, A3 => n3964, ZN => n3967
                           );
   U4383 : NAND4_X1 port map( A1 => n3970, A2 => n3969, A3 => n3968, A4 => 
                           n3967, ZN => ashr_25xAx13x);
   U4384 : AOI22_X1 port map( A1 => n5197, A2 => fromRegsPortxREG_FILE_06xx15x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx15x, ZN
                           => n3974);
   U4385 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_20xx15x,
                           B1 => n5152, B2 => fromRegsPortxREG_FILE_14xx15x, ZN
                           => n3973);
   U4386 : AOI22_X1 port map( A1 => n5367, A2 => fromRegsPortxREG_FILE_19xx15x,
                           B1 => n5167, B2 => fromRegsPortxREG_FILE_10xx15x, ZN
                           => n3972);
   U4387 : AOI22_X1 port map( A1 => n5176, A2 => fromRegsPortxREG_FILE_03xx15x,
                           B1 => n5211, B2 => fromRegsPortxREG_FILE_23xx15x, ZN
                           => n3971);
   U4388 : AND4_X1 port map( A1 => n3974, A2 => n3973, A3 => n3972, A4 => n3971
                           , ZN => n3990);
   U4389 : AOI22_X1 port map( A1 => n5260, A2 => fromRegsPortxREG_FILE_02xx15x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_11xx15x, ZN
                           => n3978);
   U4390 : AOI22_X1 port map( A1 => n5159, A2 => fromRegsPortxREG_FILE_28xx15x,
                           B1 => n5225, B2 => fromRegsPortxREG_FILE_22xx15x, ZN
                           => n3977);
   U4391 : AOI22_X1 port map( A1 => n5259, A2 => fromRegsPortxREG_FILE_21xx15x,
                           B1 => n5202, B2 => fromRegsPortxREG_FILE_12xx15x, ZN
                           => n3976);
   U4392 : AOI22_X1 port map( A1 => n5251, A2 => fromRegsPortxREG_FILE_17xx15x,
                           B1 => n5235, B2 => fromRegsPortxREG_FILE_09xx15x, ZN
                           => n3975);
   U4393 : AND4_X1 port map( A1 => n3978, A2 => n3977, A3 => n3976, A4 => n3975
                           , ZN => n3989);
   U4394 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx15x,
                           B1 => n5261, B2 => fromRegsPortxREG_FILE_27xx15x, ZN
                           => n3982);
   U4395 : AOI22_X1 port map( A1 => n5220, A2 => fromRegsPortxREG_FILE_05xx15x,
                           B1 => n5245, B2 => fromRegsPortxREG_FILE_26xx15x, ZN
                           => n3981);
   U4396 : AOI22_X1 port map( A1 => n5267, A2 => fromRegsPortxREG_FILE_25xx15x,
                           B1 => n5153, B2 => fromRegsPortxREG_FILE_29xx15x, ZN
                           => n3980);
   U4397 : NAND2_X1 port map( A1 => n5147, A2 => fromRegsPortxREG_FILE_08xx15x,
                           ZN => n3979);
   U4398 : AND4_X1 port map( A1 => n3982, A2 => n3981, A3 => n3980, A4 => n3979
                           , ZN => n3988);
   U4399 : AOI22_X1 port map( A1 => n5252, A2 => fromRegsPortxREG_FILE_04xx15x,
                           B1 => n5166, B2 => fromRegsPortxREG_FILE_18xx15x, ZN
                           => n3986);
   U4400 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx15x,
                           B1 => n5230, B2 => fromRegsPortxREG_FILE_07xx15x, ZN
                           => n3985);
   U4401 : AOI22_X1 port map( A1 => n5160, A2 => fromRegsPortxREG_FILE_15xx15x,
                           B1 => n5266, B2 => fromRegsPortxREG_FILE_24xx15x, ZN
                           => n3984);
   U4402 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx15x,
                           B1 => n5158, B2 => fromRegsPortxREG_FILE_31xx15x, ZN
                           => n3983);
   U4403 : AND4_X1 port map( A1 => n3986, A2 => n3985, A3 => n3984, A4 => n3983
                           , ZN => n3987);
   U4404 : NAND4_X1 port map( A1 => n3990, A2 => n3989, A3 => n3988, A4 => 
                           n3987, ZN => ashr_25xAx15x);
   U4405 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx16x,
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx16x, ZN
                           => n3994);
   U4406 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx16x,
                           B1 => n5202, B2 => fromRegsPortxREG_FILE_12xx16x, ZN
                           => n3993);
   U4407 : AOI22_X1 port map( A1 => n5160, A2 => fromRegsPortxREG_FILE_15xx16x,
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_28xx16x, ZN
                           => n3992);
   U4408 : AOI22_X1 port map( A1 => n5197, A2 => fromRegsPortxREG_FILE_06xx16x,
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx16x, ZN
                           => n3991);
   U4409 : AND4_X1 port map( A1 => n3994, A2 => n3993, A3 => n3992, A4 => n3991
                           , ZN => n4010);
   U4410 : AOI22_X1 port map( A1 => n5225, A2 => fromRegsPortxREG_FILE_22xx16x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx16x, ZN
                           => n3998);
   U4411 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_11xx16x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx16x, ZN
                           => n3997);
   U4412 : AOI22_X1 port map( A1 => n5153, A2 => fromRegsPortxREG_FILE_29xx16x,
                           B1 => n5253, B2 => fromRegsPortxREG_FILE_01xx16x, ZN
                           => n3996);
   U4413 : AOI22_X1 port map( A1 => n5220, A2 => fromRegsPortxREG_FILE_05xx16x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx16x, ZN
                           => n3995);
   U4414 : AND4_X1 port map( A1 => n3998, A2 => n3997, A3 => n3996, A4 => n3995
                           , ZN => n4009);
   U4415 : AOI22_X1 port map( A1 => n5176, A2 => fromRegsPortxREG_FILE_03xx16x,
                           B1 => n5260, B2 => fromRegsPortxREG_FILE_02xx16x, ZN
                           => n4002);
   U4416 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx16x,
                           B1 => n5244, B2 => fromRegsPortxREG_FILE_19xx16x, ZN
                           => n4001);
   U4417 : AOI22_X1 port map( A1 => n5251, A2 => fromRegsPortxREG_FILE_17xx16x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx16x, ZN
                           => n4000);
   U4418 : AOI22_X1 port map( A1 => n5379, A2 => fromRegsPortxREG_FILE_31xx16x,
                           B1 => n5266, B2 => fromRegsPortxREG_FILE_24xx16x, ZN
                           => n3999);
   U4419 : AND4_X1 port map( A1 => n4002, A2 => n4001, A3 => n4000, A4 => n3999
                           , ZN => n4008);
   U4420 : AOI22_X1 port map( A1 => n5211, A2 => fromRegsPortxREG_FILE_23xx16x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx16x, ZN
                           => n4006);
   U4421 : AOI22_X1 port map( A1 => n5230, A2 => fromRegsPortxREG_FILE_07xx16x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx16x, ZN
                           => n4005);
   U4422 : AOI22_X1 port map( A1 => n5267, A2 => fromRegsPortxREG_FILE_25xx16x,
                           B1 => n5268, B2 => fromRegsPortxREG_FILE_30xx16x, ZN
                           => n4004);
   U4423 : NAND2_X1 port map( A1 => n5368, A2 => fromRegsPortxREG_FILE_14xx16x,
                           ZN => n4003);
   U4424 : AND4_X1 port map( A1 => n4006, A2 => n4005, A3 => n4004, A4 => n4003
                           , ZN => n4007);
   U4425 : NAND4_X1 port map( A1 => n4010, A2 => n4009, A3 => n4008, A4 => 
                           n4007, ZN => ashr_25xAx16x);
   U4426 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx20x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx20x, ZN
                           => n4014);
   U4427 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx20x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx20x, ZN
                           => n4013);
   U4428 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx20x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx20x, ZN
                           => n4012);
   U4429 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx20x,
                           B1 => n5246, B2 => fromRegsPortxREG_FILE_13xx20x, ZN
                           => n4011);
   U4430 : AND4_X1 port map( A1 => n4014, A2 => n4013, A3 => n4012, A4 => n4011
                           , ZN => n4030);
   U4431 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx20x,
                           B1 => n5345, B2 => fromRegsPortxREG_FILE_16xx20x, ZN
                           => n4018);
   U4432 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx20x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx20x, ZN
                           => n4017);
   U4433 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx20x,
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_28xx20x, ZN
                           => n4016);
   U4434 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx20x,
                           B1 => n5202, B2 => fromRegsPortxREG_FILE_12xx20x, ZN
                           => n4015);
   U4435 : AND4_X1 port map( A1 => n4018, A2 => n4017, A3 => n4016, A4 => n4015
                           , ZN => n4029);
   U4436 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx20x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_11xx20x, ZN
                           => n4022);
   U4437 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx20x,
                           B1 => n5244, B2 => fromRegsPortxREG_FILE_19xx20x, ZN
                           => n4021);
   U4438 : AOI22_X1 port map( A1 => n5230, A2 => fromRegsPortxREG_FILE_07xx20x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_21xx20x, ZN
                           => n4020);
   U4439 : AOI22_X1 port map( A1 => n5267, A2 => fromRegsPortxREG_FILE_25xx20x,
                           B1 => n5211, B2 => fromRegsPortxREG_FILE_23xx20x, ZN
                           => n4019);
   U4440 : AND4_X1 port map( A1 => n4022, A2 => n4021, A3 => n4020, A4 => n4019
                           , ZN => n4028);
   U4441 : AOI22_X1 port map( A1 => n5379, A2 => fromRegsPortxREG_FILE_31xx20x,
                           B1 => n5266, B2 => fromRegsPortxREG_FILE_24xx20x, ZN
                           => n4026);
   U4442 : AOI22_X1 port map( A1 => n5357, A2 => fromRegsPortxREG_FILE_04xx20x,
                           B1 => n5245, B2 => fromRegsPortxREG_FILE_26xx20x, ZN
                           => n4025);
   U4443 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_02xx20x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx20x, ZN
                           => n4024);
   U4444 : NAND2_X1 port map( A1 => n5235, A2 => fromRegsPortxREG_FILE_09xx20x,
                           ZN => n4023);
   U4445 : AND4_X1 port map( A1 => n4026, A2 => n4025, A3 => n4024, A4 => n4023
                           , ZN => n4027);
   U4446 : NAND4_X1 port map( A1 => n4030, A2 => n4029, A3 => n4028, A4 => 
                           n4027, ZN => ashr_25xAx20x);
   U4447 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx21x,
                           B1 => n5379, B2 => fromRegsPortxREG_FILE_31xx21x, ZN
                           => n4034);
   U4448 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx21x,
                           B1 => n5268, B2 => fromRegsPortxREG_FILE_30xx21x, ZN
                           => n4033);
   U4449 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx21x,
                           B1 => n5245, B2 => fromRegsPortxREG_FILE_26xx21x, ZN
                           => n4032);
   U4450 : NAND2_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_27xx21x,
                           ZN => n4031);
   U4451 : AND4_X1 port map( A1 => n4034, A2 => n4033, A3 => n4032, A4 => n4031
                           , ZN => n4050);
   U4452 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_02xx21x,
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx21x, ZN
                           => n4038);
   U4453 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_24xx21x,
                           B1 => n5225, B2 => fromRegsPortxREG_FILE_22xx21x, ZN
                           => n4037);
   U4454 : AOI22_X1 port map( A1 => n5235, A2 => fromRegsPortxREG_FILE_09xx21x,
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx21x, ZN
                           => n4036);
   U4455 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx21x,
                           B1 => n5202, B2 => fromRegsPortxREG_FILE_12xx21x, ZN
                           => n4035);
   U4456 : AND4_X1 port map( A1 => n4038, A2 => n4037, A3 => n4036, A4 => n4035
                           , ZN => n4049);
   U4457 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx21x,
                           B1 => n5367, B2 => fromRegsPortxREG_FILE_19xx21x, ZN
                           => n4042);
   U4458 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx21x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx21x, ZN
                           => n4041);
   U4459 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx21x,
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_23xx21x, ZN
                           => n4040);
   U4460 : AOI22_X1 port map( A1 => n5267, A2 => fromRegsPortxREG_FILE_25xx21x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_11xx21x, ZN
                           => n4039);
   U4461 : AND4_X1 port map( A1 => n4042, A2 => n4041, A3 => n4040, A4 => n4039
                           , ZN => n4048);
   U4462 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx21x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx21x, ZN
                           => n4046);
   U4463 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx21x,
                           B1 => n5246, B2 => fromRegsPortxREG_FILE_13xx21x, ZN
                           => n4045);
   U4464 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx21x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx21x, ZN
                           => n4044);
   U4465 : AOI22_X1 port map( A1 => n5159, A2 => fromRegsPortxREG_FILE_28xx21x,
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx21x, ZN
                           => n4043);
   U4466 : AND4_X1 port map( A1 => n4046, A2 => n4045, A3 => n4044, A4 => n4043
                           , ZN => n4047);
   U4467 : NAND4_X1 port map( A1 => n4050, A2 => n4049, A3 => n4048, A4 => 
                           n4047, ZN => ashr_25xAx21x);
   U4468 : AOI22_X1 port map( A1 => n5267, A2 => fromRegsPortxREG_FILE_25xx23x,
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_06xx23x, ZN
                           => n4054);
   U4469 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx23x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx23x, ZN
                           => n4053);
   U4470 : AOI22_X1 port map( A1 => n5340, A2 => fromRegsPortxREG_FILE_09xx23x,
                           B1 => n5367, B2 => fromRegsPortxREG_FILE_19xx23x, ZN
                           => n4052);
   U4471 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx23x,
                           B1 => n5246, B2 => fromRegsPortxREG_FILE_13xx23x, ZN
                           => n4051);
   U4472 : AND4_X1 port map( A1 => n4054, A2 => n4053, A3 => n4052, A4 => n4051
                           , ZN => n4070);
   U4473 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx23x,
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx23x, ZN
                           => n4058);
   U4474 : AOI22_X1 port map( A1 => n5261, A2 => fromRegsPortxREG_FILE_27xx23x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx23x, ZN
                           => n4057);
   U4475 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx23x,
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx23x, ZN
                           => n4056);
   U4476 : AOI22_X1 port map( A1 => n5379, A2 => fromRegsPortxREG_FILE_31xx23x,
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_28xx23x, ZN
                           => n4055);
   U4477 : AND4_X1 port map( A1 => n4058, A2 => n4057, A3 => n4056, A4 => n4055
                           , ZN => n4069);
   U4478 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx23x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx23x, ZN
                           => n4062);
   U4479 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_02xx23x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx23x, ZN
                           => n4061);
   U4480 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx23x,
                           B1 => n5380, B2 => fromRegsPortxREG_FILE_01xx23x, ZN
                           => n4060);
   U4481 : AOI22_X1 port map( A1 => n5343, A2 => fromRegsPortxREG_FILE_07xx23x,
                           B1 => n5341, B2 => fromRegsPortxREG_FILE_11xx23x, ZN
                           => n4059);
   U4482 : AND4_X1 port map( A1 => n4062, A2 => n4061, A3 => n4060, A4 => n4059
                           , ZN => n4068);
   U4483 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx23x,
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_24xx23x, ZN
                           => n4066);
   U4484 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx23x,
                           B1 => n5245, B2 => fromRegsPortxREG_FILE_26xx23x, ZN
                           => n4065);
   U4485 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx23x,
                           B1 => n5351, B2 => fromRegsPortxREG_FILE_29xx23x, ZN
                           => n4064);
   U4486 : NAND2_X1 port map( A1 => n5356, A2 => fromRegsPortxREG_FILE_12xx23x,
                           ZN => n4063);
   U4487 : AND4_X1 port map( A1 => n4066, A2 => n4065, A3 => n4064, A4 => n4063
                           , ZN => n4067);
   U4488 : NAND4_X1 port map( A1 => n4070, A2 => n4069, A3 => n4068, A4 => 
                           n4067, ZN => ashr_25xAx23x);
   U4489 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx24x,
                           B1 => n5379, B2 => fromRegsPortxREG_FILE_31xx24x, ZN
                           => n4074);
   U4490 : AOI22_X1 port map( A1 => n5252, A2 => fromRegsPortxREG_FILE_04xx24x,
                           B1 => n5245, B2 => fromRegsPortxREG_FILE_26xx24x, ZN
                           => n4073);
   U4491 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx24x,
                           B1 => n5261, B2 => fromRegsPortxREG_FILE_27xx24x, ZN
                           => n4072);
   U4492 : NAND2_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx24x,
                           ZN => n4071);
   U4493 : AND4_X1 port map( A1 => n4074, A2 => n4073, A3 => n4072, A4 => n4071
                           , ZN => n4090);
   U4494 : AOI22_X1 port map( A1 => n5364, A2 => fromRegsPortxREG_FILE_18xx24x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx24x, ZN
                           => n4078);
   U4495 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_02xx24x,
                           B1 => n5246, B2 => fromRegsPortxREG_FILE_13xx24x, ZN
                           => n4077);
   U4496 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx24x,
                           B1 => n5380, B2 => fromRegsPortxREG_FILE_01xx24x, ZN
                           => n4076);
   U4497 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx24x,
                           B1 => n5341, B2 => fromRegsPortxREG_FILE_11xx24x, ZN
                           => n4075);
   U4498 : AND4_X1 port map( A1 => n4078, A2 => n4077, A3 => n4076, A4 => n4075
                           , ZN => n4089);
   U4499 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx24x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx24x, ZN
                           => n4082);
   U4500 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx24x,
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_28xx24x, ZN
                           => n4081);
   U4501 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx24x,
                           B1 => n5356, B2 => fromRegsPortxREG_FILE_12xx24x, ZN
                           => n4080);
   U4502 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx24x,
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_23xx24x, ZN
                           => n4079);
   U4503 : AND4_X1 port map( A1 => n4082, A2 => n4081, A3 => n4080, A4 => n4079
                           , ZN => n4088);
   U4504 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx24x,
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx24x, ZN
                           => n4086);
   U4505 : AOI22_X1 port map( A1 => n5342, A2 => fromRegsPortxREG_FILE_21xx24x,
                           B1 => n5367, B2 => fromRegsPortxREG_FILE_19xx24x, ZN
                           => n4085);
   U4506 : AOI22_X1 port map( A1 => n5225, A2 => fromRegsPortxREG_FILE_22xx24x,
                           B1 => n5152, B2 => fromRegsPortxREG_FILE_14xx24x, ZN
                           => n4084);
   U4507 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx24x,
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_24xx24x, ZN
                           => n4083);
   U4508 : AND4_X1 port map( A1 => n4086, A2 => n4085, A3 => n4084, A4 => n4083
                           , ZN => n4087);
   U4509 : NAND4_X1 port map( A1 => n4090, A2 => n4089, A3 => n4088, A4 => 
                           n4087, ZN => ashr_25xAx24x);
   U4510 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx25x,
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_24xx25x, ZN
                           => n4094);
   U4511 : AOI22_X1 port map( A1 => n5356, A2 => fromRegsPortxREG_FILE_12xx25x,
                           B1 => n5245, B2 => fromRegsPortxREG_FILE_26xx25x, ZN
                           => n4093);
   U4512 : NAND2_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx25x,
                           ZN => n4092);
   U4513 : AOI22_X1 port map( A1 => n5379, A2 => fromRegsPortxREG_FILE_31xx25x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx25x, ZN
                           => n4091);
   U4514 : AND4_X1 port map( A1 => n4094, A2 => n4093, A3 => n4092, A4 => n4091
                           , ZN => n4110);
   U4515 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx25x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_21xx25x, ZN
                           => n4098);
   U4516 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx25x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx25x, ZN
                           => n4097);
   U4517 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx25x,
                           B1 => n5354, B2 => fromRegsPortxREG_FILE_20xx25x, ZN
                           => n4096);
   U4518 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx25x,
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx25x, ZN
                           => n4095);
   U4519 : AND4_X1 port map( A1 => n4098, A2 => n4097, A3 => n4096, A4 => n4095
                           , ZN => n4109);
   U4520 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx25x,
                           B1 => n5246, B2 => fromRegsPortxREG_FILE_13xx25x, ZN
                           => n4102);
   U4521 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx25x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx25x, ZN
                           => n4101);
   U4522 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx25x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx25x, ZN
                           => n4100);
   U4523 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_02xx25x,
                           B1 => n5341, B2 => fromRegsPortxREG_FILE_11xx25x, ZN
                           => n4099);
   U4524 : AND4_X1 port map( A1 => n4102, A2 => n4101, A3 => n4100, A4 => n4099
                           , ZN => n4108);
   U4525 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_28xx25x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx25x, ZN
                           => n4106);
   U4526 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx25x,
                           B1 => n5367, B2 => fromRegsPortxREG_FILE_19xx25x, ZN
                           => n4105);
   U4527 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx25x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx25x, ZN
                           => n4104);
   U4528 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx25x,
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx25x, ZN
                           => n4103);
   U4529 : AND4_X1 port map( A1 => n4106, A2 => n4105, A3 => n4104, A4 => n4103
                           , ZN => n4107);
   U4530 : NAND4_X1 port map( A1 => n4110, A2 => n4109, A3 => n4108, A4 => 
                           n4107, ZN => ashr_25xAx25x);
   U4531 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx27x,
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_05xx27x, ZN
                           => n4114);
   U4532 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx27x,
                           B1 => n5355, B2 => fromRegsPortxREG_FILE_03xx27x, ZN
                           => n4113);
   U4533 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx27x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx27x, ZN
                           => n4112);
   U4534 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_28xx27x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx27x, ZN
                           => n4111);
   U4535 : AND4_X1 port map( A1 => n4114, A2 => n4113, A3 => n4112, A4 => n4111
                           , ZN => n4130);
   U4536 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx27x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_21xx27x, ZN
                           => n4118);
   U4537 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx27x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_17xx27x, ZN
                           => n4117);
   U4538 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx27x,
                           B1 => n5356, B2 => fromRegsPortxREG_FILE_12xx27x, ZN
                           => n4116);
   U4539 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_02xx27x,
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx27x, ZN
                           => n4115);
   U4540 : AND4_X1 port map( A1 => n4118, A2 => n4117, A3 => n4116, A4 => n4115
                           , ZN => n4129);
   U4541 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx27x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx27x, ZN
                           => n4122);
   U4542 : AOI22_X1 port map( A1 => n5343, A2 => fromRegsPortxREG_FILE_07xx27x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx27x, ZN
                           => n4121);
   U4543 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_11xx27x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx27x, ZN
                           => n4120);
   U4544 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx27x,
                           B1 => n5367, B2 => fromRegsPortxREG_FILE_19xx27x, ZN
                           => n4119);
   U4545 : AND4_X1 port map( A1 => n4122, A2 => n4121, A3 => n4120, A4 => n4119
                           , ZN => n4128);
   U4546 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx27x,
                           B1 => n5379, B2 => fromRegsPortxREG_FILE_31xx27x, ZN
                           => n4126);
   U4547 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_22xx27x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx27x, ZN
                           => n4125);
   U4548 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_24xx27x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx27x, ZN
                           => n4124);
   U4549 : NAND2_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx27x,
                           ZN => n4123);
   U4550 : AND4_X1 port map( A1 => n4126, A2 => n4125, A3 => n4124, A4 => n4123
                           , ZN => n4127);
   U4551 : NAND4_X1 port map( A1 => n4130, A2 => n4129, A3 => n4128, A4 => 
                           n4127, ZN => ashr_25xAx27x);
   U4552 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx28x,
                           B1 => n5356, B2 => fromRegsPortxREG_FILE_12xx28x, ZN
                           => n4134);
   U4553 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx28x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_21xx28x, ZN
                           => n4133);
   U4554 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx28x,
                           B1 => n5354, B2 => fromRegsPortxREG_FILE_20xx28x, ZN
                           => n4132);
   U4555 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx28x,
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx28x, ZN
                           => n4131);
   U4556 : AND4_X1 port map( A1 => n4134, A2 => n4133, A3 => n4132, A4 => n4131
                           , ZN => n4150);
   U4557 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx28x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx28x, ZN
                           => n4138);
   U4558 : AOI22_X1 port map( A1 => n5366, A2 => fromRegsPortxREG_FILE_13xx28x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx28x, ZN
                           => n4137);
   U4559 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx28x,
                           B1 => n5341, B2 => fromRegsPortxREG_FILE_11xx28x, ZN
                           => n4136);
   U4560 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx28x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx28x, ZN
                           => n4135);
   U4561 : AND4_X1 port map( A1 => n4138, A2 => n4137, A3 => n4136, A4 => n4135
                           , ZN => n4149);
   U4562 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx28x,
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx28x, ZN
                           => n4142);
   U4563 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx28x,
                           B1 => n5367, B2 => fromRegsPortxREG_FILE_19xx28x, ZN
                           => n4141);
   U4564 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_22xx28x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx28x, ZN
                           => n4140);
   U4565 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx28x,
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_24xx28x, ZN
                           => n4139);
   U4566 : AND4_X1 port map( A1 => n4142, A2 => n4141, A3 => n4140, A4 => n4139
                           , ZN => n4148);
   U4567 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx28x,
                           B1 => n5379, B2 => fromRegsPortxREG_FILE_31xx28x, ZN
                           => n4146);
   U4568 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_28xx28x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx28x, ZN
                           => n4145);
   U4569 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_02xx28x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx28x, ZN
                           => n4144);
   U4570 : NAND2_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx28x,
                           ZN => n4143);
   U4571 : AND4_X1 port map( A1 => n4146, A2 => n4145, A3 => n4144, A4 => n4143
                           , ZN => n4147);
   U4572 : NAND4_X1 port map( A1 => n4150, A2 => n4149, A3 => n4148, A4 => 
                           n4147, ZN => ashr_25xAx28x);
   U4573 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx29x,
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_24xx29x, ZN
                           => n4154);
   U4574 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx29x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx29x, ZN
                           => n4153);
   U4575 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx29x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx29x, ZN
                           => n4152);
   U4576 : NAND2_X1 port map( A1 => n5340, A2 => fromRegsPortxREG_FILE_09xx29x,
                           ZN => n4151);
   U4577 : AND4_X1 port map( A1 => n4154, A2 => n4153, A3 => n4152, A4 => n4151
                           , ZN => n4170);
   U4578 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx29x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx29x, ZN
                           => n4158);
   U4579 : AOI22_X1 port map( A1 => n5379, A2 => fromRegsPortxREG_FILE_31xx29x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx29x, ZN
                           => n4157);
   U4580 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx29x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx29x, ZN
                           => n4156);
   U4581 : AOI22_X1 port map( A1 => n5357, A2 => fromRegsPortxREG_FILE_04xx29x,
                           B1 => n5367, B2 => fromRegsPortxREG_FILE_19xx29x, ZN
                           => n4155);
   U4582 : AND4_X1 port map( A1 => n4158, A2 => n4157, A3 => n4156, A4 => n4155
                           , ZN => n4169);
   U4583 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx29x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_21xx29x, ZN
                           => n4162);
   U4584 : AOI22_X1 port map( A1 => n5343, A2 => fromRegsPortxREG_FILE_07xx29x,
                           B1 => n5356, B2 => fromRegsPortxREG_FILE_12xx29x, ZN
                           => n4161);
   U4585 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx29x,
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_28xx29x, ZN
                           => n4160);
   U4586 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx29x,
                           B1 => n5341, B2 => fromRegsPortxREG_FILE_11xx29x, ZN
                           => n4159);
   U4587 : AND4_X1 port map( A1 => n4162, A2 => n4161, A3 => n4160, A4 => n4159
                           , ZN => n4168);
   U4588 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx29x,
                           B1 => n5355, B2 => fromRegsPortxREG_FILE_03xx29x, ZN
                           => n4166);
   U4589 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx29x,
                           B1 => n5375, B2 => fromRegsPortxREG_FILE_02xx29x, ZN
                           => n4165);
   U4590 : AOI22_X1 port map( A1 => n5352, A2 => fromRegsPortxREG_FILE_22xx29x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx29x, ZN
                           => n4164);
   U4591 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx29x,
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_05xx29x, ZN
                           => n4163);
   U4592 : AND4_X1 port map( A1 => n4166, A2 => n4165, A3 => n4164, A4 => n4163
                           , ZN => n4167);
   U4593 : NAND4_X1 port map( A1 => n4170, A2 => n4169, A3 => n4168, A4 => 
                           n4167, ZN => ashr_25xAx29x);
   U4594 : AOI22_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_27xx30x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx30x, ZN
                           => n4174);
   U4595 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx30x,
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_05xx30x, ZN
                           => n4173);
   U4596 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_28xx30x,
                           B1 => n5367, B2 => fromRegsPortxREG_FILE_19xx30x, ZN
                           => n4172);
   U4597 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx30x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx30x, ZN
                           => n4171);
   U4598 : AND4_X1 port map( A1 => n4174, A2 => n4173, A3 => n4172, A4 => n4171
                           , ZN => n4190);
   U4599 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx30x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx30x, ZN
                           => n4178);
   U4600 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx30x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx30x, ZN
                           => n4177);
   U4601 : AOI22_X1 port map( A1 => n5160, A2 => fromRegsPortxREG_FILE_15xx30x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx30x, ZN
                           => n4176);
   U4602 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx30x,
                           B1 => n5380, B2 => fromRegsPortxREG_FILE_01xx30x, ZN
                           => n4175);
   U4603 : AND4_X1 port map( A1 => n4178, A2 => n4177, A3 => n4176, A4 => n4175
                           , ZN => n4189);
   U4604 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx30x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_21xx30x, ZN
                           => n4182);
   U4605 : AOI22_X1 port map( A1 => n5252, A2 => fromRegsPortxREG_FILE_04xx30x,
                           B1 => n5356, B2 => fromRegsPortxREG_FILE_12xx30x, ZN
                           => n4181);
   U4606 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx30x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx30x, ZN
                           => n4180);
   U4607 : AOI22_X1 port map( A1 => n5343, A2 => fromRegsPortxREG_FILE_07xx30x,
                           B1 => n5341, B2 => fromRegsPortxREG_FILE_11xx30x, ZN
                           => n4179);
   U4608 : AND4_X1 port map( A1 => n4182, A2 => n4181, A3 => n4180, A4 => n4179
                           , ZN => n4188);
   U4609 : AOI22_X1 port map( A1 => n5379, A2 => fromRegsPortxREG_FILE_31xx30x,
                           B1 => n5375, B2 => fromRegsPortxREG_FILE_02xx30x, ZN
                           => n4186);
   U4610 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx30x,
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_24xx30x, ZN
                           => n4185);
   U4611 : NAND2_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx30x,
                           ZN => n4184);
   U4612 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx30x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx30x, ZN
                           => n4183);
   U4613 : AND4_X1 port map( A1 => n4186, A2 => n4185, A3 => n4184, A4 => n4183
                           , ZN => n4187);
   U4614 : NAND4_X1 port map( A1 => n4190, A2 => n4189, A3 => n4188, A4 => 
                           n4187, ZN => ashr_25xAx30x);
   U4615 : NOR2_X1 port map( A1 => toRegsPortxDSTxx0x, A2 => n7540, ZN => n4192
                           );
   U4616 : NAND3_X1 port map( A1 => n7534, A2 => n7537, A3 => 
                           toRegsPortxDSTxx3x, ZN => n7514);
   U4617 : OR2_X1 port map( A1 => n7539, A2 => n7514, ZN => n7499);
   U4618 : INV_X1 port map( A => n7499, ZN => n4191);
   U4619 : AOI21_X1 port map( B1 => n4192, B2 => n4191, A => rst, ZN => n4193);
   U4620 : INV_X1 port map( A => n4193, ZN => IF_RegsxN698);
   U4621 : NAND2_X1 port map( A1 => n5694, A2 => fromMemoryPortxLOADEDDATAx(30)
                           , ZN => n4194);
   U4622 : NAND2_X1 port map( A1 => n4504, A2 => n4194, ZN => add_x_26xBx30x);
   U4623 : INV_X1 port map( A => add_x_26xBx30x, ZN => intadd_28xBx2x);
   U4624 : OR2_X1 port map( A1 => n5630, A2 => n5632, ZN => n5689);
   U4625 : NOR2_X1 port map( A1 => n5689, A2 => n5716, ZN => n5693);
   U4626 : NAND2_X1 port map( A1 => n5693, A2 => n6022, ZN => n5674);
   U4627 : CLKBUF_X1 port map( A => n5674, Z => n5679);
   U4628 : AOI21_X1 port map( B1 => n5693, B2 => n6020, A => n7550, ZN => n5677
                           );
   U4629 : CLKBUF_X1 port map( A => n5677, Z => n5678);
   U4630 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(21), ZN => n5737);
   U4631 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(20), A2 => n5737
                           , ZN => n4199);
   U4632 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4199,
                           ZN => n5080);
   U4633 : CLKBUF_X1 port map( A => n5080, Z => n5278);
   U4634 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(20), ZN => n6954);
   U4635 : NAND2_X1 port map( A1 => n5737, A2 => n6954, ZN => n4208);
   U4636 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4208,
                           ZN => n5013);
   U4637 : CLKBUF_X1 port map( A => n5013, Z => n5282);
   U4638 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx30x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_24xx30x, ZN
                           => n4198);
   U4639 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(23), A2 => 
                           fromMemoryPortxLOADEDDATAx(22), ZN => n4219);
   U4640 : NOR2_X1 port map( A1 => n4219, A2 => n4199, ZN => n4945);
   U4641 : CLKBUF_X1 port map( A => n4945, Z => n5280);
   U4642 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(21), A2 => n6954
                           , ZN => n4200);
   U4643 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4200,
                           ZN => n4980);
   U4644 : CLKBUF_X1 port map( A => n4980, Z => n5279);
   U4645 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx30x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx30x, ZN
                           => n4197);
   U4646 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(21), A2 => 
                           fromMemoryPortxLOADEDDATAx(20), ZN => n4201);
   U4647 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4201,
                           ZN => n5012);
   U4648 : CLKBUF_X1 port map( A => n5012, Z => n5281);
   U4649 : NOR2_X1 port map( A1 => n4219, A2 => n4208, ZN => n4978);
   U4650 : CLKBUF_X1 port map( A => n4978, Z => n5283);
   U4651 : AOI22_X1 port map( A1 => n5281, A2 => fromRegsPortxREG_FILE_27xx30x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx30x, ZN
                           => n4196);
   U4652 : NOR2_X1 port map( A1 => n4219, A2 => n4200, ZN => n4979);
   U4653 : CLKBUF_X1 port map( A => n4979, Z => n5277);
   U4654 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(22), ZN => n6995);
   U4655 : NOR3_X1 port map( A1 => n5277, A2 => n6995, A3 => n5737, ZN => n4946
                           );
   U4656 : CLKBUF_X1 port map( A => n4946, Z => n5284);
   U4657 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx30x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx30x, ZN
                           => n4195);
   U4658 : NAND4_X1 port map( A1 => n4198, A2 => n4197, A3 => n4196, A4 => 
                           n4195, ZN => n4207);
   U4659 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(23), ZN => n7033);
   U4660 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n7033
                           , ZN => n4228);
   U4661 : NOR2_X1 port map( A1 => n4199, A2 => n4228, ZN => n5052);
   U4662 : CLKBUF_X1 port map( A => n5052, Z => n5290);
   U4663 : NAND2_X1 port map( A1 => n7033, A2 => n6995, ZN => n4215);
   U4664 : NOR2_X1 port map( A1 => n4199, A2 => n4215, ZN => n5018);
   U4665 : CLKBUF_X1 port map( A => n5018, Z => n5294);
   U4666 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx30x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx30x, ZN
                           => n4205);
   U4667 : NOR2_X1 port map( A1 => n4201, A2 => n4228, ZN => n5019);
   U4668 : CLKBUF_X1 port map( A => n5019, Z => n5291);
   U4669 : NOR2_X1 port map( A1 => n4200, A2 => n4215, ZN => n4986);
   U4670 : CLKBUF_X1 port map( A => n4986, Z => n5295);
   U4671 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx30x,
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx30x, ZN
                           => n4204);
   U4672 : NOR2_X1 port map( A1 => n4208, A2 => n4228, ZN => n4985);
   U4673 : CLKBUF_X1 port map( A => n4985, Z => n5292);
   U4674 : NOR2_X1 port map( A1 => n4200, A2 => n4228, ZN => n5289);
   U4675 : CLKBUF_X1 port map( A => n5289, Z => n5119);
   U4676 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx30x,
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_22xx30x, ZN
                           => n4203);
   U4677 : NOR2_X1 port map( A1 => n4201, A2 => n4215, ZN => n5053);
   U4678 : CLKBUF_X1 port map( A => n5053, Z => n5293);
   U4679 : NAND2_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_19xx30x,
                           ZN => n4202);
   U4680 : NAND4_X1 port map( A1 => n4205, A2 => n4204, A3 => n4203, A4 => 
                           n4202, ZN => n4206);
   U4681 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4207
                           , A => n4206, ZN => n4214);
   U4682 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(24), ZN => n5314);
   U4683 : CLKBUF_X1 port map( A => n5314, Z => n7071);
   U4684 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(21), A2 => 
                           fromMemoryPortxLOADEDDATAx(20), A3 => n7071, ZN => 
                           n4218);
   U4685 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4218,
                           ZN => n4994);
   U4686 : CLKBUF_X1 port map( A => n4994, Z => n5305);
   U4687 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(21), A2 => 
                           fromMemoryPortxLOADEDDATAx(24), ZN => n4220);
   U4688 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(20), A2 => n4220
                           , ZN => n4227);
   U4689 : INV_X1 port map( A => n4227, ZN => n5091);
   U4690 : AOI22_X1 port map( A1 => n5305, A2 => fromRegsPortxREG_FILE_11xx30x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx30x, ZN
                           => n4213);
   U4691 : NAND2_X1 port map( A1 => n6954, A2 => n4220, ZN => n4225);
   U4692 : INV_X1 port map( A => n4225, ZN => n5303);
   U4693 : NAND3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(21), A2 => n7071
                           , A3 => n6954, ZN => n4224);
   U4694 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4224,
                           ZN => n5060);
   U4695 : CLKBUF_X1 port map( A => n5060, Z => n5302);
   U4696 : NOR2_X1 port map( A1 => n4219, A2 => n4224, ZN => n4995);
   U4697 : CLKBUF_X1 port map( A => n4995, Z => n5304);
   U4698 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx30x,
                           B1 => n5304, B2 => fromRegsPortxREG_FILE_14xx30x, ZN
                           => n4210);
   U4699 : NOR2_X1 port map( A1 => n4208, A2 => n4215, ZN => n4957);
   U4700 : CLKBUF_X1 port map( A => n4957, Z => n5311);
   U4701 : NOR2_X1 port map( A1 => n4219, A2 => n4218, ZN => n4993);
   U4702 : CLKBUF_X1 port map( A => n4993, Z => n5307);
   U4703 : AOI22_X1 port map( A1 => n5311, A2 => fromRegsPortxREG_FILE_16xx30x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx30x, ZN
                           => n4209);
   U4704 : NAND2_X1 port map( A1 => n4210, A2 => n4209, ZN => n4211);
   U4705 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx30x, B2 => n5303,
                           A => n4211, ZN => n4212);
   U4706 : OAI211_X1 port map( C1 => n4214, C2 => n5314, A => n4213, B => n4212
                           , ZN => n4222);
   U4707 : NOR2_X1 port map( A1 => n4215, A2 => n4224, ZN => n4760);
   U4708 : CLKBUF_X1 port map( A => n4760, Z => n5329);
   U4709 : INV_X1 port map( A => n4215, ZN => n4216);
   U4710 : NAND2_X1 port map( A1 => n4216, A2 => n4220, ZN => n4233);
   U4711 : INV_X1 port map( A => n4233, ZN => n4217);
   U4712 : NOR2_X1 port map( A1 => n5329, A2 => n4217, ZN => n4973);
   U4713 : CLKBUF_X1 port map( A => n4973, Z => n5334);
   U4714 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(23), A2 => n4218,
                           ZN => n4223);
   U4715 : AOI21_X1 port map( B1 => n4220, B2 => n4219, A => n4223, ZN => n4221
                           );
   U4716 : AND2_X1 port map( A1 => n5334, A2 => n4221, ZN => n5316);
   U4717 : NAND2_X1 port map( A1 => n4222, A2 => n5316, ZN => n4239);
   U4718 : INV_X1 port map( A => n4223, ZN => n4226);
   U4719 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4226,
                           ZN => n5036);
   U4720 : CLKBUF_X1 port map( A => n5036, Z => n5318);
   U4721 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4225,
                           ZN => n4932);
   U4722 : CLKBUF_X1 port map( A => n4932, Z => n5324);
   U4723 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx30x,
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx30x, ZN
                           => n4232);
   U4724 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(22), A2 => n4227,
                           ZN => n5035);
   U4725 : CLKBUF_X1 port map( A => n5035, Z => n5321);
   U4726 : NOR2_X1 port map( A1 => n4228, A2 => n4224, ZN => n5034);
   U4727 : CLKBUF_X1 port map( A => n5034, Z => n5319);
   U4728 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx30x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_06xx30x, ZN
                           => n4231);
   U4729 : NOR2_X1 port map( A1 => n4228, A2 => n4225, ZN => n4965);
   U4730 : CLKBUF_X1 port map( A => n4965, Z => n5320);
   U4731 : NOR2_X1 port map( A1 => n6995, A2 => n4226, ZN => n5033);
   U4732 : CLKBUF_X1 port map( A => n5033, Z => n5322);
   U4733 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx30x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx30x, ZN
                           => n4230);
   U4734 : NOR2_X1 port map( A1 => n4228, A2 => n4227, ZN => n4903);
   U4735 : CLKBUF_X1 port map( A => n4903, Z => n5323);
   U4736 : NAND2_X1 port map( A1 => n5323, A2 => fromRegsPortxREG_FILE_05xx30x,
                           ZN => n4229);
   U4737 : NAND4_X1 port map( A1 => n4232, A2 => n4231, A3 => n4230, A4 => 
                           n4229, ZN => n4237);
   U4738 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx30x,
                           ZN => n4235);
   U4739 : NOR2_X1 port map( A1 => n6954, A2 => n4233, ZN => n5072);
   U4740 : CLKBUF_X1 port map( A => n5072, Z => n5330);
   U4741 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx30x, A2 => n5330,
                           ZN => n4234);
   U4742 : NAND2_X1 port map( A1 => n4235, A2 => n4234, ZN => n4236);
   U4743 : AOI21_X1 port map( B1 => n4237, B2 => n5334, A => n4236, ZN => n4238
                           );
   U4744 : NAND2_X1 port map( A1 => n4239, A2 => n4238, ZN => n7321);
   U4745 : INV_X1 port map( A => n7321, ZN => n7487);
   U4746 : OAI22_X1 port map( A1 => n5679, A2 => intadd_28xBx2x, B1 => n5678, 
                           B2 => n7487, ZN => n4240);
   U4747 : XOR2_X1 port map( A => n7550, B => n4240, Z => 
                           DP_OP_719J14_125_1055xn38);
   U4748 : NAND2_X1 port map( A1 => n5694, A2 => fromMemoryPortxLOADEDDATAx(29)
                           , ZN => n4241);
   U4749 : NAND2_X1 port map( A1 => n4504, A2 => n4241, ZN => add_x_26xBx29x);
   U4750 : INV_X1 port map( A => add_x_26xBx29x, ZN => intadd_28xBx1x);
   U4751 : CLKBUF_X1 port map( A => n4242, Z => n5146);
   U4752 : CLKBUF_X1 port map( A => n5677, Z => n5676);
   U4753 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx29x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_24xx29x, ZN
                           => n4246);
   U4754 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx29x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx29x, ZN
                           => n4245);
   U4755 : AOI22_X1 port map( A1 => n5281, A2 => fromRegsPortxREG_FILE_27xx29x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx29x, ZN
                           => n4244);
   U4756 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx29x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx29x, ZN
                           => n4243);
   U4757 : NAND4_X1 port map( A1 => n4246, A2 => n4245, A3 => n4244, A4 => 
                           n4243, ZN => n4252);
   U4758 : AOI22_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx29x,
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx29x, ZN
                           => n4250);
   U4759 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx29x,
                           B1 => n5290, B2 => fromRegsPortxREG_FILE_21xx29x, ZN
                           => n4249);
   U4760 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx29x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx29x, ZN
                           => n4248);
   U4761 : NAND2_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_19xx29x,
                           ZN => n4247);
   U4762 : NAND4_X1 port map( A1 => n4250, A2 => n4249, A3 => n4248, A4 => 
                           n4247, ZN => n4251);
   U4763 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4252
                           , A => n4251, ZN => n4258);
   U4764 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_12xx29x,
                           B1 => n5304, B2 => fromRegsPortxREG_FILE_14xx29x, ZN
                           => n4257);
   U4765 : AOI22_X1 port map( A1 => n5305, A2 => fromRegsPortxREG_FILE_11xx29x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx29x, ZN
                           => n4254);
   U4766 : CLKBUF_X1 port map( A => n5091, Z => n5306);
   U4767 : AOI22_X1 port map( A1 => n5311, A2 => fromRegsPortxREG_FILE_16xx29x,
                           B1 => n5306, B2 => fromRegsPortxREG_FILE_13xx29x, ZN
                           => n4253);
   U4768 : NAND2_X1 port map( A1 => n4254, A2 => n4253, ZN => n4255);
   U4769 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx29x, B2 => n5302,
                           A => n4255, ZN => n4256);
   U4770 : OAI211_X1 port map( C1 => n4258, C2 => n5314, A => n4257, B => n4256
                           , ZN => n4259);
   U4771 : NAND2_X1 port map( A1 => n4259, A2 => n5316, ZN => n4269);
   U4772 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx29x,
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx29x, ZN
                           => n4263);
   U4773 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx29x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_06xx29x, ZN
                           => n4262);
   U4774 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx29x,
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx29x, ZN
                           => n4261);
   U4775 : NAND2_X1 port map( A1 => n5322, A2 => fromRegsPortxREG_FILE_07xx29x,
                           ZN => n4260);
   U4776 : NAND4_X1 port map( A1 => n4263, A2 => n4262, A3 => n4261, A4 => 
                           n4260, ZN => n4267);
   U4777 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx29x,
                           ZN => n4265);
   U4778 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx29x, A2 => n5330,
                           ZN => n4264);
   U4779 : NAND2_X1 port map( A1 => n4265, A2 => n4264, ZN => n4266);
   U4780 : AOI21_X1 port map( B1 => n4267, B2 => n5334, A => n4266, ZN => n4268
                           );
   U4781 : NAND2_X1 port map( A1 => n4269, A2 => n4268, ZN => n7252);
   U4782 : INV_X1 port map( A => n7252, ZN => n7485);
   U4783 : OAI22_X1 port map( A1 => n5679, A2 => intadd_28xBx1x, B1 => n5676, 
                           B2 => n7485, ZN => n4270);
   U4784 : XOR2_X1 port map( A => n5146, B => n4270, Z => 
                           DP_OP_719J14_125_1055xn39);
   U4785 : NAND2_X1 port map( A1 => n5694, A2 => fromMemoryPortxLOADEDDATAx(28)
                           , ZN => n4271);
   U4786 : NAND2_X1 port map( A1 => n4504, A2 => n4271, ZN => add_x_26xBx28x);
   U4787 : INV_X1 port map( A => add_x_26xBx28x, ZN => intadd_28xBx0x);
   U4788 : CLKBUF_X1 port map( A => n5677, Z => n7364);
   U4789 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx28x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx28x, ZN
                           => n4275);
   U4790 : AOI22_X1 port map( A1 => n5282, A2 => fromRegsPortxREG_FILE_24xx28x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx28x, ZN
                           => n4274);
   U4791 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx28x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_27xx28x, ZN
                           => n4273);
   U4792 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx28x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx28x, ZN
                           => n4272);
   U4793 : NAND4_X1 port map( A1 => n4275, A2 => n4274, A3 => n4273, A4 => 
                           n4272, ZN => n4281);
   U4794 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx28x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx28x, ZN
                           => n4279);
   U4795 : AOI22_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx28x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_19xx28x, ZN
                           => n4278);
   U4796 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx28x,
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx28x, ZN
                           => n4277);
   U4797 : NAND2_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx28x,
                           ZN => n4276);
   U4798 : NAND4_X1 port map( A1 => n4279, A2 => n4278, A3 => n4277, A4 => 
                           n4276, ZN => n4280);
   U4799 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4281
                           , A => n4280, ZN => n4287);
   U4800 : AOI22_X1 port map( A1 => n5306, A2 => fromRegsPortxREG_FILE_13xx28x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx28x, ZN
                           => n4286);
   U4801 : CLKBUF_X1 port map( A => n5303, Z => n5129);
   U4802 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx28x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_11xx28x, ZN
                           => n4283);
   U4803 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx28x,
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx28x, ZN
                           => n4282);
   U4804 : NAND2_X1 port map( A1 => n4283, A2 => n4282, ZN => n4284);
   U4805 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx28x, B2 => n5129,
                           A => n4284, ZN => n4285);
   U4806 : OAI211_X1 port map( C1 => n4287, C2 => n7071, A => n4286, B => n4285
                           , ZN => n4288);
   U4807 : NAND2_X1 port map( A1 => n4288, A2 => n5316, ZN => n4298);
   U4808 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx28x,
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx28x, ZN
                           => n4292);
   U4809 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx28x,
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx28x, ZN
                           => n4291);
   U4810 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx28x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx28x, ZN
                           => n4290);
   U4811 : NAND2_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx28x,
                           ZN => n4289);
   U4812 : NAND4_X1 port map( A1 => n4292, A2 => n4291, A3 => n4290, A4 => 
                           n4289, ZN => n4296);
   U4813 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx28x,
                           ZN => n4294);
   U4814 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx28x, A2 => n5330,
                           ZN => n4293);
   U4815 : NAND2_X1 port map( A1 => n4294, A2 => n4293, ZN => n4295);
   U4816 : AOI21_X1 port map( B1 => n4296, B2 => n5334, A => n4295, ZN => n4297
                           );
   U4817 : NAND2_X1 port map( A1 => n4298, A2 => n4297, ZN => n7242);
   U4818 : INV_X1 port map( A => n7242, ZN => n7484);
   U4819 : OAI22_X1 port map( A1 => n5679, A2 => intadd_28xBx0x, B1 => n7364, 
                           B2 => n7484, ZN => n4299);
   U4820 : XOR2_X1 port map( A => n7550, B => n4299, Z => 
                           DP_OP_719J14_125_1055xn40);
   U4821 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx27x,
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_29xx27x, ZN
                           => n4303);
   U4822 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx27x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx27x, ZN
                           => n4302);
   U4823 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_26xx27x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_27xx27x, ZN
                           => n4301);
   U4824 : AOI22_X1 port map( A1 => n5282, A2 => fromRegsPortxREG_FILE_24xx27x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx27x, ZN
                           => n4300);
   U4825 : NAND4_X1 port map( A1 => n4303, A2 => n4302, A3 => n4301, A4 => 
                           n4300, ZN => n4309);
   U4826 : AOI22_X1 port map( A1 => n5295, A2 => fromRegsPortxREG_FILE_18xx27x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_19xx27x, ZN
                           => n4307);
   U4827 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx27x,
                           B1 => n5289, B2 => fromRegsPortxREG_FILE_22xx27x, ZN
                           => n4306);
   U4828 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx27x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx27x, ZN
                           => n4305);
   U4829 : NAND2_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx27x,
                           ZN => n4304);
   U4830 : NAND4_X1 port map( A1 => n4307, A2 => n4306, A3 => n4305, A4 => 
                           n4304, ZN => n4308);
   U4831 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4309
                           , A => n4308, ZN => n4315);
   U4832 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx27x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx27x, ZN
                           => n4314);
   U4833 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx27x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx27x, ZN
                           => n4311);
   U4834 : AOI22_X1 port map( A1 => n5305, A2 => fromRegsPortxREG_FILE_11xx27x,
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx27x, ZN
                           => n4310);
   U4835 : NAND2_X1 port map( A1 => n4311, A2 => n4310, ZN => n4312);
   U4836 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx27x, B2 => n5303,
                           A => n4312, ZN => n4313);
   U4837 : OAI211_X1 port map( C1 => n4315, C2 => n5314, A => n4314, B => n4313
                           , ZN => n4316);
   U4838 : NAND2_X1 port map( A1 => n4316, A2 => n5316, ZN => n4326);
   U4839 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx27x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx27x, ZN
                           => n4320);
   U4840 : AOI22_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx27x,
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx27x, ZN
                           => n4319);
   U4841 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx27x,
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx27x, ZN
                           => n4318);
   U4842 : NAND2_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx27x,
                           ZN => n4317);
   U4843 : NAND4_X1 port map( A1 => n4320, A2 => n4319, A3 => n4318, A4 => 
                           n4317, ZN => n4324);
   U4844 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx27x,
                           ZN => n4322);
   U4845 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx27x, A2 => n5330,
                           ZN => n4321);
   U4846 : NAND2_X1 port map( A1 => n4322, A2 => n4321, ZN => n4323);
   U4847 : AOI21_X1 port map( B1 => n4324, B2 => n5334, A => n4323, ZN => n4325
                           );
   U4848 : NAND2_X1 port map( A1 => n4326, A2 => n4325, ZN => n7183);
   U4849 : INV_X1 port map( A => n7183, ZN => n7483);
   U4850 : CLKBUF_X1 port map( A => n5674, Z => n5675);
   U4851 : INV_X1 port map( A => add_x_26xBx27x, ZN => n7168);
   U4852 : OAI22_X1 port map( A1 => n7483, A2 => n5678, B1 => n5675, B2 => 
                           n7168, ZN => n4327);
   U4853 : XOR2_X1 port map( A => n7550, B => n4327, Z => 
                           DP_OP_719J14_125_1055xn41);
   U4854 : NAND2_X1 port map( A1 => n5694, A2 => fromMemoryPortxLOADEDDATAx(26)
                           , ZN => n4328);
   U4855 : NAND2_X1 port map( A1 => n4504, A2 => n4328, ZN => add_x_26xBx26x);
   U4856 : INV_X1 port map( A => add_x_26xBx26x, ZN => n7126);
   U4857 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx26x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx26x, ZN
                           => n4332);
   U4858 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx26x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx26x, ZN
                           => n4331);
   U4859 : AOI22_X1 port map( A1 => n5282, A2 => fromRegsPortxREG_FILE_24xx26x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_27xx26x, ZN
                           => n4330);
   U4860 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx26x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx26x, ZN
                           => n4329);
   U4861 : NAND4_X1 port map( A1 => n4332, A2 => n4331, A3 => n4330, A4 => 
                           n4329, ZN => n4338);
   U4862 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx26x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_19xx26x, ZN
                           => n4336);
   U4863 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx26x,
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_23xx26x, ZN
                           => n4335);
   U4864 : AOI22_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx26x,
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx26x, ZN
                           => n4334);
   U4865 : NAND2_X1 port map( A1 => n5294, A2 => fromRegsPortxREG_FILE_17xx26x,
                           ZN => n4333);
   U4866 : NAND4_X1 port map( A1 => n4336, A2 => n4335, A3 => n4334, A4 => 
                           n4333, ZN => n4337);
   U4867 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4338
                           , A => n4337, ZN => n4344);
   U4868 : AOI22_X1 port map( A1 => n5305, A2 => fromRegsPortxREG_FILE_11xx26x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx26x, ZN
                           => n4343);
   U4869 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx26x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx26x, ZN
                           => n4340);
   U4870 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx26x,
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx26x, ZN
                           => n4339);
   U4871 : NAND2_X1 port map( A1 => n4340, A2 => n4339, ZN => n4341);
   U4872 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx26x, B2 => n5303,
                           A => n4341, ZN => n4342);
   U4873 : OAI211_X1 port map( C1 => n4344, C2 => n5314, A => n4343, B => n4342
                           , ZN => n4345);
   U4874 : NAND2_X1 port map( A1 => n4345, A2 => n5316, ZN => n4355);
   U4875 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx26x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx26x, ZN
                           => n4349);
   U4876 : AOI22_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx26x,
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx26x, ZN
                           => n4348);
   U4877 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx26x,
                           B1 => n5318, B2 => fromRegsPortxREG_FILE_03xx26x, ZN
                           => n4347);
   U4878 : NAND2_X1 port map( A1 => n5323, A2 => fromRegsPortxREG_FILE_05xx26x,
                           ZN => n4346);
   U4879 : NAND4_X1 port map( A1 => n4349, A2 => n4348, A3 => n4347, A4 => 
                           n4346, ZN => n4353);
   U4880 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx26x,
                           ZN => n4351);
   U4881 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx26x, A2 => n5330,
                           ZN => n4350);
   U4882 : NAND2_X1 port map( A1 => n4351, A2 => n4350, ZN => n4352);
   U4883 : AOI21_X1 port map( B1 => n4353, B2 => n5334, A => n4352, ZN => n4354
                           );
   U4884 : NAND2_X1 port map( A1 => n4355, A2 => n4354, ZN => n7120);
   U4885 : INV_X1 port map( A => n7120, ZN => n7482);
   U4886 : OAI22_X1 port map( A1 => n5679, A2 => n7126, B1 => n5676, B2 => 
                           n7482, ZN => n4356);
   U4887 : XOR2_X1 port map( A => n5146, B => n4356, Z => 
                           DP_OP_719J14_125_1055xn42);
   U4888 : NAND2_X1 port map( A1 => n5694, A2 => fromMemoryPortxLOADEDDATAx(25)
                           , ZN => n4357);
   U4889 : NAND2_X1 port map( A1 => n4504, A2 => n4357, ZN => add_x_26xBx25x);
   U4890 : INV_X1 port map( A => add_x_26xBx25x, ZN => n7080);
   U4891 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx25x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx25x, ZN
                           => n4361);
   U4892 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx25x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_24xx25x, ZN
                           => n4360);
   U4893 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx25x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx25x, ZN
                           => n4359);
   U4894 : AOI22_X1 port map( A1 => n5281, A2 => fromRegsPortxREG_FILE_27xx25x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx25x, ZN
                           => n4358);
   U4895 : NAND4_X1 port map( A1 => n4361, A2 => n4360, A3 => n4359, A4 => 
                           n4358, ZN => n4367);
   U4896 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx25x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_19xx25x, ZN
                           => n4365);
   U4897 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx25x,
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx25x, ZN
                           => n4364);
   U4898 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx25x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx25x, ZN
                           => n4363);
   U4899 : NAND2_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_22xx25x,
                           ZN => n4362);
   U4900 : NAND4_X1 port map( A1 => n4365, A2 => n4364, A3 => n4363, A4 => 
                           n4362, ZN => n4366);
   U4901 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4367
                           , A => n4366, ZN => n4373);
   U4902 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx25x,
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx25x, ZN
                           => n4372);
   U4903 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx25x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx25x, ZN
                           => n4369);
   U4904 : AOI22_X1 port map( A1 => n5305, A2 => fromRegsPortxREG_FILE_11xx25x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx25x, ZN
                           => n4368);
   U4905 : NAND2_X1 port map( A1 => n4369, A2 => n4368, ZN => n4370);
   U4906 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx25x, B2 => n5303,
                           A => n4370, ZN => n4371);
   U4907 : OAI211_X1 port map( C1 => n4373, C2 => n5314, A => n4372, B => n4371
                           , ZN => n4374);
   U4908 : NAND2_X1 port map( A1 => n4374, A2 => n5316, ZN => n4384);
   U4909 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx25x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_06xx25x, ZN
                           => n4378);
   U4910 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx25x,
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx25x, ZN
                           => n4377);
   U4911 : AOI22_X1 port map( A1 => n5323, A2 => fromRegsPortxREG_FILE_05xx25x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx25x, ZN
                           => n4376);
   U4912 : NAND2_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx25x,
                           ZN => n4375);
   U4913 : NAND4_X1 port map( A1 => n4378, A2 => n4377, A3 => n4376, A4 => 
                           n4375, ZN => n4382);
   U4914 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx25x,
                           ZN => n4380);
   U4915 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx25x, A2 => n5330,
                           ZN => n4379);
   U4916 : NAND2_X1 port map( A1 => n4380, A2 => n4379, ZN => n4381);
   U4917 : AOI21_X1 port map( B1 => n4382, B2 => n5334, A => n4381, ZN => n4383
                           );
   U4918 : NAND2_X1 port map( A1 => n4384, A2 => n4383, ZN => n7097);
   U4919 : INV_X1 port map( A => n7097, ZN => n7481);
   U4920 : OAI22_X1 port map( A1 => n5679, A2 => n7080, B1 => n7364, B2 => 
                           n7481, ZN => n4385);
   U4921 : XOR2_X1 port map( A => n7550, B => n4385, Z => 
                           DP_OP_719J14_125_1055xn43);
   U4922 : NAND2_X1 port map( A1 => n5694, A2 => fromMemoryPortxLOADEDDATAx(24)
                           , ZN => n4386);
   U4923 : NAND2_X1 port map( A1 => n4504, A2 => n4386, ZN => add_x_26xBx24x);
   U4924 : INV_X1 port map( A => add_x_26xBx24x, ZN => intadd_26xBx7x);
   U4925 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_26xx24x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_24xx24x, ZN
                           => n4390);
   U4926 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx24x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx24x, ZN
                           => n4389);
   U4927 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx24x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_27xx24x, ZN
                           => n4388);
   U4928 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx24x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx24x, ZN
                           => n4387);
   U4929 : NAND4_X1 port map( A1 => n4390, A2 => n4389, A3 => n4388, A4 => 
                           n4387, ZN => n4396);
   U4930 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx24x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx24x, ZN
                           => n4394);
   U4931 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx24x,
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_23xx24x, ZN
                           => n4393);
   U4932 : AOI22_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_22xx24x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_19xx24x, ZN
                           => n4392);
   U4933 : NAND2_X1 port map( A1 => n5295, A2 => fromRegsPortxREG_FILE_18xx24x,
                           ZN => n4391);
   U4934 : NAND4_X1 port map( A1 => n4394, A2 => n4393, A3 => n4392, A4 => 
                           n4391, ZN => n4395);
   U4935 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4396
                           , A => n4395, ZN => n4402);
   U4936 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx24x,
                           B1 => n5303, B2 => fromRegsPortxREG_FILE_12xx24x, ZN
                           => n4401);
   U4937 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx24x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx24x, ZN
                           => n4398);
   U4938 : AOI22_X1 port map( A1 => n5311, A2 => fromRegsPortxREG_FILE_16xx24x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx24x, ZN
                           => n4397);
   U4939 : NAND2_X1 port map( A1 => n4398, A2 => n4397, ZN => n4399);
   U4940 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_11xx24x, B2 => n5305,
                           A => n4399, ZN => n4400);
   U4941 : OAI211_X1 port map( C1 => n4402, C2 => n5314, A => n4401, B => n4400
                           , ZN => n4403);
   U4942 : NAND2_X1 port map( A1 => n4403, A2 => n5316, ZN => n4413);
   U4943 : AOI22_X1 port map( A1 => n5324, A2 => fromRegsPortxREG_FILE_08xx24x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx24x, ZN
                           => n4407);
   U4944 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx24x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_06xx24x, ZN
                           => n4406);
   U4945 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx24x,
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx24x, ZN
                           => n4405);
   U4946 : NAND2_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx24x,
                           ZN => n4404);
   U4947 : NAND4_X1 port map( A1 => n4407, A2 => n4406, A3 => n4405, A4 => 
                           n4404, ZN => n4411);
   U4948 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx24x,
                           ZN => n4409);
   U4949 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx24x, A2 => n5330,
                           ZN => n4408);
   U4950 : NAND2_X1 port map( A1 => n4409, A2 => n4408, ZN => n4410);
   U4951 : AOI21_X1 port map( B1 => n4411, B2 => n5334, A => n4410, ZN => n4412
                           );
   U4952 : NAND2_X1 port map( A1 => n4413, A2 => n4412, ZN => n7053);
   U4953 : INV_X1 port map( A => n7053, ZN => n7480);
   U4954 : OAI22_X1 port map( A1 => n7480, A2 => n5678, B1 => n5675, B2 => 
                           intadd_26xBx7x, ZN => n4414);
   U4955 : XOR2_X1 port map( A => n7550, B => n4414, Z => 
                           DP_OP_719J14_125_1055xn44);
   U4956 : NAND2_X1 port map( A1 => n4504, A2 => n7033, ZN => n4415);
   U4957 : AND2_X1 port map( A1 => n4445, A2 => n4415, ZN => add_x_26xBx23x);
   U4958 : INV_X1 port map( A => add_x_26xBx23x, ZN => intadd_26xBx6x);
   U4959 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx23x,
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_29xx23x, ZN
                           => n4419);
   U4960 : AOI22_X1 port map( A1 => n5282, A2 => fromRegsPortxREG_FILE_24xx23x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_27xx23x, ZN
                           => n4418);
   U4961 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx23x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx23x, ZN
                           => n4417);
   U4962 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_26xx23x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx23x, ZN
                           => n4416);
   U4963 : NAND4_X1 port map( A1 => n4419, A2 => n4418, A3 => n4417, A4 => 
                           n4416, ZN => n4425);
   U4964 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx23x,
                           B1 => n5019, B2 => fromRegsPortxREG_FILE_23xx23x, ZN
                           => n4423);
   U4965 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx23x,
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_22xx23x, ZN
                           => n4422);
   U4966 : AOI22_X1 port map( A1 => n5295, A2 => fromRegsPortxREG_FILE_18xx23x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx23x, ZN
                           => n4421);
   U4967 : NAND2_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_19xx23x,
                           ZN => n4420);
   U4968 : NAND4_X1 port map( A1 => n4423, A2 => n4422, A3 => n4421, A4 => 
                           n4420, ZN => n4424);
   U4969 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4425
                           , A => n4424, ZN => n4431);
   U4970 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx23x,
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx23x, ZN
                           => n4430);
   U4971 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx23x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx23x, ZN
                           => n4427);
   U4972 : AOI22_X1 port map( A1 => n5305, A2 => fromRegsPortxREG_FILE_11xx23x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx23x, ZN
                           => n4426);
   U4973 : NAND2_X1 port map( A1 => n4427, A2 => n4426, ZN => n4428);
   U4974 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx23x, B2 => n5129,
                           A => n4428, ZN => n4429);
   U4975 : OAI211_X1 port map( C1 => n4431, C2 => n7071, A => n4430, B => n4429
                           , ZN => n4432);
   U4976 : NAND2_X1 port map( A1 => n4432, A2 => n5316, ZN => n4442);
   U4977 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx23x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_06xx23x, ZN
                           => n4436);
   U4978 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx23x,
                           B1 => n4903, B2 => fromRegsPortxREG_FILE_05xx23x, ZN
                           => n4435);
   U4979 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx23x,
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx23x, ZN
                           => n4434);
   U4980 : NAND2_X1 port map( A1 => n5322, A2 => fromRegsPortxREG_FILE_07xx23x,
                           ZN => n4433);
   U4981 : NAND4_X1 port map( A1 => n4436, A2 => n4435, A3 => n4434, A4 => 
                           n4433, ZN => n4440);
   U4982 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx23x,
                           ZN => n4438);
   U4983 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx23x, A2 => n5330,
                           ZN => n4437);
   U4984 : NAND2_X1 port map( A1 => n4438, A2 => n4437, ZN => n4439);
   U4985 : AOI21_X1 port map( B1 => n4440, B2 => n5334, A => n4439, ZN => n4441
                           );
   U4986 : NAND2_X1 port map( A1 => n4442, A2 => n4441, ZN => n7009);
   U4987 : INV_X1 port map( A => n7009, ZN => n7479);
   U4988 : OAI22_X1 port map( A1 => n7479, A2 => n5678, B1 => n5675, B2 => 
                           intadd_26xBx6x, ZN => n4443);
   U4989 : XOR2_X1 port map( A => n5146, B => n4443, Z => 
                           DP_OP_719J14_125_1055xn45);
   U4990 : NAND2_X1 port map( A1 => n4504, A2 => n6995, ZN => n4444);
   U4991 : AND2_X1 port map( A1 => n4445, A2 => n4444, ZN => add_x_26xBx22x);
   U4992 : INV_X1 port map( A => add_x_26xBx22x, ZN => intadd_26xBx5x);
   U4993 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_26xx22x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_24xx22x, ZN
                           => n4449);
   U4994 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx22x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_27xx22x, ZN
                           => n4448);
   U4995 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx22x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx22x, ZN
                           => n4447);
   U4996 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx22x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx22x, ZN
                           => n4446);
   U4997 : NAND4_X1 port map( A1 => n4449, A2 => n4448, A3 => n4447, A4 => 
                           n4446, ZN => n4455);
   U4998 : AOI22_X1 port map( A1 => n5295, A2 => fromRegsPortxREG_FILE_18xx22x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_19xx22x, ZN
                           => n4453);
   U4999 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx22x,
                           B1 => n5290, B2 => fromRegsPortxREG_FILE_21xx22x, ZN
                           => n4452);
   U5000 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx22x,
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_22xx22x, ZN
                           => n4451);
   U5001 : NAND2_X1 port map( A1 => n5294, A2 => fromRegsPortxREG_FILE_17xx22x,
                           ZN => n4450);
   U5002 : NAND4_X1 port map( A1 => n4453, A2 => n4452, A3 => n4451, A4 => 
                           n4450, ZN => n4454);
   U5003 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4455
                           , A => n4454, ZN => n4461);
   U5004 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx22x,
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx22x, ZN
                           => n4460);
   U5005 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx22x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_11xx22x, ZN
                           => n4457);
   U5006 : AOI22_X1 port map( A1 => n5306, A2 => fromRegsPortxREG_FILE_13xx22x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx22x, ZN
                           => n4456);
   U5007 : NAND2_X1 port map( A1 => n4457, A2 => n4456, ZN => n4458);
   U5008 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx22x, B2 => n5129,
                           A => n4458, ZN => n4459);
   U5009 : OAI211_X1 port map( C1 => n4461, C2 => n7071, A => n4460, B => n4459
                           , ZN => n4462);
   U5010 : CLKBUF_X1 port map( A => n5316, Z => n5133);
   U5011 : NAND2_X1 port map( A1 => n4462, A2 => n5133, ZN => n4472);
   U5012 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx22x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx22x, ZN
                           => n4466);
   U5013 : AOI22_X1 port map( A1 => n4932, A2 => fromRegsPortxREG_FILE_08xx22x,
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx22x, ZN
                           => n4465);
   U5014 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx22x,
                           B1 => n5036, B2 => fromRegsPortxREG_FILE_03xx22x, ZN
                           => n4464);
   U5015 : NAND2_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx22x,
                           ZN => n4463);
   U5016 : NAND4_X1 port map( A1 => n4466, A2 => n4465, A3 => n4464, A4 => 
                           n4463, ZN => n4470);
   U5017 : NAND2_X1 port map( A1 => n4760, A2 => fromRegsPortxREG_FILE_02xx22x,
                           ZN => n4468);
   U5018 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx22x, A2 => n5330,
                           ZN => n4467);
   U5019 : NAND2_X1 port map( A1 => n4468, A2 => n4467, ZN => n4469);
   U5020 : AOI21_X1 port map( B1 => n4470, B2 => n5334, A => n4469, ZN => n4471
                           );
   U5021 : NAND2_X1 port map( A1 => n4472, A2 => n4471, ZN => n6958);
   U5022 : INV_X1 port map( A => n6958, ZN => n7478);
   U5023 : OAI22_X1 port map( A1 => n5674, A2 => intadd_26xBx5x, B1 => n5676, 
                           B2 => n7478, ZN => n4473);
   U5024 : XOR2_X1 port map( A => n5146, B => n4473, Z => 
                           DP_OP_719J14_125_1055xn46);
   U5025 : NAND2_X1 port map( A1 => n5694, A2 => fromMemoryPortxLOADEDDATAx(21)
                           , ZN => n4474);
   U5026 : NAND2_X1 port map( A1 => n4504, A2 => n4474, ZN => add_x_26xBx21x);
   U5027 : INV_X1 port map( A => add_x_26xBx21x, ZN => intadd_26xBx4x);
   U5028 : AOI22_X1 port map( A1 => n5013, A2 => fromRegsPortxREG_FILE_24xx21x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx21x, ZN
                           => n4478);
   U5029 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx21x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx21x, ZN
                           => n4477);
   U5030 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx21x,
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_29xx21x, ZN
                           => n4476);
   U5031 : AOI22_X1 port map( A1 => n5281, A2 => fromRegsPortxREG_FILE_27xx21x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx21x, ZN
                           => n4475);
   U5032 : NAND4_X1 port map( A1 => n4478, A2 => n4477, A3 => n4476, A4 => 
                           n4475, ZN => n4484);
   U5033 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx21x,
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_22xx21x, ZN
                           => n4482);
   U5034 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx21x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_19xx21x, ZN
                           => n4481);
   U5035 : AOI22_X1 port map( A1 => n4986, A2 => fromRegsPortxREG_FILE_18xx21x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx21x, ZN
                           => n4480);
   U5036 : NAND2_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx21x,
                           ZN => n4479);
   U5037 : NAND4_X1 port map( A1 => n4482, A2 => n4481, A3 => n4480, A4 => 
                           n4479, ZN => n4483);
   U5038 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4484
                           , A => n4483, ZN => n4490);
   U5039 : AOI22_X1 port map( A1 => n5305, A2 => fromRegsPortxREG_FILE_11xx21x,
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx21x, ZN
                           => n4489);
   U5040 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx21x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx21x, ZN
                           => n4486);
   U5041 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_12xx21x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx21x, ZN
                           => n4485);
   U5042 : NAND2_X1 port map( A1 => n4486, A2 => n4485, ZN => n4487);
   U5043 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx21x, B2 => n5302,
                           A => n4487, ZN => n4488);
   U5044 : OAI211_X1 port map( C1 => n4490, C2 => n7071, A => n4489, B => n4488
                           , ZN => n4491);
   U5045 : NAND2_X1 port map( A1 => n4491, A2 => n5133, ZN => n4501);
   U5046 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx21x,
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_06xx21x, ZN
                           => n4495);
   U5047 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx21x,
                           B1 => n4903, B2 => fromRegsPortxREG_FILE_05xx21x, ZN
                           => n4494);
   U5048 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx21x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx21x, ZN
                           => n4493);
   U5049 : NAND2_X1 port map( A1 => n4932, A2 => fromRegsPortxREG_FILE_08xx21x,
                           ZN => n4492);
   U5050 : NAND4_X1 port map( A1 => n4495, A2 => n4494, A3 => n4493, A4 => 
                           n4492, ZN => n4499);
   U5051 : NAND2_X1 port map( A1 => n4760, A2 => fromRegsPortxREG_FILE_02xx21x,
                           ZN => n4497);
   U5052 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx21x, A2 => n5330,
                           ZN => n4496);
   U5053 : NAND2_X1 port map( A1 => n4497, A2 => n4496, ZN => n4498);
   U5054 : AOI21_X1 port map( B1 => n4499, B2 => n5334, A => n4498, ZN => n4500
                           );
   U5055 : NAND2_X1 port map( A1 => n4501, A2 => n4500, ZN => n5720);
   U5056 : INV_X1 port map( A => n5720, ZN => n7477);
   U5057 : OAI22_X1 port map( A1 => n5674, A2 => intadd_26xBx4x, B1 => n5677, 
                           B2 => n7477, ZN => n4502);
   U5058 : XOR2_X1 port map( A => n5146, B => n4502, Z => 
                           DP_OP_719J14_125_1055xn47);
   U5059 : NAND2_X1 port map( A1 => n5694, A2 => fromMemoryPortxLOADEDDATAx(20)
                           , ZN => n4503);
   U5060 : NAND2_X1 port map( A1 => n4504, A2 => n4503, ZN => add_x_26xBx20x);
   U5061 : INV_X1 port map( A => add_x_26xBx20x, ZN => intadd_26xBx3x);
   U5062 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx20x,
                           B1 => n5013, B2 => fromRegsPortxREG_FILE_24xx20x, ZN
                           => n4508);
   U5063 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx20x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx20x, ZN
                           => n4507);
   U5064 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx20x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_27xx20x, ZN
                           => n4506);
   U5065 : AOI22_X1 port map( A1 => n5284, A2 => fromRegsPortxREG_FILE_31xx20x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx20x, ZN
                           => n4505);
   U5066 : NAND4_X1 port map( A1 => n4508, A2 => n4507, A3 => n4506, A4 => 
                           n4505, ZN => n4514);
   U5067 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx20x,
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_22xx20x, ZN
                           => n4512);
   U5068 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx20x,
                           B1 => n4986, B2 => fromRegsPortxREG_FILE_18xx20x, ZN
                           => n4511);
   U5069 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx20x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_19xx20x, ZN
                           => n4510);
   U5070 : NAND2_X1 port map( A1 => n5294, A2 => fromRegsPortxREG_FILE_17xx20x,
                           ZN => n4509);
   U5071 : NAND4_X1 port map( A1 => n4512, A2 => n4511, A3 => n4510, A4 => 
                           n4509, ZN => n4513);
   U5072 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4514
                           , A => n4513, ZN => n4520);
   U5073 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx20x,
                           B1 => n4957, B2 => fromRegsPortxREG_FILE_16xx20x, ZN
                           => n4519);
   U5074 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx20x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx20x, ZN
                           => n4516);
   U5075 : AOI22_X1 port map( A1 => n5305, A2 => fromRegsPortxREG_FILE_11xx20x,
                           B1 => n5306, B2 => fromRegsPortxREG_FILE_13xx20x, ZN
                           => n4515);
   U5076 : NAND2_X1 port map( A1 => n4516, A2 => n4515, ZN => n4517);
   U5077 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx20x, B2 => n5129,
                           A => n4517, ZN => n4518);
   U5078 : OAI211_X1 port map( C1 => n4520, C2 => n7071, A => n4519, B => n4518
                           , ZN => n4521);
   U5079 : NAND2_X1 port map( A1 => n4521, A2 => n5133, ZN => n4531);
   U5080 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx20x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx20x, ZN
                           => n4525);
   U5081 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx20x,
                           B1 => n4903, B2 => fromRegsPortxREG_FILE_05xx20x, ZN
                           => n4524);
   U5082 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx20x,
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx20x, ZN
                           => n4523);
   U5083 : NAND2_X1 port map( A1 => n5034, A2 => fromRegsPortxREG_FILE_06xx20x,
                           ZN => n4522);
   U5084 : NAND4_X1 port map( A1 => n4525, A2 => n4524, A3 => n4523, A4 => 
                           n4522, ZN => n4529);
   U5085 : NAND2_X1 port map( A1 => n4760, A2 => fromRegsPortxREG_FILE_02xx20x,
                           ZN => n4527);
   U5086 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx20x, A2 => n5330,
                           ZN => n4526);
   U5087 : NAND2_X1 port map( A1 => n4527, A2 => n4526, ZN => n4528);
   U5088 : AOI21_X1 port map( B1 => n4529, B2 => n5334, A => n4528, ZN => n4530
                           );
   U5089 : NAND2_X1 port map( A1 => n4531, A2 => n4530, ZN => n6933);
   U5090 : INV_X1 port map( A => n6933, ZN => n7476);
   U5091 : OAI22_X1 port map( A1 => n5674, A2 => intadd_26xBx3x, B1 => n7364, 
                           B2 => n7476, ZN => n4532);
   U5092 : XOR2_X1 port map( A => n5146, B => n4532, Z => 
                           DP_OP_719J14_125_1055xn48);
   U5093 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(31), A2 => n4533,
                           ZN => n4769);
   U5094 : AOI21_X1 port map( B1 => n4768, B2 => fromMemoryPortxLOADEDDATAx(31)
                           , A => n4769, ZN => n5653);
   U5095 : NAND2_X1 port map( A1 => n7445, A2 => fromMemoryPortxLOADEDDATAx(3),
                           ZN => n5642);
   U5096 : NAND2_X1 port map( A1 => n5642, A2 => n4534, ZN => n5651);
   U5097 : NAND2_X1 port map( A1 => n5651, A2 => fromMemoryPortxLOADEDDATAx(19)
                           , ZN => n4535);
   U5098 : NAND2_X1 port map( A1 => n5653, A2 => n4535, ZN => add_x_26xBx19x);
   U5099 : INV_X1 port map( A => add_x_26xBx19x, ZN => intadd_26xBx2x);
   U5100 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_26xx19x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_24xx19x, ZN
                           => n4539);
   U5101 : AOI22_X1 port map( A1 => n4945, A2 => fromRegsPortxREG_FILE_29xx19x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_27xx19x, ZN
                           => n4538);
   U5102 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx19x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx19x, ZN
                           => n4537);
   U5103 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx19x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx19x, ZN
                           => n4536);
   U5104 : NAND4_X1 port map( A1 => n4539, A2 => n4538, A3 => n4537, A4 => 
                           n4536, ZN => n4545);
   U5105 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx19x,
                           B1 => n5290, B2 => fromRegsPortxREG_FILE_21xx19x, ZN
                           => n4543);
   U5106 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx19x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx19x, ZN
                           => n4542);
   U5107 : AOI22_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx19x,
                           B1 => n4986, B2 => fromRegsPortxREG_FILE_18xx19x, ZN
                           => n4541);
   U5108 : NAND2_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_19xx19x,
                           ZN => n4540);
   U5109 : NAND4_X1 port map( A1 => n4543, A2 => n4542, A3 => n4541, A4 => 
                           n4540, ZN => n4544);
   U5110 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4545
                           , A => n4544, ZN => n4551);
   U5111 : AOI22_X1 port map( A1 => n5306, A2 => fromRegsPortxREG_FILE_13xx19x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx19x, ZN
                           => n4550);
   U5112 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx19x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_11xx19x, ZN
                           => n4547);
   U5113 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_12xx19x,
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx19x, ZN
                           => n4546);
   U5114 : NAND2_X1 port map( A1 => n4547, A2 => n4546, ZN => n4548);
   U5115 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx19x, B2 => n5302,
                           A => n4548, ZN => n4549);
   U5116 : OAI211_X1 port map( C1 => n4551, C2 => n7071, A => n4550, B => n4549
                           , ZN => n4552);
   U5117 : NAND2_X1 port map( A1 => n4552, A2 => n5133, ZN => n4562);
   U5118 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx19x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx19x, ZN
                           => n4556);
   U5119 : AOI22_X1 port map( A1 => n5034, A2 => fromRegsPortxREG_FILE_06xx19x,
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx19x, ZN
                           => n4555);
   U5120 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx19x,
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx19x, ZN
                           => n4554);
   U5121 : NAND2_X1 port map( A1 => n5036, A2 => fromRegsPortxREG_FILE_03xx19x,
                           ZN => n4553);
   U5122 : NAND4_X1 port map( A1 => n4556, A2 => n4555, A3 => n4554, A4 => 
                           n4553, ZN => n4560);
   U5123 : NAND2_X1 port map( A1 => n4760, A2 => fromRegsPortxREG_FILE_02xx19x,
                           ZN => n4558);
   U5124 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx19x, A2 => n5330,
                           ZN => n4557);
   U5125 : NAND2_X1 port map( A1 => n4558, A2 => n4557, ZN => n4559);
   U5126 : AOI21_X1 port map( B1 => n4560, B2 => n5334, A => n4559, ZN => n4561
                           );
   U5127 : NAND2_X1 port map( A1 => n4562, A2 => n4561, ZN => n6888);
   U5128 : INV_X1 port map( A => n6888, ZN => n7475);
   U5129 : OAI22_X1 port map( A1 => n5674, A2 => intadd_26xBx2x, B1 => n7364, 
                           B2 => n7475, ZN => n4563);
   U5130 : XOR2_X1 port map( A => n7550, B => n4563, Z => 
                           DP_OP_719J14_125_1055xn49);
   U5131 : NAND2_X1 port map( A1 => n5651, A2 => fromMemoryPortxLOADEDDATAx(18)
                           , ZN => n4564);
   U5132 : NAND2_X1 port map( A1 => n5653, A2 => n4564, ZN => add_x_26xBx18x);
   U5133 : INV_X1 port map( A => add_x_26xBx18x, ZN => intadd_26xBx1x);
   U5134 : AOI22_X1 port map( A1 => n5013, A2 => fromRegsPortxREG_FILE_24xx18x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx18x, ZN
                           => n4568);
   U5135 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx18x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx18x, ZN
                           => n4567);
   U5136 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx18x,
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_27xx18x, ZN
                           => n4566);
   U5137 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx18x,
                           B1 => n4946, B2 => fromRegsPortxREG_FILE_31xx18x, ZN
                           => n4565);
   U5138 : NAND4_X1 port map( A1 => n4568, A2 => n4567, A3 => n4566, A4 => 
                           n4565, ZN => n4574);
   U5139 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx18x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx18x, ZN
                           => n4572);
   U5140 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx18x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_19xx18x, ZN
                           => n4571);
   U5141 : AOI22_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx18x,
                           B1 => n4986, B2 => fromRegsPortxREG_FILE_18xx18x, ZN
                           => n4570);
   U5142 : NAND2_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx18x,
                           ZN => n4569);
   U5143 : NAND4_X1 port map( A1 => n4572, A2 => n4571, A3 => n4570, A4 => 
                           n4569, ZN => n4573);
   U5144 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4574
                           , A => n4573, ZN => n4580);
   U5145 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_12xx18x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx18x, ZN
                           => n4579);
   U5146 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx18x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_11xx18x, ZN
                           => n4576);
   U5147 : AOI22_X1 port map( A1 => n4957, A2 => fromRegsPortxREG_FILE_16xx18x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx18x, ZN
                           => n4575);
   U5148 : NAND2_X1 port map( A1 => n4576, A2 => n4575, ZN => n4577);
   U5149 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx18x, B2 => n5060,
                           A => n4577, ZN => n4578);
   U5150 : OAI211_X1 port map( C1 => n4580, C2 => n7071, A => n4579, B => n4578
                           , ZN => n4581);
   U5151 : NAND2_X1 port map( A1 => n4581, A2 => n5133, ZN => n4591);
   U5152 : AOI22_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx18x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx18x, ZN
                           => n4585);
   U5153 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx18x,
                           B1 => n4932, B2 => fromRegsPortxREG_FILE_08xx18x, ZN
                           => n4584);
   U5154 : AOI22_X1 port map( A1 => n5035, A2 => fromRegsPortxREG_FILE_09xx18x,
                           B1 => n5036, B2 => fromRegsPortxREG_FILE_03xx18x, ZN
                           => n4583);
   U5155 : NAND2_X1 port map( A1 => n4903, A2 => fromRegsPortxREG_FILE_05xx18x,
                           ZN => n4582);
   U5156 : NAND4_X1 port map( A1 => n4585, A2 => n4584, A3 => n4583, A4 => 
                           n4582, ZN => n4589);
   U5157 : NAND2_X1 port map( A1 => n4760, A2 => fromRegsPortxREG_FILE_02xx18x,
                           ZN => n4587);
   U5158 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx18x, A2 => n5330,
                           ZN => n4586);
   U5159 : NAND2_X1 port map( A1 => n4587, A2 => n4586, ZN => n4588);
   U5160 : AOI21_X1 port map( B1 => n4589, B2 => n5334, A => n4588, ZN => n4590
                           );
   U5161 : NAND2_X1 port map( A1 => n4591, A2 => n4590, ZN => n6861);
   U5162 : INV_X1 port map( A => n6861, ZN => n7474);
   U5163 : OAI22_X1 port map( A1 => n7474, A2 => n5676, B1 => n5675, B2 => 
                           intadd_26xBx1x, ZN => n4592);
   U5164 : XOR2_X1 port map( A => n5146, B => n4592, Z => 
                           DP_OP_719J14_125_1055xn50);
   U5165 : NAND2_X1 port map( A1 => n5651, A2 => fromMemoryPortxLOADEDDATAx(17)
                           , ZN => n4593);
   U5166 : NAND2_X1 port map( A1 => n5653, A2 => n4593, ZN => add_x_26xBx17x);
   U5167 : INV_X1 port map( A => add_x_26xBx17x, ZN => intadd_26xBx0x);
   U5168 : AOI22_X1 port map( A1 => n4980, A2 => fromRegsPortxREG_FILE_26xx17x,
                           B1 => n5013, B2 => fromRegsPortxREG_FILE_24xx17x, ZN
                           => n4597);
   U5169 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx17x,
                           B1 => n5012, B2 => fromRegsPortxREG_FILE_27xx17x, ZN
                           => n4596);
   U5170 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx17x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx17x, ZN
                           => n4595);
   U5171 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx17x,
                           B1 => n4946, B2 => fromRegsPortxREG_FILE_31xx17x, ZN
                           => n4594);
   U5172 : NAND4_X1 port map( A1 => n4597, A2 => n4596, A3 => n4595, A4 => 
                           n4594, ZN => n4603);
   U5173 : AOI22_X1 port map( A1 => n4986, A2 => fromRegsPortxREG_FILE_18xx17x,
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_19xx17x, ZN
                           => n4601);
   U5174 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx17x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx17x, ZN
                           => n4600);
   U5175 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx17x,
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_22xx17x, ZN
                           => n4599);
   U5176 : NAND2_X1 port map( A1 => n4985, A2 => fromRegsPortxREG_FILE_20xx17x,
                           ZN => n4598);
   U5177 : NAND4_X1 port map( A1 => n4601, A2 => n4600, A3 => n4599, A4 => 
                           n4598, ZN => n4602);
   U5178 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4603
                           , A => n4602, ZN => n4609);
   U5179 : AOI22_X1 port map( A1 => n5306, A2 => fromRegsPortxREG_FILE_13xx17x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx17x, ZN
                           => n4608);
   U5180 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx17x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_11xx17x, ZN
                           => n4605);
   U5181 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_12xx17x,
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx17x, ZN
                           => n4604);
   U5182 : NAND2_X1 port map( A1 => n4605, A2 => n4604, ZN => n4606);
   U5183 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx17x, B2 => n5060,
                           A => n4606, ZN => n4607);
   U5184 : OAI211_X1 port map( C1 => n4609, C2 => n5314, A => n4608, B => n4607
                           , ZN => n4610);
   U5185 : NAND2_X1 port map( A1 => n4610, A2 => n5133, ZN => n4620);
   U5186 : AOI22_X1 port map( A1 => n4932, A2 => fromRegsPortxREG_FILE_08xx17x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx17x, ZN
                           => n4614);
   U5187 : AOI22_X1 port map( A1 => n5035, A2 => fromRegsPortxREG_FILE_09xx17x,
                           B1 => n5034, B2 => fromRegsPortxREG_FILE_06xx17x, ZN
                           => n4613);
   U5188 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx17x,
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx17x, ZN
                           => n4612);
   U5189 : NAND2_X1 port map( A1 => n4965, A2 => fromRegsPortxREG_FILE_04xx17x,
                           ZN => n4611);
   U5190 : NAND4_X1 port map( A1 => n4614, A2 => n4613, A3 => n4612, A4 => 
                           n4611, ZN => n4618);
   U5191 : NAND2_X1 port map( A1 => n4760, A2 => fromRegsPortxREG_FILE_02xx17x,
                           ZN => n4616);
   U5192 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx17x, A2 => n5330,
                           ZN => n4615);
   U5193 : NAND2_X1 port map( A1 => n4616, A2 => n4615, ZN => n4617);
   U5194 : AOI21_X1 port map( B1 => n4618, B2 => n5334, A => n4617, ZN => n4619
                           );
   U5195 : NAND2_X1 port map( A1 => n4620, A2 => n4619, ZN => n6806);
   U5196 : INV_X1 port map( A => n6806, ZN => n7473);
   U5197 : OAI22_X1 port map( A1 => n5679, A2 => intadd_26xBx0x, B1 => n7364, 
                           B2 => n7473, ZN => n4621);
   U5198 : XOR2_X1 port map( A => n5146, B => n4621, Z => 
                           DP_OP_719J14_125_1055xn51);
   U5199 : NAND2_X1 port map( A1 => n5651, A2 => fromMemoryPortxLOADEDDATAx(16)
                           , ZN => n4622);
   U5200 : NAND2_X1 port map( A1 => n5653, A2 => n4622, ZN => add_x_26xBx16x);
   U5201 : INV_X1 port map( A => add_x_26xBx16x, ZN => n6783);
   U5202 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx16x,
                           B1 => n5012, B2 => fromRegsPortxREG_FILE_27xx16x, ZN
                           => n4626);
   U5203 : AOI22_X1 port map( A1 => n4980, A2 => fromRegsPortxREG_FILE_26xx16x,
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx16x, ZN
                           => n4625);
   U5204 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx16x,
                           B1 => n5013, B2 => fromRegsPortxREG_FILE_24xx16x, ZN
                           => n4624);
   U5205 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx16x,
                           B1 => n4946, B2 => fromRegsPortxREG_FILE_31xx16x, ZN
                           => n4623);
   U5206 : NAND4_X1 port map( A1 => n4626, A2 => n4625, A3 => n4624, A4 => 
                           n4623, ZN => n4632);
   U5207 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx16x,
                           B1 => n5019, B2 => fromRegsPortxREG_FILE_23xx16x, ZN
                           => n4630);
   U5208 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx16x,
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_19xx16x, ZN
                           => n4629);
   U5209 : AOI22_X1 port map( A1 => n4986, A2 => fromRegsPortxREG_FILE_18xx16x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx16x, ZN
                           => n4628);
   U5210 : NAND2_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx16x,
                           ZN => n4627);
   U5211 : NAND4_X1 port map( A1 => n4630, A2 => n4629, A3 => n4628, A4 => 
                           n4627, ZN => n4631);
   U5212 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4632
                           , A => n4631, ZN => n4638);
   U5213 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx16x,
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx16x, ZN
                           => n4637);
   U5214 : AOI22_X1 port map( A1 => n5305, A2 => fromRegsPortxREG_FILE_11xx16x,
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx16x, ZN
                           => n4634);
   U5215 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_12xx16x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx16x, ZN
                           => n4633);
   U5216 : NAND2_X1 port map( A1 => n4634, A2 => n4633, ZN => n4635);
   U5217 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx16x, B2 => n5060,
                           A => n4635, ZN => n4636);
   U5218 : OAI211_X1 port map( C1 => n4638, C2 => n7071, A => n4637, B => n4636
                           , ZN => n4639);
   U5219 : NAND2_X1 port map( A1 => n4639, A2 => n5133, ZN => n4649);
   U5220 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx16x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx16x, ZN
                           => n4643);
   U5221 : AOI22_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx16x,
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx16x, ZN
                           => n4642);
   U5222 : AOI22_X1 port map( A1 => n5035, A2 => fromRegsPortxREG_FILE_09xx16x,
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx16x, ZN
                           => n4641);
   U5223 : NAND2_X1 port map( A1 => n5036, A2 => fromRegsPortxREG_FILE_03xx16x,
                           ZN => n4640);
   U5224 : NAND4_X1 port map( A1 => n4643, A2 => n4642, A3 => n4641, A4 => 
                           n4640, ZN => n4647);
   U5225 : NAND2_X1 port map( A1 => n4760, A2 => fromRegsPortxREG_FILE_02xx16x,
                           ZN => n4645);
   U5226 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx16x, A2 => n5330,
                           ZN => n4644);
   U5227 : NAND2_X1 port map( A1 => n4645, A2 => n4644, ZN => n4646);
   U5228 : AOI21_X1 port map( B1 => n4647, B2 => n5334, A => n4646, ZN => n4648
                           );
   U5229 : NAND2_X1 port map( A1 => n4649, A2 => n4648, ZN => n6777);
   U5230 : INV_X1 port map( A => n6777, ZN => n7472);
   U5231 : OAI22_X1 port map( A1 => n5674, A2 => n6783, B1 => n7364, B2 => 
                           n7472, ZN => n4650);
   U5232 : XOR2_X1 port map( A => n7550, B => n4650, Z => 
                           DP_OP_719J14_125_1055xn52);
   U5233 : NAND2_X1 port map( A1 => n5651, A2 => fromMemoryPortxLOADEDDATAx(15)
                           , ZN => n4651);
   U5234 : NAND2_X1 port map( A1 => n5653, A2 => n4651, ZN => add_x_26xBx15x);
   U5235 : INV_X1 port map( A => add_x_26xBx15x, ZN => n6743);
   U5236 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx15x,
                           B1 => n5012, B2 => fromRegsPortxREG_FILE_27xx15x, ZN
                           => n4655);
   U5237 : AOI22_X1 port map( A1 => n4945, A2 => fromRegsPortxREG_FILE_29xx15x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_24xx15x, ZN
                           => n4654);
   U5238 : AOI22_X1 port map( A1 => n4980, A2 => fromRegsPortxREG_FILE_26xx15x,
                           B1 => n4978, B2 => fromRegsPortxREG_FILE_28xx15x, ZN
                           => n4653);
   U5239 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx15x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx15x, ZN
                           => n4652);
   U5240 : NAND4_X1 port map( A1 => n4655, A2 => n4654, A3 => n4653, A4 => 
                           n4652, ZN => n4661);
   U5241 : AOI22_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx15x,
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx15x, ZN
                           => n4659);
   U5242 : AOI22_X1 port map( A1 => n4985, A2 => fromRegsPortxREG_FILE_20xx15x,
                           B1 => n5019, B2 => fromRegsPortxREG_FILE_23xx15x, ZN
                           => n4658);
   U5243 : AOI22_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_19xx15x,
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx15x, ZN
                           => n4657);
   U5244 : NAND2_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx15x,
                           ZN => n4656);
   U5245 : NAND4_X1 port map( A1 => n4659, A2 => n4658, A3 => n4657, A4 => 
                           n4656, ZN => n4660);
   U5246 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4661
                           , A => n4660, ZN => n4667);
   U5247 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx15x,
                           B1 => n4957, B2 => fromRegsPortxREG_FILE_16xx15x, ZN
                           => n4666);
   U5248 : AOI22_X1 port map( A1 => n4995, A2 => fromRegsPortxREG_FILE_14xx15x,
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_11xx15x, ZN
                           => n4663);
   U5249 : AOI22_X1 port map( A1 => n5306, A2 => fromRegsPortxREG_FILE_13xx15x,
                           B1 => n4993, B2 => fromRegsPortxREG_FILE_15xx15x, ZN
                           => n4662);
   U5250 : NAND2_X1 port map( A1 => n4663, A2 => n4662, ZN => n4664);
   U5251 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx15x, B2 => n5303,
                           A => n4664, ZN => n4665);
   U5252 : OAI211_X1 port map( C1 => n4667, C2 => n5314, A => n4666, B => n4665
                           , ZN => n4668);
   U5253 : NAND2_X1 port map( A1 => n4668, A2 => n5133, ZN => n4678);
   U5254 : AOI22_X1 port map( A1 => n5035, A2 => fromRegsPortxREG_FILE_09xx15x,
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx15x, ZN
                           => n4672);
   U5255 : AOI22_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx15x,
                           B1 => n4932, B2 => fromRegsPortxREG_FILE_08xx15x, ZN
                           => n4671);
   U5256 : AOI22_X1 port map( A1 => n4965, A2 => fromRegsPortxREG_FILE_04xx15x,
                           B1 => n4903, B2 => fromRegsPortxREG_FILE_05xx15x, ZN
                           => n4670);
   U5257 : NAND2_X1 port map( A1 => n5036, A2 => fromRegsPortxREG_FILE_03xx15x,
                           ZN => n4669);
   U5258 : NAND4_X1 port map( A1 => n4672, A2 => n4671, A3 => n4670, A4 => 
                           n4669, ZN => n4676);
   U5259 : NAND2_X1 port map( A1 => n4760, A2 => fromRegsPortxREG_FILE_02xx15x,
                           ZN => n4674);
   U5260 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx15x, A2 => n5330,
                           ZN => n4673);
   U5261 : NAND2_X1 port map( A1 => n4674, A2 => n4673, ZN => n4675);
   U5262 : AOI21_X1 port map( B1 => n4676, B2 => n4973, A => n4675, ZN => n4677
                           );
   U5263 : NAND2_X1 port map( A1 => n4678, A2 => n4677, ZN => n6739);
   U5264 : INV_X1 port map( A => n6739, ZN => n7471);
   U5265 : OAI22_X1 port map( A1 => n5674, A2 => n6743, B1 => n7364, B2 => 
                           n7471, ZN => n4679);
   U5266 : XOR2_X1 port map( A => n5146, B => n4679, Z => 
                           DP_OP_719J14_125_1055xn53);
   U5267 : NAND2_X1 port map( A1 => n5651, A2 => fromMemoryPortxLOADEDDATAx(14)
                           , ZN => n4680);
   U5268 : NAND2_X1 port map( A1 => n5653, A2 => n4680, ZN => add_x_26xBx14x);
   U5269 : INV_X1 port map( A => add_x_26xBx14x, ZN => intadd_27xBx3x);
   U5270 : AOI22_X1 port map( A1 => n4979, A2 => fromRegsPortxREG_FILE_30xx14x,
                           B1 => n5278, B2 => fromRegsPortxREG_FILE_25xx14x, ZN
                           => n4684);
   U5271 : AOI22_X1 port map( A1 => n4980, A2 => fromRegsPortxREG_FILE_26xx14x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_24xx14x, ZN
                           => n4683);
   U5272 : AOI22_X1 port map( A1 => n4945, A2 => fromRegsPortxREG_FILE_29xx14x,
                           B1 => n4978, B2 => fromRegsPortxREG_FILE_28xx14x, ZN
                           => n4682);
   U5273 : AOI22_X1 port map( A1 => n5281, A2 => fromRegsPortxREG_FILE_27xx14x,
                           B1 => n4946, B2 => fromRegsPortxREG_FILE_31xx14x, ZN
                           => n4681);
   U5274 : NAND4_X1 port map( A1 => n4684, A2 => n4683, A3 => n4682, A4 => 
                           n4681, ZN => n4690);
   U5275 : AOI22_X1 port map( A1 => n4986, A2 => fromRegsPortxREG_FILE_18xx14x,
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_19xx14x, ZN
                           => n4688);
   U5276 : AOI22_X1 port map( A1 => n5052, A2 => fromRegsPortxREG_FILE_21xx14x,
                           B1 => n5018, B2 => fromRegsPortxREG_FILE_17xx14x, ZN
                           => n4687);
   U5277 : AOI22_X1 port map( A1 => n5019, A2 => fromRegsPortxREG_FILE_23xx14x,
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_22xx14x, ZN
                           => n4686);
   U5278 : NAND2_X1 port map( A1 => n4985, A2 => fromRegsPortxREG_FILE_20xx14x,
                           ZN => n4685);
   U5279 : NAND4_X1 port map( A1 => n4688, A2 => n4687, A3 => n4686, A4 => 
                           n4685, ZN => n4689);
   U5280 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4690
                           , A => n4689, ZN => n4696);
   U5281 : AOI22_X1 port map( A1 => n4995, A2 => fromRegsPortxREG_FILE_14xx14x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx14x, ZN
                           => n4695);
   U5282 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx14x,
                           B1 => n4993, B2 => fromRegsPortxREG_FILE_15xx14x, ZN
                           => n4692);
   U5283 : AOI22_X1 port map( A1 => n4994, A2 => fromRegsPortxREG_FILE_11xx14x,
                           B1 => n4957, B2 => fromRegsPortxREG_FILE_16xx14x, ZN
                           => n4691);
   U5284 : NAND2_X1 port map( A1 => n4692, A2 => n4691, ZN => n4693);
   U5285 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx14x, B2 => n5303,
                           A => n4693, ZN => n4694);
   U5286 : OAI211_X1 port map( C1 => n4696, C2 => n5314, A => n4695, B => n4694
                           , ZN => n4697);
   U5287 : NAND2_X1 port map( A1 => n4697, A2 => n5133, ZN => n4707);
   U5288 : AOI22_X1 port map( A1 => n4903, A2 => fromRegsPortxREG_FILE_05xx14x,
                           B1 => n5033, B2 => fromRegsPortxREG_FILE_07xx14x, ZN
                           => n4701);
   U5289 : AOI22_X1 port map( A1 => n4965, A2 => fromRegsPortxREG_FILE_04xx14x,
                           B1 => n5034, B2 => fromRegsPortxREG_FILE_06xx14x, ZN
                           => n4700);
   U5290 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx14x,
                           B1 => n4932, B2 => fromRegsPortxREG_FILE_08xx14x, ZN
                           => n4699);
   U5291 : NAND2_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx14x,
                           ZN => n4698);
   U5292 : NAND4_X1 port map( A1 => n4701, A2 => n4700, A3 => n4699, A4 => 
                           n4698, ZN => n4705);
   U5293 : NAND2_X1 port map( A1 => n4760, A2 => fromRegsPortxREG_FILE_02xx14x,
                           ZN => n4703);
   U5294 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx14x, A2 => n5330,
                           ZN => n4702);
   U5295 : NAND2_X1 port map( A1 => n4703, A2 => n4702, ZN => n4704);
   U5296 : AOI21_X1 port map( B1 => n4705, B2 => n4973, A => n4704, ZN => n4706
                           );
   U5297 : NAND2_X1 port map( A1 => n4707, A2 => n4706, ZN => n6693);
   U5298 : INV_X1 port map( A => n6693, ZN => n7470);
   U5299 : OAI22_X1 port map( A1 => n5674, A2 => intadd_27xBx3x, B1 => n7364, 
                           B2 => n7470, ZN => n4708);
   U5300 : XOR2_X1 port map( A => n5146, B => n4708, Z => 
                           DP_OP_719J14_125_1055xn54);
   U5301 : NAND2_X1 port map( A1 => n5651, A2 => fromMemoryPortxLOADEDDATAx(13)
                           , ZN => n4709);
   U5302 : NAND2_X1 port map( A1 => n5653, A2 => n4709, ZN => add_x_26xBx13x);
   U5303 : INV_X1 port map( A => add_x_26xBx13x, ZN => intadd_27xBx2x);
   U5304 : AOI22_X1 port map( A1 => n5278, A2 => fromRegsPortxREG_FILE_25xx13x,
                           B1 => n5012, B2 => fromRegsPortxREG_FILE_27xx13x, ZN
                           => n4713);
   U5305 : AOI22_X1 port map( A1 => n4979, A2 => fromRegsPortxREG_FILE_30xx13x,
                           B1 => n4980, B2 => fromRegsPortxREG_FILE_26xx13x, ZN
                           => n4712);
   U5306 : AOI22_X1 port map( A1 => n4945, A2 => fromRegsPortxREG_FILE_29xx13x,
                           B1 => n4978, B2 => fromRegsPortxREG_FILE_28xx13x, ZN
                           => n4711);
   U5307 : AOI22_X1 port map( A1 => n5282, A2 => fromRegsPortxREG_FILE_24xx13x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx13x, ZN
                           => n4710);
   U5308 : NAND4_X1 port map( A1 => n4713, A2 => n4712, A3 => n4711, A4 => 
                           n4710, ZN => n4719);
   U5309 : AOI22_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx13x,
                           B1 => n5018, B2 => fromRegsPortxREG_FILE_17xx13x, ZN
                           => n4717);
   U5310 : AOI22_X1 port map( A1 => n4985, A2 => fromRegsPortxREG_FILE_20xx13x,
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx13x, ZN
                           => n4716);
   U5311 : AOI22_X1 port map( A1 => n5052, A2 => fromRegsPortxREG_FILE_21xx13x,
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_19xx13x, ZN
                           => n4715);
   U5312 : NAND2_X1 port map( A1 => n5019, A2 => fromRegsPortxREG_FILE_23xx13x,
                           ZN => n4714);
   U5313 : NAND4_X1 port map( A1 => n4717, A2 => n4716, A3 => n4715, A4 => 
                           n4714, ZN => n4718);
   U5314 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4719
                           , A => n4718, ZN => n4725);
   U5315 : AOI22_X1 port map( A1 => n4957, A2 => fromRegsPortxREG_FILE_16xx13x,
                           B1 => n4993, B2 => fromRegsPortxREG_FILE_15xx13x, ZN
                           => n4724);
   U5316 : AOI22_X1 port map( A1 => n4995, A2 => fromRegsPortxREG_FILE_14xx13x,
                           B1 => n4994, B2 => fromRegsPortxREG_FILE_11xx13x, ZN
                           => n4721);
   U5317 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_12xx13x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx13x, ZN
                           => n4720);
   U5318 : NAND2_X1 port map( A1 => n4721, A2 => n4720, ZN => n4722);
   U5319 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx13x, B2 => n5302,
                           A => n4722, ZN => n4723);
   U5320 : OAI211_X1 port map( C1 => n4725, C2 => n5314, A => n4724, B => n4723
                           , ZN => n4726);
   U5321 : NAND2_X1 port map( A1 => n4726, A2 => n5133, ZN => n4736);
   U5322 : AOI22_X1 port map( A1 => n4965, A2 => fromRegsPortxREG_FILE_04xx13x,
                           B1 => n5033, B2 => fromRegsPortxREG_FILE_07xx13x, ZN
                           => n4730);
   U5323 : AOI22_X1 port map( A1 => n5035, A2 => fromRegsPortxREG_FILE_09xx13x,
                           B1 => n4932, B2 => fromRegsPortxREG_FILE_08xx13x, ZN
                           => n4729);
   U5324 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx13x,
                           B1 => n4903, B2 => fromRegsPortxREG_FILE_05xx13x, ZN
                           => n4728);
   U5325 : NAND2_X1 port map( A1 => n5034, A2 => fromRegsPortxREG_FILE_06xx13x,
                           ZN => n4727);
   U5326 : NAND4_X1 port map( A1 => n4730, A2 => n4729, A3 => n4728, A4 => 
                           n4727, ZN => n4734);
   U5327 : NAND2_X1 port map( A1 => n4760, A2 => fromRegsPortxREG_FILE_02xx13x,
                           ZN => n4732);
   U5328 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx13x, A2 => n5330,
                           ZN => n4731);
   U5329 : NAND2_X1 port map( A1 => n4732, A2 => n4731, ZN => n4733);
   U5330 : AOI21_X1 port map( B1 => n4734, B2 => n4973, A => n4733, ZN => n4735
                           );
   U5331 : NAND2_X1 port map( A1 => n4736, A2 => n4735, ZN => n6669);
   U5332 : INV_X1 port map( A => n6669, ZN => n7469);
   U5333 : OAI22_X1 port map( A1 => n5674, A2 => intadd_27xBx2x, B1 => n7364, 
                           B2 => n7469, ZN => n4737);
   U5334 : XOR2_X1 port map( A => n7550, B => n4737, Z => 
                           DP_OP_719J14_125_1055xn55);
   U5335 : NAND2_X1 port map( A1 => n5651, A2 => fromMemoryPortxLOADEDDATAx(12)
                           , ZN => n4738);
   U5336 : NAND2_X1 port map( A1 => n5653, A2 => n4738, ZN => add_x_26xBx12x);
   U5337 : INV_X1 port map( A => add_x_26xBx12x, ZN => intadd_27xBx1x);
   U5338 : AOI22_X1 port map( A1 => n4979, A2 => fromRegsPortxREG_FILE_30xx12x,
                           B1 => n4980, B2 => fromRegsPortxREG_FILE_26xx12x, ZN
                           => n4742);
   U5339 : AOI22_X1 port map( A1 => n5281, A2 => fromRegsPortxREG_FILE_27xx12x,
                           B1 => n4978, B2 => fromRegsPortxREG_FILE_28xx12x, ZN
                           => n4741);
   U5340 : AOI22_X1 port map( A1 => n5080, A2 => fromRegsPortxREG_FILE_25xx12x,
                           B1 => n4945, B2 => fromRegsPortxREG_FILE_29xx12x, ZN
                           => n4740);
   U5341 : AOI22_X1 port map( A1 => n5013, A2 => fromRegsPortxREG_FILE_24xx12x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx12x, ZN
                           => n4739);
   U5342 : NAND4_X1 port map( A1 => n4742, A2 => n4741, A3 => n4740, A4 => 
                           n4739, ZN => n4748);
   U5343 : AOI22_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_19xx12x,
                           B1 => n5018, B2 => fromRegsPortxREG_FILE_17xx12x, ZN
                           => n4746);
   U5344 : AOI22_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx12x,
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx12x, ZN
                           => n4745);
   U5345 : AOI22_X1 port map( A1 => n4985, A2 => fromRegsPortxREG_FILE_20xx12x,
                           B1 => n5019, B2 => fromRegsPortxREG_FILE_23xx12x, ZN
                           => n4744);
   U5346 : NAND2_X1 port map( A1 => n5052, A2 => fromRegsPortxREG_FILE_21xx12x,
                           ZN => n4743);
   U5347 : NAND4_X1 port map( A1 => n4746, A2 => n4745, A3 => n4744, A4 => 
                           n4743, ZN => n4747);
   U5348 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4748
                           , A => n4747, ZN => n4754);
   U5349 : AOI22_X1 port map( A1 => n4994, A2 => fromRegsPortxREG_FILE_11xx12x,
                           B1 => n4957, B2 => fromRegsPortxREG_FILE_16xx12x, ZN
                           => n4753);
   U5350 : AOI22_X1 port map( A1 => n5060, A2 => fromRegsPortxREG_FILE_10xx12x,
                           B1 => n4993, B2 => fromRegsPortxREG_FILE_15xx12x, ZN
                           => n4750);
   U5351 : AOI22_X1 port map( A1 => n4995, A2 => fromRegsPortxREG_FILE_14xx12x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx12x, ZN
                           => n4749);
   U5352 : NAND2_X1 port map( A1 => n4750, A2 => n4749, ZN => n4751);
   U5353 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx12x, B2 => n5129,
                           A => n4751, ZN => n4752);
   U5354 : OAI211_X1 port map( C1 => n4754, C2 => n5314, A => n4753, B => n4752
                           , ZN => n4755);
   U5355 : NAND2_X1 port map( A1 => n4755, A2 => n5133, ZN => n4766);
   U5356 : AOI22_X1 port map( A1 => n5035, A2 => fromRegsPortxREG_FILE_09xx12x,
                           B1 => n5033, B2 => fromRegsPortxREG_FILE_07xx12x, ZN
                           => n4759);
   U5357 : AOI22_X1 port map( A1 => n4965, A2 => fromRegsPortxREG_FILE_04xx12x,
                           B1 => n5034, B2 => fromRegsPortxREG_FILE_06xx12x, ZN
                           => n4758);
   U5358 : AOI22_X1 port map( A1 => n4932, A2 => fromRegsPortxREG_FILE_08xx12x,
                           B1 => n4903, B2 => fromRegsPortxREG_FILE_05xx12x, ZN
                           => n4757);
   U5359 : NAND2_X1 port map( A1 => n5036, A2 => fromRegsPortxREG_FILE_03xx12x,
                           ZN => n4756);
   U5360 : NAND4_X1 port map( A1 => n4759, A2 => n4758, A3 => n4757, A4 => 
                           n4756, ZN => n4764);
   U5361 : NAND2_X1 port map( A1 => n4760, A2 => fromRegsPortxREG_FILE_02xx12x,
                           ZN => n4762);
   U5362 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx12x, A2 => n5072,
                           ZN => n4761);
   U5363 : NAND2_X1 port map( A1 => n4762, A2 => n4761, ZN => n4763);
   U5364 : AOI21_X1 port map( B1 => n4764, B2 => n4973, A => n4763, ZN => n4765
                           );
   U5365 : NAND2_X1 port map( A1 => n4766, A2 => n4765, ZN => n6626);
   U5366 : INV_X1 port map( A => n6626, ZN => n7468);
   U5367 : OAI22_X1 port map( A1 => n7468, A2 => n5676, B1 => n5675, B2 => 
                           intadd_27xBx1x, ZN => n4767);
   U5368 : XOR2_X1 port map( A => n5146, B => n4767, Z => 
                           DP_OP_719J14_125_1055xn56);
   U5369 : NAND2_X1 port map( A1 => n4768, A2 => fromMemoryPortxLOADEDDATAx(7),
                           ZN => n4773);
   U5370 : INV_X1 port map( A => n4769, ZN => n4770);
   U5371 : OAI21_X1 port map( B1 => n5642, B2 => n6954, A => n4770, ZN => n4771
                           );
   U5372 : INV_X1 port map( A => n4771, ZN => n4772);
   U5373 : NAND2_X1 port map( A1 => n4773, A2 => n4772, ZN => add_x_26xBx11x);
   U5374 : INV_X1 port map( A => add_x_26xBx11x, ZN => intadd_27xBx0x);
   U5375 : AOI22_X1 port map( A1 => n5080, A2 => fromRegsPortxREG_FILE_25xx11x,
                           B1 => n4978, B2 => fromRegsPortxREG_FILE_28xx11x, ZN
                           => n4777);
   U5376 : AOI22_X1 port map( A1 => n4979, A2 => fromRegsPortxREG_FILE_30xx11x,
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx11x, ZN
                           => n4776);
   U5377 : AOI22_X1 port map( A1 => n4945, A2 => fromRegsPortxREG_FILE_29xx11x,
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_24xx11x, ZN
                           => n4775);
   U5378 : AOI22_X1 port map( A1 => n5281, A2 => fromRegsPortxREG_FILE_27xx11x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx11x, ZN
                           => n4774);
   U5379 : NAND4_X1 port map( A1 => n4777, A2 => n4776, A3 => n4775, A4 => 
                           n4774, ZN => n4783);
   U5380 : AOI22_X1 port map( A1 => n4986, A2 => fromRegsPortxREG_FILE_18xx11x,
                           B1 => n5018, B2 => fromRegsPortxREG_FILE_17xx11x, ZN
                           => n4781);
   U5381 : AOI22_X1 port map( A1 => n5052, A2 => fromRegsPortxREG_FILE_21xx11x,
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_19xx11x, ZN
                           => n4780);
   U5382 : AOI22_X1 port map( A1 => n5019, A2 => fromRegsPortxREG_FILE_23xx11x,
                           B1 => n5289, B2 => fromRegsPortxREG_FILE_22xx11x, ZN
                           => n4779);
   U5383 : NAND2_X1 port map( A1 => n4985, A2 => fromRegsPortxREG_FILE_20xx11x,
                           ZN => n4778);
   U5384 : NAND4_X1 port map( A1 => n4781, A2 => n4780, A3 => n4779, A4 => 
                           n4778, ZN => n4782);
   U5385 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4783
                           , A => n4782, ZN => n4789);
   U5386 : AOI22_X1 port map( A1 => n4957, A2 => fromRegsPortxREG_FILE_16xx11x,
                           B1 => n4993, B2 => fromRegsPortxREG_FILE_15xx11x, ZN
                           => n4788);
   U5387 : AOI22_X1 port map( A1 => n5060, A2 => fromRegsPortxREG_FILE_10xx11x,
                           B1 => n4994, B2 => fromRegsPortxREG_FILE_11xx11x, ZN
                           => n4785);
   U5388 : AOI22_X1 port map( A1 => n4995, A2 => fromRegsPortxREG_FILE_14xx11x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx11x, ZN
                           => n4784);
   U5389 : NAND2_X1 port map( A1 => n4785, A2 => n4784, ZN => n4786);
   U5390 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx11x, B2 => n5129,
                           A => n4786, ZN => n4787);
   U5391 : OAI211_X1 port map( C1 => n4789, C2 => n5314, A => n4788, B => n4787
                           , ZN => n4790);
   U5392 : NAND2_X1 port map( A1 => n4790, A2 => n5316, ZN => n4800);
   U5393 : AOI22_X1 port map( A1 => n4965, A2 => fromRegsPortxREG_FILE_04xx11x,
                           B1 => n5036, B2 => fromRegsPortxREG_FILE_03xx11x, ZN
                           => n4794);
   U5394 : AOI22_X1 port map( A1 => n5035, A2 => fromRegsPortxREG_FILE_09xx11x,
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx11x, ZN
                           => n4793);
   U5395 : AOI22_X1 port map( A1 => n4932, A2 => fromRegsPortxREG_FILE_08xx11x,
                           B1 => n5033, B2 => fromRegsPortxREG_FILE_07xx11x, ZN
                           => n4792);
   U5396 : NAND2_X1 port map( A1 => n5034, A2 => fromRegsPortxREG_FILE_06xx11x,
                           ZN => n4791);
   U5397 : NAND4_X1 port map( A1 => n4794, A2 => n4793, A3 => n4792, A4 => 
                           n4791, ZN => n4798);
   U5398 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx11x,
                           ZN => n4796);
   U5399 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx11x, A2 => n5072,
                           ZN => n4795);
   U5400 : NAND2_X1 port map( A1 => n4796, A2 => n4795, ZN => n4797);
   U5401 : AOI21_X1 port map( B1 => n4798, B2 => n4973, A => n4797, ZN => n4799
                           );
   U5402 : NAND2_X1 port map( A1 => n4800, A2 => n4799, ZN => n6553);
   U5403 : INV_X1 port map( A => n6553, ZN => n7467);
   U5404 : OAI22_X1 port map( A1 => n5674, A2 => intadd_27xBx0x, B1 => n7364, 
                           B2 => n7467, ZN => n4801);
   U5405 : XOR2_X1 port map( A => n5146, B => n4801, Z => 
                           DP_OP_719J14_125_1055xn57);
   U5406 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(30), A2 => n4944,
                           ZN => add_x_26xBx10x);
   U5407 : INV_X1 port map( A => add_x_26xBx10x, ZN => n5814);
   U5408 : AOI22_X1 port map( A1 => n5080, A2 => fromRegsPortxREG_FILE_25xx10x,
                           B1 => n4980, B2 => fromRegsPortxREG_FILE_26xx10x, ZN
                           => n4805);
   U5409 : AOI22_X1 port map( A1 => n4979, A2 => fromRegsPortxREG_FILE_30xx10x,
                           B1 => n5012, B2 => fromRegsPortxREG_FILE_27xx10x, ZN
                           => n4804);
   U5410 : AOI22_X1 port map( A1 => n5013, A2 => fromRegsPortxREG_FILE_24xx10x,
                           B1 => n4978, B2 => fromRegsPortxREG_FILE_28xx10x, ZN
                           => n4803);
   U5411 : AOI22_X1 port map( A1 => n4945, A2 => fromRegsPortxREG_FILE_29xx10x,
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx10x, ZN
                           => n4802);
   U5412 : NAND4_X1 port map( A1 => n4805, A2 => n4804, A3 => n4803, A4 => 
                           n4802, ZN => n4811);
   U5413 : AOI22_X1 port map( A1 => n4985, A2 => fromRegsPortxREG_FILE_20xx10x,
                           B1 => n5289, B2 => fromRegsPortxREG_FILE_22xx10x, ZN
                           => n4809);
   U5414 : AOI22_X1 port map( A1 => n5019, A2 => fromRegsPortxREG_FILE_23xx10x,
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_19xx10x, ZN
                           => n4808);
   U5415 : AOI22_X1 port map( A1 => n5052, A2 => fromRegsPortxREG_FILE_21xx10x,
                           B1 => n5018, B2 => fromRegsPortxREG_FILE_17xx10x, ZN
                           => n4807);
   U5416 : NAND2_X1 port map( A1 => n5295, A2 => fromRegsPortxREG_FILE_18xx10x,
                           ZN => n4806);
   U5417 : NAND4_X1 port map( A1 => n4809, A2 => n4808, A3 => n4807, A4 => 
                           n4806, ZN => n4810);
   U5418 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4811
                           , A => n4810, ZN => n4817);
   U5419 : AOI22_X1 port map( A1 => n4994, A2 => fromRegsPortxREG_FILE_11xx10x,
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx10x, ZN
                           => n4816);
   U5420 : AOI22_X1 port map( A1 => n5060, A2 => fromRegsPortxREG_FILE_10xx10x,
                           B1 => n4993, B2 => fromRegsPortxREG_FILE_15xx10x, ZN
                           => n4813);
   U5421 : AOI22_X1 port map( A1 => n4995, A2 => fromRegsPortxREG_FILE_14xx10x,
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx10x, ZN
                           => n4812);
   U5422 : NAND2_X1 port map( A1 => n4813, A2 => n4812, ZN => n4814);
   U5423 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx10x, B2 => n5129,
                           A => n4814, ZN => n4815);
   U5424 : OAI211_X1 port map( C1 => n4817, C2 => n5314, A => n4816, B => n4815
                           , ZN => n4818);
   U5425 : NAND2_X1 port map( A1 => n4818, A2 => n5316, ZN => n4828);
   U5426 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx10x,
                           B1 => n4903, B2 => fromRegsPortxREG_FILE_05xx10x, ZN
                           => n4822);
   U5427 : AOI22_X1 port map( A1 => n5034, A2 => fromRegsPortxREG_FILE_06xx10x,
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx10x, ZN
                           => n4821);
   U5428 : AOI22_X1 port map( A1 => n4965, A2 => fromRegsPortxREG_FILE_04xx10x,
                           B1 => n5033, B2 => fromRegsPortxREG_FILE_07xx10x, ZN
                           => n4820);
   U5429 : NAND2_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx10x,
                           ZN => n4819);
   U5430 : NAND4_X1 port map( A1 => n4822, A2 => n4821, A3 => n4820, A4 => 
                           n4819, ZN => n4826);
   U5431 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx10x,
                           ZN => n4824);
   U5432 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx10x, A2 => n5072,
                           ZN => n4823);
   U5433 : NAND2_X1 port map( A1 => n4824, A2 => n4823, ZN => n4825);
   U5434 : AOI21_X1 port map( B1 => n4826, B2 => n4973, A => n4825, ZN => n4827
                           );
   U5435 : NAND2_X1 port map( A1 => n4828, A2 => n4827, ZN => n6530);
   U5436 : INV_X1 port map( A => n6530, ZN => n7466);
   U5437 : OAI22_X1 port map( A1 => n5674, A2 => n5814, B1 => n7364, B2 => 
                           n7466, ZN => n4829);
   U5438 : XOR2_X1 port map( A => n7550, B => n4829, Z => 
                           DP_OP_719J14_125_1055xn58);
   U5439 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(29), A2 => n4944,
                           ZN => add_x_26xBx9x);
   U5440 : AOI22_X1 port map( A1 => n4945, A2 => fromRegsPortxREG_FILE_29xx9x, 
                           B1 => n5012, B2 => fromRegsPortxREG_FILE_27xx9x, ZN 
                           => n4833);
   U5441 : AOI22_X1 port map( A1 => n5080, A2 => fromRegsPortxREG_FILE_25xx9x, 
                           B1 => n4978, B2 => fromRegsPortxREG_FILE_28xx9x, ZN 
                           => n4832);
   U5442 : AOI22_X1 port map( A1 => n4979, A2 => fromRegsPortxREG_FILE_30xx9x, 
                           B1 => n4980, B2 => fromRegsPortxREG_FILE_26xx9x, ZN 
                           => n4831);
   U5443 : AOI22_X1 port map( A1 => n5282, A2 => fromRegsPortxREG_FILE_24xx9x, 
                           B1 => n4946, B2 => fromRegsPortxREG_FILE_31xx9x, ZN 
                           => n4830);
   U5444 : NAND4_X1 port map( A1 => n4833, A2 => n4832, A3 => n4831, A4 => 
                           n4830, ZN => n4839);
   U5445 : AOI22_X1 port map( A1 => n5052, A2 => fromRegsPortxREG_FILE_21xx9x, 
                           B1 => n5018, B2 => fromRegsPortxREG_FILE_17xx9x, ZN 
                           => n4837);
   U5446 : AOI22_X1 port map( A1 => n4986, A2 => fromRegsPortxREG_FILE_18xx9x, 
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_19xx9x, ZN 
                           => n4836);
   U5447 : AOI22_X1 port map( A1 => n5019, A2 => fromRegsPortxREG_FILE_23xx9x, 
                           B1 => n5289, B2 => fromRegsPortxREG_FILE_22xx9x, ZN 
                           => n4835);
   U5448 : NAND2_X1 port map( A1 => n4985, A2 => fromRegsPortxREG_FILE_20xx9x, 
                           ZN => n4834);
   U5449 : NAND4_X1 port map( A1 => n4837, A2 => n4836, A3 => n4835, A4 => 
                           n4834, ZN => n4838);
   U5450 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4839
                           , A => n4838, ZN => n4845);
   U5451 : AOI22_X1 port map( A1 => n4995, A2 => fromRegsPortxREG_FILE_14xx9x, 
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx9x, ZN 
                           => n4844);
   U5452 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx9x, 
                           B1 => n4993, B2 => fromRegsPortxREG_FILE_15xx9x, ZN 
                           => n4841);
   U5453 : AOI22_X1 port map( A1 => n4994, A2 => fromRegsPortxREG_FILE_11xx9x, 
                           B1 => n4957, B2 => fromRegsPortxREG_FILE_16xx9x, ZN 
                           => n4840);
   U5454 : NAND2_X1 port map( A1 => n4841, A2 => n4840, ZN => n4842);
   U5455 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx9x, B2 => n5303, 
                           A => n4842, ZN => n4843);
   U5456 : OAI211_X1 port map( C1 => n4845, C2 => n5314, A => n4844, B => n4843
                           , ZN => n4846);
   U5457 : NAND2_X1 port map( A1 => n4846, A2 => n5316, ZN => n4856);
   U5458 : AOI22_X1 port map( A1 => n4932, A2 => fromRegsPortxREG_FILE_08xx9x, 
                           B1 => n5033, B2 => fromRegsPortxREG_FILE_07xx9x, ZN 
                           => n4850);
   U5459 : AOI22_X1 port map( A1 => n4965, A2 => fromRegsPortxREG_FILE_04xx9x, 
                           B1 => n4903, B2 => fromRegsPortxREG_FILE_05xx9x, ZN 
                           => n4849);
   U5460 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx9x, 
                           B1 => n5034, B2 => fromRegsPortxREG_FILE_06xx9x, ZN 
                           => n4848);
   U5461 : NAND2_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx9x, 
                           ZN => n4847);
   U5462 : NAND4_X1 port map( A1 => n4850, A2 => n4849, A3 => n4848, A4 => 
                           n4847, ZN => n4854);
   U5463 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx9x, 
                           ZN => n4852);
   U5464 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx9x, A2 => n5072, 
                           ZN => n4851);
   U5465 : NAND2_X1 port map( A1 => n4852, A2 => n4851, ZN => n4853);
   U5466 : AOI21_X1 port map( B1 => n4854, B2 => n4973, A => n4853, ZN => n4855
                           );
   U5467 : NAND2_X1 port map( A1 => n4856, A2 => n4855, ZN => n6480);
   U5468 : INV_X1 port map( A => n6480, ZN => n7465);
   U5469 : INV_X1 port map( A => add_x_26xBx9x, ZN => n6476);
   U5470 : OAI22_X1 port map( A1 => n7465, A2 => n5677, B1 => n5675, B2 => 
                           n6476, ZN => n4857);
   U5471 : XOR2_X1 port map( A => n5146, B => n4857, Z => 
                           DP_OP_719J14_125_1055xn59);
   U5472 : INV_X1 port map( A => add_x_26xBx8x, ZN => n5587);
   U5473 : AOI22_X1 port map( A1 => n5013, A2 => fromRegsPortxREG_FILE_24xx8x, 
                           B1 => n4978, B2 => fromRegsPortxREG_FILE_28xx8x, ZN 
                           => n4861);
   U5474 : AOI22_X1 port map( A1 => n4979, A2 => fromRegsPortxREG_FILE_30xx8x, 
                           B1 => n4980, B2 => fromRegsPortxREG_FILE_26xx8x, ZN 
                           => n4860);
   U5475 : AOI22_X1 port map( A1 => n4945, A2 => fromRegsPortxREG_FILE_29xx8x, 
                           B1 => n5012, B2 => fromRegsPortxREG_FILE_27xx8x, ZN 
                           => n4859);
   U5476 : AOI22_X1 port map( A1 => n5080, A2 => fromRegsPortxREG_FILE_25xx8x, 
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx8x, ZN 
                           => n4858);
   U5477 : NAND4_X1 port map( A1 => n4861, A2 => n4860, A3 => n4859, A4 => 
                           n4858, ZN => n4867);
   U5478 : AOI22_X1 port map( A1 => n4985, A2 => fromRegsPortxREG_FILE_20xx8x, 
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx8x, ZN 
                           => n4865);
   U5479 : AOI22_X1 port map( A1 => n5019, A2 => fromRegsPortxREG_FILE_23xx8x, 
                           B1 => n5018, B2 => fromRegsPortxREG_FILE_17xx8x, ZN 
                           => n4864);
   U5480 : AOI22_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx8x, 
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_19xx8x, ZN 
                           => n4863);
   U5481 : NAND2_X1 port map( A1 => n5052, A2 => fromRegsPortxREG_FILE_21xx8x, 
                           ZN => n4862);
   U5482 : NAND4_X1 port map( A1 => n4865, A2 => n4864, A3 => n4863, A4 => 
                           n4862, ZN => n4866);
   U5483 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4867
                           , A => n4866, ZN => n4873);
   U5484 : AOI22_X1 port map( A1 => n4995, A2 => fromRegsPortxREG_FILE_14xx8x, 
                           B1 => n4957, B2 => fromRegsPortxREG_FILE_16xx8x, ZN 
                           => n4872);
   U5485 : AOI22_X1 port map( A1 => n4994, A2 => fromRegsPortxREG_FILE_11xx8x, 
                           B1 => n4993, B2 => fromRegsPortxREG_FILE_15xx8x, ZN 
                           => n4869);
   U5486 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_12xx8x, 
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx8x, ZN 
                           => n4868);
   U5487 : NAND2_X1 port map( A1 => n4869, A2 => n4868, ZN => n4870);
   U5488 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx8x, B2 => n5302, 
                           A => n4870, ZN => n4871);
   U5489 : OAI211_X1 port map( C1 => n4873, C2 => n5314, A => n4872, B => n4871
                           , ZN => n4874);
   U5490 : NAND2_X1 port map( A1 => n4874, A2 => n5316, ZN => n4884);
   U5491 : AOI22_X1 port map( A1 => n5035, A2 => fromRegsPortxREG_FILE_09xx8x, 
                           B1 => n5036, B2 => fromRegsPortxREG_FILE_03xx8x, ZN 
                           => n4878);
   U5492 : AOI22_X1 port map( A1 => n4965, A2 => fromRegsPortxREG_FILE_04xx8x, 
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx8x, ZN 
                           => n4877);
   U5493 : AOI22_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx8x, 
                           B1 => n5033, B2 => fromRegsPortxREG_FILE_07xx8x, ZN 
                           => n4876);
   U5494 : NAND2_X1 port map( A1 => n4903, A2 => fromRegsPortxREG_FILE_05xx8x, 
                           ZN => n4875);
   U5495 : NAND4_X1 port map( A1 => n4878, A2 => n4877, A3 => n4876, A4 => 
                           n4875, ZN => n4882);
   U5496 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx8x, 
                           ZN => n4880);
   U5497 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx8x, A2 => n5072, 
                           ZN => n4879);
   U5498 : NAND2_X1 port map( A1 => n4880, A2 => n4879, ZN => n4881);
   U5499 : AOI21_X1 port map( B1 => n4882, B2 => n4973, A => n4881, ZN => n4883
                           );
   U5500 : NAND2_X1 port map( A1 => n4884, A2 => n4883, ZN => n6421);
   U5501 : INV_X1 port map( A => n6421, ZN => n7464);
   U5502 : OAI22_X1 port map( A1 => n5674, A2 => n5587, B1 => n7364, B2 => 
                           n7464, ZN => n4885);
   U5503 : XOR2_X1 port map( A => n5146, B => n4885, Z => 
                           DP_OP_719J14_125_1055xn60);
   U5504 : INV_X1 port map( A => add_x_26xBx7x, ZN => n6394);
   U5505 : AOI22_X1 port map( A1 => n5080, A2 => fromRegsPortxREG_FILE_25xx7x, 
                           B1 => n4978, B2 => fromRegsPortxREG_FILE_28xx7x, ZN 
                           => n4889);
   U5506 : AOI22_X1 port map( A1 => n4980, A2 => fromRegsPortxREG_FILE_26xx7x, 
                           B1 => n5012, B2 => fromRegsPortxREG_FILE_27xx7x, ZN 
                           => n4888);
   U5507 : AOI22_X1 port map( A1 => n4979, A2 => fromRegsPortxREG_FILE_30xx7x, 
                           B1 => n4945, B2 => fromRegsPortxREG_FILE_29xx7x, ZN 
                           => n4887);
   U5508 : AOI22_X1 port map( A1 => n5013, A2 => fromRegsPortxREG_FILE_24xx7x, 
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx7x, ZN 
                           => n4886);
   U5509 : NAND4_X1 port map( A1 => n4889, A2 => n4888, A3 => n4887, A4 => 
                           n4886, ZN => n4895);
   U5510 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx7x, 
                           B1 => n5290, B2 => fromRegsPortxREG_FILE_21xx7x, ZN 
                           => n4893);
   U5511 : AOI22_X1 port map( A1 => n4986, A2 => fromRegsPortxREG_FILE_18xx7x, 
                           B1 => n5018, B2 => fromRegsPortxREG_FILE_17xx7x, ZN 
                           => n4892);
   U5512 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx7x, 
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_19xx7x, ZN 
                           => n4891);
   U5513 : NAND2_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_22xx7x, 
                           ZN => n4890);
   U5514 : NAND4_X1 port map( A1 => n4893, A2 => n4892, A3 => n4891, A4 => 
                           n4890, ZN => n4894);
   U5515 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4895
                           , A => n4894, ZN => n4901);
   U5516 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_12xx7x, 
                           B1 => n4993, B2 => fromRegsPortxREG_FILE_15xx7x, ZN 
                           => n4900);
   U5517 : AOI22_X1 port map( A1 => n5060, A2 => fromRegsPortxREG_FILE_10xx7x, 
                           B1 => n4994, B2 => fromRegsPortxREG_FILE_11xx7x, ZN 
                           => n4897);
   U5518 : AOI22_X1 port map( A1 => n4957, A2 => fromRegsPortxREG_FILE_16xx7x, 
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx7x, ZN 
                           => n4896);
   U5519 : NAND2_X1 port map( A1 => n4897, A2 => n4896, ZN => n4898);
   U5520 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_14xx7x, B2 => n4995, 
                           A => n4898, ZN => n4899);
   U5521 : OAI211_X1 port map( C1 => n4901, C2 => n5314, A => n4900, B => n4899
                           , ZN => n4902);
   U5522 : NAND2_X1 port map( A1 => n4902, A2 => n5316, ZN => n4913);
   U5523 : AOI22_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx7x, 
                           B1 => n5033, B2 => fromRegsPortxREG_FILE_07xx7x, ZN 
                           => n4907);
   U5524 : AOI22_X1 port map( A1 => n5035, A2 => fromRegsPortxREG_FILE_09xx7x, 
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx7x, ZN 
                           => n4906);
   U5525 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx7x, 
                           B1 => n5036, B2 => fromRegsPortxREG_FILE_03xx7x, ZN 
                           => n4905);
   U5526 : NAND2_X1 port map( A1 => n4903, A2 => fromRegsPortxREG_FILE_05xx7x, 
                           ZN => n4904);
   U5527 : NAND4_X1 port map( A1 => n4907, A2 => n4906, A3 => n4905, A4 => 
                           n4904, ZN => n4911);
   U5528 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx7x, 
                           ZN => n4909);
   U5529 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx7x, A2 => n5072, 
                           ZN => n4908);
   U5530 : NAND2_X1 port map( A1 => n4909, A2 => n4908, ZN => n4910);
   U5531 : AOI21_X1 port map( B1 => n4911, B2 => n4973, A => n4910, ZN => n4912
                           );
   U5532 : NAND2_X1 port map( A1 => n4913, A2 => n4912, ZN => n6377);
   U5533 : INV_X1 port map( A => n6377, ZN => n7463);
   U5534 : OAI22_X1 port map( A1 => n5675, A2 => n6394, B1 => n7364, B2 => 
                           n7463, ZN => n4914);
   U5535 : XOR2_X1 port map( A => n7550, B => n4914, Z => 
                           DP_OP_719J14_125_1055xn61);
   U5536 : AOI22_X1 port map( A1 => n4979, A2 => fromRegsPortxREG_FILE_30xx6x, 
                           B1 => n4978, B2 => fromRegsPortxREG_FILE_28xx6x, ZN 
                           => n4918);
   U5537 : AOI22_X1 port map( A1 => n5013, A2 => fromRegsPortxREG_FILE_24xx6x, 
                           B1 => n5012, B2 => fromRegsPortxREG_FILE_27xx6x, ZN 
                           => n4917);
   U5538 : AOI22_X1 port map( A1 => n5080, A2 => fromRegsPortxREG_FILE_25xx6x, 
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx6x, ZN 
                           => n4916);
   U5539 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx6x, 
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx6x, ZN 
                           => n4915);
   U5540 : NAND4_X1 port map( A1 => n4918, A2 => n4917, A3 => n4916, A4 => 
                           n4915, ZN => n4924);
   U5541 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx6x, 
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx6x, ZN 
                           => n4922);
   U5542 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx6x, 
                           B1 => n5290, B2 => fromRegsPortxREG_FILE_21xx6x, ZN 
                           => n4921);
   U5543 : AOI22_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_19xx6x, 
                           B1 => n5018, B2 => fromRegsPortxREG_FILE_17xx6x, ZN 
                           => n4920);
   U5544 : NAND2_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_22xx6x, 
                           ZN => n4919);
   U5545 : NAND4_X1 port map( A1 => n4922, A2 => n4921, A3 => n4920, A4 => 
                           n4919, ZN => n4923);
   U5546 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4924
                           , A => n4923, ZN => n4930);
   U5547 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx6x, 
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx6x, ZN 
                           => n4929);
   U5548 : AOI22_X1 port map( A1 => n5060, A2 => fromRegsPortxREG_FILE_10xx6x, 
                           B1 => n4994, B2 => fromRegsPortxREG_FILE_11xx6x, ZN 
                           => n4926);
   U5549 : AOI22_X1 port map( A1 => n5306, A2 => fromRegsPortxREG_FILE_13xx6x, 
                           B1 => n4993, B2 => fromRegsPortxREG_FILE_15xx6x, ZN 
                           => n4925);
   U5550 : NAND2_X1 port map( A1 => n4926, A2 => n4925, ZN => n4927);
   U5551 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx6x, B2 => n5129, 
                           A => n4927, ZN => n4928);
   U5552 : OAI211_X1 port map( C1 => n4930, C2 => n5314, A => n4929, B => n4928
                           , ZN => n4931);
   U5553 : NAND2_X1 port map( A1 => n4931, A2 => n5316, ZN => n4942);
   U5554 : AOI22_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx6x, 
                           B1 => n5033, B2 => fromRegsPortxREG_FILE_07xx6x, ZN 
                           => n4936);
   U5555 : AOI22_X1 port map( A1 => n5035, A2 => fromRegsPortxREG_FILE_09xx6x, 
                           B1 => n4965, B2 => fromRegsPortxREG_FILE_04xx6x, ZN 
                           => n4935);
   U5556 : AOI22_X1 port map( A1 => n4932, A2 => fromRegsPortxREG_FILE_08xx6x, 
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx6x, ZN 
                           => n4934);
   U5557 : NAND2_X1 port map( A1 => n5036, A2 => fromRegsPortxREG_FILE_03xx6x, 
                           ZN => n4933);
   U5558 : NAND4_X1 port map( A1 => n4936, A2 => n4935, A3 => n4934, A4 => 
                           n4933, ZN => n4940);
   U5559 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx6x, 
                           ZN => n4938);
   U5560 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx6x, A2 => n5072, 
                           ZN => n4937);
   U5561 : NAND2_X1 port map( A1 => n4938, A2 => n4937, ZN => n4939);
   U5562 : AOI21_X1 port map( B1 => n4940, B2 => n4973, A => n4939, ZN => n4941
                           );
   U5563 : NAND2_X1 port map( A1 => n4942, A2 => n4941, ZN => n6326);
   U5564 : INV_X1 port map( A => n6326, ZN => n7462);
   U5565 : INV_X1 port map( A => add_x_26xBx6x, ZN => n6332);
   U5566 : OAI22_X1 port map( A1 => n5676, A2 => n7462, B1 => n5675, B2 => 
                           n6332, ZN => n4943);
   U5567 : XOR2_X1 port map( A => n5146, B => n4943, Z => 
                           DP_OP_719J14_125_1055xn62);
   U5568 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(25), A2 => n4944,
                           ZN => add_x_26xBx5x);
   U5569 : AOI22_X1 port map( A1 => n4979, A2 => fromRegsPortxREG_FILE_30xx5x, 
                           B1 => n5012, B2 => fromRegsPortxREG_FILE_27xx5x, ZN 
                           => n4950);
   U5570 : AOI22_X1 port map( A1 => n5080, A2 => fromRegsPortxREG_FILE_25xx5x, 
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_24xx5x, ZN 
                           => n4949);
   U5571 : AOI22_X1 port map( A1 => n4945, A2 => fromRegsPortxREG_FILE_29xx5x, 
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx5x, ZN 
                           => n4948);
   U5572 : AOI22_X1 port map( A1 => n4946, A2 => fromRegsPortxREG_FILE_31xx5x, 
                           B1 => n4978, B2 => fromRegsPortxREG_FILE_28xx5x, ZN 
                           => n4947);
   U5573 : NAND4_X1 port map( A1 => n4950, A2 => n4949, A3 => n4948, A4 => 
                           n4947, ZN => n4956);
   U5574 : AOI22_X1 port map( A1 => n4985, A2 => fromRegsPortxREG_FILE_20xx5x, 
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_19xx5x, ZN 
                           => n4954);
   U5575 : AOI22_X1 port map( A1 => n5052, A2 => fromRegsPortxREG_FILE_21xx5x, 
                           B1 => n5018, B2 => fromRegsPortxREG_FILE_17xx5x, ZN 
                           => n4953);
   U5576 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx5x, 
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx5x, ZN 
                           => n4952);
   U5577 : NAND2_X1 port map( A1 => n5289, A2 => fromRegsPortxREG_FILE_22xx5x, 
                           ZN => n4951);
   U5578 : NAND4_X1 port map( A1 => n4954, A2 => n4953, A3 => n4952, A4 => 
                           n4951, ZN => n4955);
   U5579 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4956
                           , A => n4955, ZN => n4963);
   U5580 : AOI22_X1 port map( A1 => n4957, A2 => fromRegsPortxREG_FILE_16xx5x, 
                           B1 => n4993, B2 => fromRegsPortxREG_FILE_15xx5x, ZN 
                           => n4962);
   U5581 : AOI22_X1 port map( A1 => n4995, A2 => fromRegsPortxREG_FILE_14xx5x, 
                           B1 => n4994, B2 => fromRegsPortxREG_FILE_11xx5x, ZN 
                           => n4959);
   U5582 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_12xx5x, 
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx5x, ZN 
                           => n4958);
   U5583 : NAND2_X1 port map( A1 => n4959, A2 => n4958, ZN => n4960);
   U5584 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx5x, B2 => n5060, 
                           A => n4960, ZN => n4961);
   U5585 : OAI211_X1 port map( C1 => n4963, C2 => n5314, A => n4962, B => n4961
                           , ZN => n4964);
   U5586 : NAND2_X1 port map( A1 => n4964, A2 => n5316, ZN => n4976);
   U5587 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx5x, 
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx5x, ZN 
                           => n4969);
   U5588 : AOI22_X1 port map( A1 => n5034, A2 => fromRegsPortxREG_FILE_06xx5x, 
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx5x, ZN 
                           => n4968);
   U5589 : AOI22_X1 port map( A1 => n4965, A2 => fromRegsPortxREG_FILE_04xx5x, 
                           B1 => n5033, B2 => fromRegsPortxREG_FILE_07xx5x, ZN 
                           => n4967);
   U5590 : NAND2_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx5x, 
                           ZN => n4966);
   U5591 : NAND4_X1 port map( A1 => n4969, A2 => n4968, A3 => n4967, A4 => 
                           n4966, ZN => n4974);
   U5592 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx5x, 
                           ZN => n4971);
   U5593 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx5x, A2 => n5072, 
                           ZN => n4970);
   U5594 : NAND2_X1 port map( A1 => n4971, A2 => n4970, ZN => n4972);
   U5595 : AOI21_X1 port map( B1 => n4974, B2 => n4973, A => n4972, ZN => n4975
                           );
   U5596 : NAND2_X1 port map( A1 => n4976, A2 => n4975, ZN => n5402);
   U5597 : INV_X1 port map( A => n5402, ZN => n7461);
   U5598 : INV_X1 port map( A => add_x_26xBx5x, ZN => n6283);
   U5599 : OAI22_X1 port map( A1 => n7461, A2 => n5678, B1 => n5675, B2 => 
                           n6283, ZN => n4977);
   U5600 : XOR2_X1 port map( A => n5146, B => n4977, Z => 
                           DP_OP_719J14_125_1055xn63);
   U5601 : AOI22_X1 port map( A1 => n4979, A2 => fromRegsPortxREG_FILE_30xx4x, 
                           B1 => n4978, B2 => fromRegsPortxREG_FILE_28xx4x, ZN 
                           => n4984);
   U5602 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx4x, 
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_24xx4x, ZN 
                           => n4983);
   U5603 : AOI22_X1 port map( A1 => n5080, A2 => fromRegsPortxREG_FILE_25xx4x, 
                           B1 => n5012, B2 => fromRegsPortxREG_FILE_27xx4x, ZN 
                           => n4982);
   U5604 : AOI22_X1 port map( A1 => n4980, A2 => fromRegsPortxREG_FILE_26xx4x, 
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx4x, ZN 
                           => n4981);
   U5605 : NAND4_X1 port map( A1 => n4984, A2 => n4983, A3 => n4982, A4 => 
                           n4981, ZN => n4992);
   U5606 : AOI22_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx4x, 
                           B1 => n5018, B2 => fromRegsPortxREG_FILE_17xx4x, ZN 
                           => n4990);
   U5607 : AOI22_X1 port map( A1 => n4985, A2 => fromRegsPortxREG_FILE_20xx4x, 
                           B1 => n5291, B2 => fromRegsPortxREG_FILE_23xx4x, ZN 
                           => n4989);
   U5608 : AOI22_X1 port map( A1 => n4986, A2 => fromRegsPortxREG_FILE_18xx4x, 
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_19xx4x, ZN 
                           => n4988);
   U5609 : NAND2_X1 port map( A1 => n5052, A2 => fromRegsPortxREG_FILE_21xx4x, 
                           ZN => n4987);
   U5610 : NAND4_X1 port map( A1 => n4990, A2 => n4989, A3 => n4988, A4 => 
                           n4987, ZN => n4991);
   U5611 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n4992
                           , A => n4991, ZN => n5001);
   U5612 : AOI22_X1 port map( A1 => n5306, A2 => fromRegsPortxREG_FILE_13xx4x, 
                           B1 => n4993, B2 => fromRegsPortxREG_FILE_15xx4x, ZN 
                           => n5000);
   U5613 : AOI22_X1 port map( A1 => n4995, A2 => fromRegsPortxREG_FILE_14xx4x, 
                           B1 => n4994, B2 => fromRegsPortxREG_FILE_11xx4x, ZN 
                           => n4997);
   U5614 : AOI22_X1 port map( A1 => n5129, A2 => fromRegsPortxREG_FILE_12xx4x, 
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx4x, ZN 
                           => n4996);
   U5615 : NAND2_X1 port map( A1 => n4997, A2 => n4996, ZN => n4998);
   U5616 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_10xx4x, B2 => n5302, 
                           A => n4998, ZN => n4999);
   U5617 : OAI211_X1 port map( C1 => n5001, C2 => n5314, A => n5000, B => n4999
                           , ZN => n5010);
   U5618 : AOI22_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx4x, 
                           B1 => n5033, B2 => fromRegsPortxREG_FILE_07xx4x, ZN 
                           => n5005);
   U5619 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx4x, 
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx4x, ZN 
                           => n5004);
   U5620 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx4x, 
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx4x, ZN 
                           => n5003);
   U5621 : NAND2_X1 port map( A1 => n5036, A2 => fromRegsPortxREG_FILE_03xx4x, 
                           ZN => n5002);
   U5622 : NAND4_X1 port map( A1 => n5005, A2 => n5004, A3 => n5003, A4 => 
                           n5002, ZN => n5006);
   U5623 : NAND2_X1 port map( A1 => n5006, A2 => n5334, ZN => n5008);
   U5624 : AOI22_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx4x, 
                           B1 => n5072, B2 => fromRegsPortxREG_FILE_01xx4x, ZN 
                           => n5007);
   U5625 : NAND2_X1 port map( A1 => n5008, A2 => n5007, ZN => n5009);
   U5626 : AOI21_X2 port map( B1 => n5010, B2 => n5316, A => n5009, ZN => n7192
                           );
   U5627 : INV_X1 port map( A => ashr_25xSHx4x, ZN => n7331);
   U5628 : OAI22_X1 port map( A1 => n7192, A2 => n5676, B1 => n5675, B2 => 
                           n7331, ZN => n5011);
   U5629 : XOR2_X1 port map( A => n7550, B => n5011, Z => 
                           DP_OP_719J14_125_1055xn64);
   U5630 : AOI22_X1 port map( A1 => n5013, A2 => fromRegsPortxREG_FILE_24xx3x, 
                           B1 => n5012, B2 => fromRegsPortxREG_FILE_27xx3x, ZN 
                           => n5017);
   U5631 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx3x, 
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx3x, ZN 
                           => n5016);
   U5632 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx3x, 
                           B1 => n5278, B2 => fromRegsPortxREG_FILE_25xx3x, ZN 
                           => n5015);
   U5633 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_26xx3x, 
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx3x, ZN 
                           => n5014);
   U5634 : NAND4_X1 port map( A1 => n5017, A2 => n5016, A3 => n5015, A4 => 
                           n5014, ZN => n5025);
   U5635 : AOI22_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx3x, 
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_19xx3x, ZN 
                           => n5023);
   U5636 : AOI22_X1 port map( A1 => n5052, A2 => fromRegsPortxREG_FILE_21xx3x, 
                           B1 => n5018, B2 => fromRegsPortxREG_FILE_17xx3x, ZN 
                           => n5022);
   U5637 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx3x, 
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx3x, ZN 
                           => n5021);
   U5638 : NAND2_X1 port map( A1 => n5019, A2 => fromRegsPortxREG_FILE_23xx3x, 
                           ZN => n5020);
   U5639 : NAND4_X1 port map( A1 => n5023, A2 => n5022, A3 => n5021, A4 => 
                           n5020, ZN => n5024);
   U5640 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5025
                           , A => n5024, ZN => n5031);
   U5641 : AOI22_X1 port map( A1 => n5306, A2 => fromRegsPortxREG_FILE_13xx3x, 
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx3x, ZN 
                           => n5030);
   U5642 : AOI22_X1 port map( A1 => n5060, A2 => fromRegsPortxREG_FILE_10xx3x, 
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_11xx3x, ZN 
                           => n5027);
   U5643 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx3x, 
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx3x, ZN 
                           => n5026);
   U5644 : NAND2_X1 port map( A1 => n5027, A2 => n5026, ZN => n5028);
   U5645 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx3x, B2 => n5129, 
                           A => n5028, ZN => n5029);
   U5646 : OAI211_X1 port map( C1 => n5031, C2 => n5314, A => n5030, B => n5029
                           , ZN => n5032);
   U5647 : NAND2_X1 port map( A1 => n5032, A2 => n5316, ZN => n5046);
   U5648 : AOI22_X1 port map( A1 => n5324, A2 => fromRegsPortxREG_FILE_08xx3x, 
                           B1 => n5033, B2 => fromRegsPortxREG_FILE_07xx3x, ZN 
                           => n5040);
   U5649 : AOI22_X1 port map( A1 => n5035, A2 => fromRegsPortxREG_FILE_09xx3x, 
                           B1 => n5034, B2 => fromRegsPortxREG_FILE_06xx3x, ZN 
                           => n5039);
   U5650 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx3x, 
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx3x, ZN 
                           => n5038);
   U5651 : NAND2_X1 port map( A1 => n5036, A2 => fromRegsPortxREG_FILE_03xx3x, 
                           ZN => n5037);
   U5652 : NAND4_X1 port map( A1 => n5040, A2 => n5039, A3 => n5038, A4 => 
                           n5037, ZN => n5044);
   U5653 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx3x, 
                           ZN => n5042);
   U5654 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx3x, A2 => n5072, 
                           ZN => n5041);
   U5655 : NAND2_X1 port map( A1 => n5042, A2 => n5041, ZN => n5043);
   U5656 : AOI21_X1 port map( B1 => n5044, B2 => n5334, A => n5043, ZN => n5045
                           );
   U5657 : NAND2_X2 port map( A1 => n5046, A2 => n5045, ZN => n7207);
   U5658 : INV_X2 port map( A => n7207, ZN => n7376);
   U5659 : OAI22_X1 port map( A1 => n7376, A2 => n7364, B1 => n5675, B2 => 
                           intadd_29xBx2x, ZN => n5047);
   U5660 : XOR2_X1 port map( A => n5146, B => n5047, Z => 
                           DP_OP_719J14_125_1055xn65);
   U5661 : AOI22_X1 port map( A1 => n5080, A2 => fromRegsPortxREG_FILE_25xx2x, 
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx2x, ZN 
                           => n5051);
   U5662 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx2x, 
                           B1 => n5280, B2 => fromRegsPortxREG_FILE_29xx2x, ZN 
                           => n5050);
   U5663 : AOI22_X1 port map( A1 => n5282, A2 => fromRegsPortxREG_FILE_24xx2x, 
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx2x, ZN 
                           => n5049);
   U5664 : AOI22_X1 port map( A1 => n5281, A2 => fromRegsPortxREG_FILE_27xx2x, 
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx2x, ZN 
                           => n5048);
   U5665 : NAND4_X1 port map( A1 => n5051, A2 => n5050, A3 => n5049, A4 => 
                           n5048, ZN => n5059);
   U5666 : AOI22_X1 port map( A1 => n5052, A2 => fromRegsPortxREG_FILE_21xx2x, 
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx2x, ZN 
                           => n5057);
   U5667 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx2x, 
                           B1 => n5289, B2 => fromRegsPortxREG_FILE_22xx2x, ZN 
                           => n5056);
   U5668 : AOI22_X1 port map( A1 => n5295, A2 => fromRegsPortxREG_FILE_18xx2x, 
                           B1 => n5053, B2 => fromRegsPortxREG_FILE_19xx2x, ZN 
                           => n5055);
   U5669 : NAND2_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx2x, 
                           ZN => n5054);
   U5670 : NAND4_X1 port map( A1 => n5057, A2 => n5056, A3 => n5055, A4 => 
                           n5054, ZN => n5058);
   U5671 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5059
                           , A => n5058, ZN => n5066);
   U5672 : AOI22_X1 port map( A1 => n5303, A2 => fromRegsPortxREG_FILE_12xx2x, 
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx2x, ZN 
                           => n5065);
   U5673 : AOI22_X1 port map( A1 => n5060, A2 => fromRegsPortxREG_FILE_10xx2x, 
                           B1 => n5304, B2 => fromRegsPortxREG_FILE_14xx2x, ZN 
                           => n5062);
   U5674 : AOI22_X1 port map( A1 => n5311, A2 => fromRegsPortxREG_FILE_16xx2x, 
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx2x, ZN 
                           => n5061);
   U5675 : NAND2_X1 port map( A1 => n5062, A2 => n5061, ZN => n5063);
   U5676 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_11xx2x, B2 => n5305, 
                           A => n5063, ZN => n5064);
   U5677 : OAI211_X1 port map( C1 => n5066, C2 => n5314, A => n5065, B => n5064
                           , ZN => n5067);
   U5678 : NAND2_X1 port map( A1 => n5067, A2 => n5316, ZN => n5078);
   U5679 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx2x, 
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx2x, ZN 
                           => n5071);
   U5680 : AOI22_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx2x, 
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx2x, ZN 
                           => n5070);
   U5681 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx2x, 
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx2x, ZN 
                           => n5069);
   U5682 : NAND2_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx2x, 
                           ZN => n5068);
   U5683 : NAND4_X1 port map( A1 => n5071, A2 => n5070, A3 => n5069, A4 => 
                           n5068, ZN => n5076);
   U5684 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx2x, 
                           ZN => n5074);
   U5685 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx2x, A2 => n5072, 
                           ZN => n5073);
   U5686 : NAND2_X1 port map( A1 => n5074, A2 => n5073, ZN => n5075);
   U5687 : AOI21_X1 port map( B1 => n5076, B2 => n5334, A => n5075, ZN => n5077
                           );
   U5688 : NAND2_X1 port map( A1 => n5078, A2 => n5077, ZN => n6900);
   U5689 : CLKBUF_X1 port map( A => n6900, Z => n7309);
   U5690 : OAI22_X1 port map( A1 => n7311, A2 => n5678, B1 => n5675, B2 => 
                           intadd_29xBx1x, ZN => n5079);
   U5691 : XOR2_X1 port map( A => n7550, B => n5079, Z => 
                           DP_OP_719J14_125_1055xn66);
   U5692 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx1x, 
                           B1 => n5281, B2 => fromRegsPortxREG_FILE_27xx1x, ZN 
                           => n5084);
   U5693 : AOI22_X1 port map( A1 => n5279, A2 => fromRegsPortxREG_FILE_26xx1x, 
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx1x, ZN 
                           => n5083);
   U5694 : AOI22_X1 port map( A1 => n5080, A2 => fromRegsPortxREG_FILE_25xx1x, 
                           B1 => n5282, B2 => fromRegsPortxREG_FILE_24xx1x, ZN 
                           => n5082);
   U5695 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx1x, 
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx1x, ZN 
                           => n5081);
   U5696 : NAND4_X1 port map( A1 => n5084, A2 => n5083, A3 => n5082, A4 => 
                           n5081, ZN => n5090);
   U5697 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx1x, 
                           B1 => n5293, B2 => fromRegsPortxREG_FILE_19xx1x, ZN 
                           => n5088);
   U5698 : AOI22_X1 port map( A1 => n5290, A2 => fromRegsPortxREG_FILE_21xx1x, 
                           B1 => n5119, B2 => fromRegsPortxREG_FILE_22xx1x, ZN 
                           => n5087);
   U5699 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx1x, 
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx1x, ZN 
                           => n5086);
   U5700 : NAND2_X1 port map( A1 => n5295, A2 => fromRegsPortxREG_FILE_18xx1x, 
                           ZN => n5085);
   U5701 : NAND4_X1 port map( A1 => n5088, A2 => n5087, A3 => n5086, A4 => 
                           n5085, ZN => n5089);
   U5702 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5090
                           , A => n5089, ZN => n5097);
   U5703 : AOI22_X1 port map( A1 => n5305, A2 => fromRegsPortxREG_FILE_11xx1x, 
                           B1 => n5091, B2 => fromRegsPortxREG_FILE_13xx1x, ZN 
                           => n5096);
   U5704 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx1x, 
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx1x, ZN 
                           => n5093);
   U5705 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx1x, 
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx1x, ZN 
                           => n5092);
   U5706 : NAND2_X1 port map( A1 => n5093, A2 => n5092, ZN => n5094);
   U5707 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx1x, B2 => n5129, 
                           A => n5094, ZN => n5095);
   U5708 : OAI211_X1 port map( C1 => n5097, C2 => n5314, A => n5096, B => n5095
                           , ZN => n5098);
   U5709 : NAND2_X1 port map( A1 => n5098, A2 => n5133, ZN => n5108);
   U5710 : AOI22_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx1x, 
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx1x, ZN 
                           => n5102);
   U5711 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx1x, 
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx1x, ZN 
                           => n5101);
   U5712 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx1x, 
                           B1 => n5319, B2 => fromRegsPortxREG_FILE_06xx1x, ZN 
                           => n5100);
   U5713 : NAND2_X1 port map( A1 => n5323, A2 => fromRegsPortxREG_FILE_05xx1x, 
                           ZN => n5099);
   U5714 : NAND4_X1 port map( A1 => n5102, A2 => n5101, A3 => n5100, A4 => 
                           n5099, ZN => n5106);
   U5715 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx1x, 
                           ZN => n5104);
   U5716 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx1x, A2 => n5330, 
                           ZN => n5103);
   U5717 : NAND2_X1 port map( A1 => n5104, A2 => n5103, ZN => n5105);
   U5718 : AOI21_X1 port map( B1 => n5106, B2 => n5334, A => n5105, ZN => n5107
                           );
   U5719 : NAND2_X2 port map( A1 => n5108, A2 => n5107, ZN => n7402);
   U5720 : INV_X2 port map( A => n7402, ZN => n7304);
   U5721 : OAI22_X1 port map( A1 => intadd_29xBx0x, A2 => n5675, B1 => n7364, 
                           B2 => n7304, ZN => n5109);
   U5722 : XOR2_X1 port map( A => n7550, B => n5109, Z => 
                           DP_OP_719J14_125_1055xn67);
   U5723 : NAND2_X1 port map( A1 => n7460, A2 => fromMemoryPortxLOADEDDATAx(7),
                           ZN => n5114);
   U5724 : AND2_X1 port map( A1 => n7452, A2 => n5110, ZN => n5111);
   U5725 : NAND2_X1 port map( A1 => n5715, A2 => n5111, ZN => n5112);
   U5726 : NAND2_X1 port map( A1 => n5112, A2 => fromMemoryPortxLOADEDDATAx(20)
                           , ZN => n5113);
   U5727 : NAND2_X2 port map( A1 => n5114, A2 => n5113, ZN => n7412);
   U5728 : INV_X1 port map( A => n7412, ZN => n7333);
   U5729 : AOI22_X1 port map( A1 => n5281, A2 => fromRegsPortxREG_FILE_27xx0x, 
                           B1 => n5283, B2 => fromRegsPortxREG_FILE_28xx0x, ZN 
                           => n5118);
   U5730 : AOI22_X1 port map( A1 => n5280, A2 => fromRegsPortxREG_FILE_29xx0x, 
                           B1 => n5279, B2 => fromRegsPortxREG_FILE_26xx0x, ZN 
                           => n5117);
   U5731 : AOI22_X1 port map( A1 => n5277, A2 => fromRegsPortxREG_FILE_30xx0x, 
                           B1 => n5278, B2 => fromRegsPortxREG_FILE_25xx0x, ZN 
                           => n5116);
   U5732 : AOI22_X1 port map( A1 => n5282, A2 => fromRegsPortxREG_FILE_24xx0x, 
                           B1 => n5284, B2 => fromRegsPortxREG_FILE_31xx0x, ZN 
                           => n5115);
   U5733 : NAND4_X1 port map( A1 => n5118, A2 => n5117, A3 => n5116, A4 => 
                           n5115, ZN => n5125);
   U5734 : AOI22_X1 port map( A1 => n5119, A2 => fromRegsPortxREG_FILE_22xx0x, 
                           B1 => n5295, B2 => fromRegsPortxREG_FILE_18xx0x, ZN 
                           => n5123);
   U5735 : AOI22_X1 port map( A1 => n5291, A2 => fromRegsPortxREG_FILE_23xx0x, 
                           B1 => n5290, B2 => fromRegsPortxREG_FILE_21xx0x, ZN 
                           => n5122);
   U5736 : AOI22_X1 port map( A1 => n5292, A2 => fromRegsPortxREG_FILE_20xx0x, 
                           B1 => n5294, B2 => fromRegsPortxREG_FILE_17xx0x, ZN 
                           => n5121);
   U5737 : NAND2_X1 port map( A1 => n5293, A2 => fromRegsPortxREG_FILE_19xx0x, 
                           ZN => n5120);
   U5738 : NAND4_X1 port map( A1 => n5123, A2 => n5122, A3 => n5121, A4 => 
                           n5120, ZN => n5124);
   U5739 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5125
                           , A => n5124, ZN => n5132);
   U5740 : AOI22_X1 port map( A1 => n5306, A2 => fromRegsPortxREG_FILE_13xx0x, 
                           B1 => n5307, B2 => fromRegsPortxREG_FILE_15xx0x, ZN 
                           => n5131);
   U5741 : AOI22_X1 port map( A1 => n5302, A2 => fromRegsPortxREG_FILE_10xx0x, 
                           B1 => n5305, B2 => fromRegsPortxREG_FILE_11xx0x, ZN 
                           => n5127);
   U5742 : AOI22_X1 port map( A1 => n5304, A2 => fromRegsPortxREG_FILE_14xx0x, 
                           B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx0x, ZN 
                           => n5126);
   U5743 : NAND2_X1 port map( A1 => n5127, A2 => n5126, ZN => n5128);
   U5744 : AOI21_X1 port map( B1 => fromRegsPortxREG_FILE_12xx0x, B2 => n5129, 
                           A => n5128, ZN => n5130);
   U5745 : OAI211_X1 port map( C1 => n5132, C2 => n7071, A => n5131, B => n5130
                           , ZN => n5134);
   U5746 : NAND2_X1 port map( A1 => n5134, A2 => n5133, ZN => n5144);
   U5747 : AOI22_X1 port map( A1 => n5318, A2 => fromRegsPortxREG_FILE_03xx0x, 
                           B1 => n5324, B2 => fromRegsPortxREG_FILE_08xx0x, ZN 
                           => n5138);
   U5748 : AOI22_X1 port map( A1 => n5319, A2 => fromRegsPortxREG_FILE_06xx0x, 
                           B1 => n5323, B2 => fromRegsPortxREG_FILE_05xx0x, ZN 
                           => n5137);
   U5749 : AOI22_X1 port map( A1 => n5320, A2 => fromRegsPortxREG_FILE_04xx0x, 
                           B1 => n5322, B2 => fromRegsPortxREG_FILE_07xx0x, ZN 
                           => n5136);
   U5750 : NAND2_X1 port map( A1 => n5321, A2 => fromRegsPortxREG_FILE_09xx0x, 
                           ZN => n5135);
   U5751 : NAND4_X1 port map( A1 => n5138, A2 => n5137, A3 => n5136, A4 => 
                           n5135, ZN => n5142);
   U5752 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx0x, 
                           ZN => n5140);
   U5753 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx0x, A2 => n5330, 
                           ZN => n5139);
   U5754 : NAND2_X1 port map( A1 => n5140, A2 => n5139, ZN => n5141);
   U5755 : AOI21_X1 port map( B1 => n5142, B2 => n5334, A => n5141, ZN => n5143
                           );
   U5756 : NAND2_X1 port map( A1 => n5144, A2 => n5143, ZN => n7086);
   U5757 : CLKBUF_X1 port map( A => n7086, Z => n7267);
   U5758 : OAI22_X1 port map( A1 => n5674, A2 => n7333, B1 => n5676, B2 => 
                           n7209, ZN => n5145);
   U5759 : XOR2_X1 port map( A => n5146, B => n5145, Z => 
                           DP_OP_719J14_125_1055xn68);
   U5760 : XOR2_X1 port map( A => n7551, B => n7321, Z => 
                           DP_OP_679J14_122_3096xn38);
   U5761 : XOR2_X1 port map( A => n7551, B => n7252, Z => 
                           DP_OP_679J14_122_3096xn39);
   U5762 : XOR2_X1 port map( A => n7551, B => n7242, Z => 
                           DP_OP_679J14_122_3096xn40);
   U5763 : XOR2_X1 port map( A => n7551, B => n7183, Z => 
                           DP_OP_679J14_122_3096xn41);
   U5764 : XOR2_X1 port map( A => n7551, B => n7120, Z => 
                           DP_OP_679J14_122_3096xn42);
   U5765 : XOR2_X1 port map( A => n7551, B => n7097, Z => 
                           DP_OP_679J14_122_3096xn43);
   U5766 : XOR2_X1 port map( A => n7551, B => n7053, Z => 
                           DP_OP_679J14_122_3096xn44);
   U5767 : XOR2_X1 port map( A => n5680, B => n7009, Z => 
                           DP_OP_679J14_122_3096xn45);
   U5768 : XOR2_X1 port map( A => n5680, B => n6958, Z => 
                           DP_OP_679J14_122_3096xn46);
   U5769 : XOR2_X1 port map( A => n5680, B => n5720, Z => 
                           DP_OP_679J14_122_3096xn47);
   U5770 : XOR2_X1 port map( A => n5680, B => n6933, Z => 
                           DP_OP_679J14_122_3096xn48);
   U5771 : XOR2_X1 port map( A => n5680, B => n6888, Z => 
                           DP_OP_679J14_122_3096xn49);
   U5772 : XOR2_X1 port map( A => n5680, B => n6861, Z => 
                           DP_OP_679J14_122_3096xn50);
   U5773 : XOR2_X1 port map( A => n7551, B => n6806, Z => 
                           DP_OP_679J14_122_3096xn51);
   U5774 : XOR2_X1 port map( A => n7551, B => n6777, Z => 
                           DP_OP_679J14_122_3096xn52);
   U5775 : XOR2_X1 port map( A => n7551, B => n6739, Z => 
                           DP_OP_679J14_122_3096xn53);
   U5776 : XOR2_X1 port map( A => n7551, B => n6693, Z => 
                           DP_OP_679J14_122_3096xn54);
   U5777 : XOR2_X1 port map( A => n7551, B => n6669, Z => 
                           DP_OP_679J14_122_3096xn55);
   U5778 : XOR2_X1 port map( A => n7551, B => n6626, Z => 
                           DP_OP_679J14_122_3096xn56);
   U5779 : XOR2_X1 port map( A => n7551, B => n6553, Z => 
                           DP_OP_679J14_122_3096xn57);
   U5780 : XOR2_X1 port map( A => n7551, B => n6530, Z => 
                           DP_OP_679J14_122_3096xn58);
   U5781 : XOR2_X1 port map( A => n7551, B => n6480, Z => 
                           DP_OP_679J14_122_3096xn59);
   U5782 : XOR2_X1 port map( A => n7551, B => n6421, Z => 
                           DP_OP_679J14_122_3096xn60);
   U5783 : XOR2_X1 port map( A => n7551, B => n6377, Z => 
                           DP_OP_679J14_122_3096xn61);
   U5784 : XOR2_X1 port map( A => n7551, B => n6326, Z => 
                           DP_OP_679J14_122_3096xn62);
   U5785 : XOR2_X1 port map( A => n7551, B => n5402, Z => 
                           DP_OP_679J14_122_3096xn63);
   U5786 : INV_X1 port map( A => n7192, ZN => n7349);
   U5787 : XOR2_X1 port map( A => n7551, B => n7349, Z => 
                           DP_OP_679J14_122_3096xn64);
   U5788 : XOR2_X1 port map( A => n7551, B => n7207, Z => 
                           DP_OP_679J14_122_3096xn65);
   U5789 : CLKBUF_X1 port map( A => n6900, Z => n6110);
   U5790 : XOR2_X1 port map( A => n7551, B => n6110, Z => 
                           DP_OP_679J14_122_3096xn66);
   U5791 : XOR2_X1 port map( A => n7551, B => n5711, Z => 
                           DP_OP_679J14_122_3096xn67);
   U5792 : CLKBUF_X1 port map( A => n7086, Z => n7399);
   U5793 : XOR2_X1 port map( A => n7551, B => n7399, Z => 
                           DP_OP_679J14_122_3096xn68);
   U5794 : INV_X1 port map( A => ashr_25xAx1x, ZN => intadd_29xAx0x);
   U5795 : INV_X1 port map( A => ashr_25xAx30x, ZN => intadd_28xAx2x);
   U5796 : INV_X1 port map( A => ashr_25xAx29x, ZN => intadd_28xAx1x);
   U5797 : INV_X1 port map( A => ashr_25xAx28x, ZN => intadd_28xAx0x);
   U5798 : AOI22_X1 port map( A1 => n5251, A2 => fromRegsPortxREG_FILE_17xx14x,
                           B1 => n5266, B2 => fromRegsPortxREG_FILE_24xx14x, ZN
                           => n5151);
   U5799 : AOI22_X1 port map( A1 => n5147, A2 => fromRegsPortxREG_FILE_08xx14x,
                           B1 => n5261, B2 => fromRegsPortxREG_FILE_27xx14x, ZN
                           => n5150);
   U5800 : NAND2_X1 port map( A1 => n5356, A2 => fromRegsPortxREG_FILE_12xx14x,
                           ZN => n5149);
   U5801 : AOI22_X1 port map( A1 => n5267, A2 => fromRegsPortxREG_FILE_25xx14x,
                           B1 => n5339, B2 => fromRegsPortxREG_FILE_30xx14x, ZN
                           => n5148);
   U5802 : AND4_X1 port map( A1 => n5151, A2 => n5150, A3 => n5149, A4 => n5148
                           , ZN => n5175);
   U5803 : AOI22_X1 port map( A1 => n5365, A2 => fromRegsPortxREG_FILE_26xx14x,
                           B1 => n5152, B2 => fromRegsPortxREG_FILE_14xx14x, ZN
                           => n5157);
   U5804 : AOI22_X1 port map( A1 => n5259, A2 => fromRegsPortxREG_FILE_21xx14x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx14x, ZN
                           => n5156);
   U5805 : AOI22_X1 port map( A1 => n5176, A2 => fromRegsPortxREG_FILE_03xx14x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx14x, ZN
                           => n5155);
   U5806 : AOI22_X1 port map( A1 => n5153, A2 => fromRegsPortxREG_FILE_29xx14x,
                           B1 => n5211, B2 => fromRegsPortxREG_FILE_23xx14x, ZN
                           => n5154);
   U5807 : AND4_X1 port map( A1 => n5157, A2 => n5156, A3 => n5155, A4 => n5154
                           , ZN => n5174);
   U5808 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx14x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_11xx14x, ZN
                           => n5164);
   U5809 : AOI22_X1 port map( A1 => n5158, A2 => fromRegsPortxREG_FILE_31xx14x,
                           B1 => n5357, B2 => fromRegsPortxREG_FILE_04xx14x, ZN
                           => n5163);
   U5810 : AOI22_X1 port map( A1 => n5159, A2 => fromRegsPortxREG_FILE_28xx14x,
                           B1 => n5225, B2 => fromRegsPortxREG_FILE_22xx14x, ZN
                           => n5162);
   U5811 : AOI22_X1 port map( A1 => n5197, A2 => fromRegsPortxREG_FILE_06xx14x,
                           B1 => n5160, B2 => fromRegsPortxREG_FILE_15xx14x, ZN
                           => n5161);
   U5812 : AND4_X1 port map( A1 => n5164, A2 => n5163, A3 => n5162, A4 => n5161
                           , ZN => n5173);
   U5813 : AOI22_X1 port map( A1 => n5165, A2 => fromRegsPortxREG_FILE_20xx14x,
                           B1 => n5220, B2 => fromRegsPortxREG_FILE_05xx14x, ZN
                           => n5171);
   U5814 : AOI22_X1 port map( A1 => n5367, A2 => fromRegsPortxREG_FILE_19xx14x,
                           B1 => n5166, B2 => fromRegsPortxREG_FILE_18xx14x, ZN
                           => n5170);
   U5815 : AOI22_X1 port map( A1 => n5260, A2 => fromRegsPortxREG_FILE_02xx14x,
                           B1 => n5167, B2 => fromRegsPortxREG_FILE_10xx14x, ZN
                           => n5169);
   U5816 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx14x,
                           B1 => n5230, B2 => fromRegsPortxREG_FILE_07xx14x, ZN
                           => n5168);
   U5817 : AND4_X1 port map( A1 => n5171, A2 => n5170, A3 => n5169, A4 => n5168
                           , ZN => n5172);
   U5818 : NAND4_X1 port map( A1 => n5175, A2 => n5174, A3 => n5173, A4 => 
                           n5172, ZN => ashr_25xAx14x);
   U5819 : INV_X1 port map( A => ashr_25xAx14x, ZN => intadd_27xAx3x);
   U5820 : INV_X1 port map( A => ashr_25xAx13x, ZN => intadd_27xAx2x);
   U5821 : INV_X1 port map( A => ashr_25xAx24x, ZN => intadd_26xAx7x);
   U5822 : INV_X1 port map( A => ashr_25xAx23x, ZN => intadd_26xAx6x);
   U5823 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx22x,
                           B1 => n5176, B2 => fromRegsPortxREG_FILE_03xx22x, ZN
                           => n5180);
   U5824 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx22x,
                           B1 => n5220, B2 => fromRegsPortxREG_FILE_05xx22x, ZN
                           => n5179);
   U5825 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx22x,
                           B1 => n5367, B2 => fromRegsPortxREG_FILE_19xx22x, ZN
                           => n5178);
   U5826 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx22x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx22x, ZN
                           => n5177);
   U5827 : AND4_X1 port map( A1 => n5180, A2 => n5179, A3 => n5178, A4 => n5177
                           , ZN => n5196);
   U5828 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx22x,
                           B1 => n5345, B2 => fromRegsPortxREG_FILE_16xx22x, ZN
                           => n5184);
   U5829 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx22x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_17xx22x, ZN
                           => n5183);
   U5830 : AOI22_X1 port map( A1 => n5267, A2 => fromRegsPortxREG_FILE_25xx22x,
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_28xx22x, ZN
                           => n5182);
   U5831 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_02xx22x,
                           B1 => n5356, B2 => fromRegsPortxREG_FILE_12xx22x, ZN
                           => n5181);
   U5832 : AND4_X1 port map( A1 => n5184, A2 => n5183, A3 => n5182, A4 => n5181
                           , ZN => n5195);
   U5833 : AOI22_X1 port map( A1 => n5225, A2 => fromRegsPortxREG_FILE_22xx22x,
                           B1 => n5246, B2 => fromRegsPortxREG_FILE_13xx22x, ZN
                           => n5188);
   U5834 : AOI22_X1 port map( A1 => n5376, A2 => fromRegsPortxREG_FILE_24xx22x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx22x, ZN
                           => n5187);
   U5835 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx22x,
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx22x, ZN
                           => n5186);
   U5836 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_11xx22x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx22x, ZN
                           => n5185);
   U5837 : AND4_X1 port map( A1 => n5188, A2 => n5187, A3 => n5186, A4 => n5185
                           , ZN => n5194);
   U5838 : AOI22_X1 port map( A1 => n5379, A2 => fromRegsPortxREG_FILE_31xx22x,
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx22x, ZN
                           => n5192);
   U5839 : AOI22_X1 port map( A1 => n5357, A2 => fromRegsPortxREG_FILE_04xx22x,
                           B1 => n5365, B2 => fromRegsPortxREG_FILE_26xx22x, ZN
                           => n5191);
   U5840 : AOI22_X1 port map( A1 => n5235, A2 => fromRegsPortxREG_FILE_09xx22x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx22x, ZN
                           => n5190);
   U5841 : NAND2_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx22x,
                           ZN => n5189);
   U5842 : AND4_X1 port map( A1 => n5192, A2 => n5191, A3 => n5190, A4 => n5189
                           , ZN => n5193);
   U5843 : NAND4_X1 port map( A1 => n5196, A2 => n5195, A3 => n5194, A4 => 
                           n5193, ZN => ashr_25xAx22x);
   U5844 : INV_X1 port map( A => ashr_25xAx22x, ZN => intadd_26xAx5x);
   U5845 : INV_X1 port map( A => ashr_25xAx21x, ZN => intadd_26xAx4x);
   U5846 : INV_X1 port map( A => ashr_25xAx20x, ZN => intadd_26xAx3x);
   U5847 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx19x,
                           B1 => n5197, B2 => fromRegsPortxREG_FILE_06xx19x, ZN
                           => n5201);
   U5848 : AOI22_X1 port map( A1 => n5379, A2 => fromRegsPortxREG_FILE_31xx19x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx19x, ZN
                           => n5200);
   U5849 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_11xx19x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx19x, ZN
                           => n5199);
   U5850 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_28xx19x,
                           B1 => n5244, B2 => fromRegsPortxREG_FILE_19xx19x, ZN
                           => n5198);
   U5851 : AND4_X1 port map( A1 => n5201, A2 => n5200, A3 => n5199, A4 => n5198
                           , ZN => n5219);
   U5852 : AOI22_X1 port map( A1 => n5261, A2 => fromRegsPortxREG_FILE_27xx19x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx19x, ZN
                           => n5206);
   U5853 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx19x,
                           B1 => n5251, B2 => fromRegsPortxREG_FILE_17xx19x, ZN
                           => n5205);
   U5854 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx19x,
                           B1 => n5252, B2 => fromRegsPortxREG_FILE_04xx19x, ZN
                           => n5204);
   U5855 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx19x,
                           B1 => n5202, B2 => fromRegsPortxREG_FILE_12xx19x, ZN
                           => n5203);
   U5856 : AND4_X1 port map( A1 => n5206, A2 => n5205, A3 => n5204, A4 => n5203
                           , ZN => n5218);
   U5857 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_02xx19x,
                           B1 => n5246, B2 => fromRegsPortxREG_FILE_13xx19x, ZN
                           => n5210);
   U5858 : AOI22_X1 port map( A1 => n5365, A2 => fromRegsPortxREG_FILE_26xx19x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx19x, ZN
                           => n5209);
   U5859 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx19x,
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx19x, ZN
                           => n5208);
   U5860 : AOI22_X1 port map( A1 => n5267, A2 => fromRegsPortxREG_FILE_25xx19x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx19x, ZN
                           => n5207);
   U5861 : AND4_X1 port map( A1 => n5210, A2 => n5209, A3 => n5208, A4 => n5207
                           , ZN => n5217);
   U5862 : AOI22_X1 port map( A1 => n5354, A2 => fromRegsPortxREG_FILE_20xx19x,
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx19x, ZN
                           => n5215);
   U5863 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx19x,
                           B1 => n5266, B2 => fromRegsPortxREG_FILE_24xx19x, ZN
                           => n5214);
   U5864 : NAND2_X1 port map( A1 => n5211, A2 => fromRegsPortxREG_FILE_23xx19x,
                           ZN => n5213);
   U5865 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx19x,
                           B1 => n5268, B2 => fromRegsPortxREG_FILE_30xx19x, ZN
                           => n5212);
   U5866 : AND4_X1 port map( A1 => n5215, A2 => n5214, A3 => n5213, A4 => n5212
                           , ZN => n5216);
   U5867 : NAND4_X1 port map( A1 => n5219, A2 => n5218, A3 => n5217, A4 => 
                           n5216, ZN => ashr_25xAx19x);
   U5868 : INV_X1 port map( A => ashr_25xAx19x, ZN => intadd_26xAx2x);
   U5869 : AOI22_X1 port map( A1 => n5267, A2 => fromRegsPortxREG_FILE_25xx18x,
                           B1 => n5220, B2 => fromRegsPortxREG_FILE_05xx18x, ZN
                           => n5224);
   U5870 : AOI22_X1 port map( A1 => n5379, A2 => fromRegsPortxREG_FILE_31xx18x,
                           B1 => n5375, B2 => fromRegsPortxREG_FILE_02xx18x, ZN
                           => n5223);
   U5871 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx18x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx18x, ZN
                           => n5222);
   U5872 : AOI22_X1 port map( A1 => n5350, A2 => fromRegsPortxREG_FILE_17xx18x,
                           B1 => n5369, B2 => fromRegsPortxREG_FILE_10xx18x, ZN
                           => n5221);
   U5873 : AND4_X1 port map( A1 => n5224, A2 => n5223, A3 => n5222, A4 => n5221
                           , ZN => n5243);
   U5874 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx18x,
                           B1 => n5356, B2 => fromRegsPortxREG_FILE_12xx18x, ZN
                           => n5229);
   U5875 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx18x,
                           B1 => n5225, B2 => fromRegsPortxREG_FILE_22xx18x, ZN
                           => n5228);
   U5876 : AOI22_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_01xx18x,
                           B1 => n5354, B2 => fromRegsPortxREG_FILE_20xx18x, ZN
                           => n5227);
   U5877 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx18x,
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_28xx18x, ZN
                           => n5226);
   U5878 : AND4_X1 port map( A1 => n5229, A2 => n5228, A3 => n5227, A4 => n5226
                           , ZN => n5242);
   U5879 : AOI22_X1 port map( A1 => n5367, A2 => fromRegsPortxREG_FILE_19xx18x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx18x, ZN
                           => n5234);
   U5880 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx18x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx18x, ZN
                           => n5233);
   U5881 : AOI22_X1 port map( A1 => n5230, A2 => fromRegsPortxREG_FILE_07xx18x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_21xx18x, ZN
                           => n5232);
   U5882 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx18x,
                           B1 => n5341, B2 => fromRegsPortxREG_FILE_11xx18x, ZN
                           => n5231);
   U5883 : AND4_X1 port map( A1 => n5234, A2 => n5233, A3 => n5232, A4 => n5231
                           , ZN => n5241);
   U5884 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx18x,
                           B1 => n5266, B2 => fromRegsPortxREG_FILE_24xx18x, ZN
                           => n5239);
   U5885 : AOI22_X1 port map( A1 => n5252, A2 => fromRegsPortxREG_FILE_04xx18x,
                           B1 => n5353, B2 => fromRegsPortxREG_FILE_27xx18x, ZN
                           => n5238);
   U5886 : AOI22_X1 port map( A1 => n5235, A2 => fromRegsPortxREG_FILE_09xx18x,
                           B1 => n5245, B2 => fromRegsPortxREG_FILE_26xx18x, ZN
                           => n5237);
   U5887 : NAND2_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx18x,
                           ZN => n5236);
   U5888 : AND4_X1 port map( A1 => n5239, A2 => n5238, A3 => n5237, A4 => n5236
                           , ZN => n5240);
   U5889 : NAND4_X1 port map( A1 => n5243, A2 => n5242, A3 => n5241, A4 => 
                           n5240, ZN => ashr_25xAx18x);
   U5890 : INV_X1 port map( A => ashr_25xAx18x, ZN => intadd_26xAx1x);
   U5891 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx17x,
                           B1 => n5244, B2 => fromRegsPortxREG_FILE_19xx17x, ZN
                           => n5250);
   U5892 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx17x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx17x, ZN
                           => n5249);
   U5893 : AOI22_X1 port map( A1 => n5245, A2 => fromRegsPortxREG_FILE_26xx17x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx17x, ZN
                           => n5248);
   U5894 : AOI22_X1 port map( A1 => n5356, A2 => fromRegsPortxREG_FILE_12xx17x,
                           B1 => n5246, B2 => fromRegsPortxREG_FILE_13xx17x, ZN
                           => n5247);
   U5895 : AND4_X1 port map( A1 => n5250, A2 => n5249, A3 => n5248, A4 => n5247
                           , ZN => n5276);
   U5896 : AOI22_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx17x,
                           B1 => n5251, B2 => fromRegsPortxREG_FILE_17xx17x, ZN
                           => n5257);
   U5897 : AOI22_X1 port map( A1 => n5379, A2 => fromRegsPortxREG_FILE_31xx17x,
                           B1 => n5252, B2 => fromRegsPortxREG_FILE_04xx17x, ZN
                           => n5256);
   U5898 : AOI22_X1 port map( A1 => n5253, A2 => fromRegsPortxREG_FILE_01xx17x,
                           B1 => n5354, B2 => fromRegsPortxREG_FILE_20xx17x, ZN
                           => n5255);
   U5899 : AOI22_X1 port map( A1 => n5374, A2 => fromRegsPortxREG_FILE_05xx17x,
                           B1 => n5377, B2 => fromRegsPortxREG_FILE_28xx17x, ZN
                           => n5254);
   U5900 : AND4_X1 port map( A1 => n5257, A2 => n5256, A3 => n5255, A4 => n5254
                           , ZN => n5275);
   U5901 : AOI22_X1 port map( A1 => n5338, A2 => fromRegsPortxREG_FILE_23xx17x,
                           B1 => n5258, B2 => fromRegsPortxREG_FILE_11xx17x, ZN
                           => n5265);
   U5902 : AOI22_X1 port map( A1 => n5260, A2 => fromRegsPortxREG_FILE_02xx17x,
                           B1 => n5259, B2 => fromRegsPortxREG_FILE_21xx17x, ZN
                           => n5264);
   U5903 : AOI22_X1 port map( A1 => n5261, A2 => fromRegsPortxREG_FILE_27xx17x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx17x, ZN
                           => n5263);
   U5904 : AOI22_X1 port map( A1 => n5362, A2 => fromRegsPortxREG_FILE_06xx17x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx17x, ZN
                           => n5262);
   U5905 : AND4_X1 port map( A1 => n5265, A2 => n5264, A3 => n5263, A4 => n5262
                           , ZN => n5274);
   U5906 : AOI22_X1 port map( A1 => n5344, A2 => fromRegsPortxREG_FILE_15xx17x,
                           B1 => n5343, B2 => fromRegsPortxREG_FILE_07xx17x, ZN
                           => n5272);
   U5907 : AOI22_X1 port map( A1 => n5267, A2 => fromRegsPortxREG_FILE_25xx17x,
                           B1 => n5266, B2 => fromRegsPortxREG_FILE_24xx17x, ZN
                           => n5271);
   U5908 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx17x,
                           B1 => n5268, B2 => fromRegsPortxREG_FILE_30xx17x, ZN
                           => n5270);
   U5909 : NAND2_X1 port map( A1 => n5369, A2 => fromRegsPortxREG_FILE_10xx17x,
                           ZN => n5269);
   U5910 : AND4_X1 port map( A1 => n5272, A2 => n5271, A3 => n5270, A4 => n5269
                           , ZN => n5273);
   U5911 : NAND4_X1 port map( A1 => n5276, A2 => n5275, A3 => n5274, A4 => 
                           n5273, ZN => ashr_25xAx17x);
   U5912 : INV_X1 port map( A => ashr_25xAx17x, ZN => intadd_26xAx0x);
   U5913 : NAND2_X1 port map( A1 => n7538, A2 => n7509, ZN => n5952);
   U5914 : INV_X1 port map( A => n5952, ZN => n5827);
   U5915 : INV_X1 port map( A => n5827, ZN => n5936);
   U5916 : NAND2_X1 port map( A1 => n5739, A2 => n7535, ZN => n5740);
   U5917 : NOR4_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(2), A2 => n5936, 
                           A3 => n6361, A4 => n5740, ZN => n5443);
   U5918 : AND2_X1 port map( A1 => n5443, A2 => n5741, ZN => n5659);
   U5919 : INV_X1 port map( A => n5659, ZN => n5625);
   U5920 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_25xx31x, A2 => n5278,
                           B1 => fromRegsPortxREG_FILE_30xx31x, B2 => n5277, ZN
                           => n5288);
   U5921 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_29xx31x, A2 => n5280,
                           B1 => fromRegsPortxREG_FILE_26xx31x, B2 => n5279, ZN
                           => n5287);
   U5922 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_24xx31x, A2 => n5282,
                           B1 => fromRegsPortxREG_FILE_27xx31x, B2 => n5281, ZN
                           => n5286);
   U5923 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_31xx31x, A2 => n5284,
                           B1 => fromRegsPortxREG_FILE_28xx31x, B2 => n5283, ZN
                           => n5285);
   U5924 : NAND4_X1 port map( A1 => n5288, A2 => n5287, A3 => n5286, A4 => 
                           n5285, ZN => n5301);
   U5925 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_21xx31x, A2 => n5290,
                           B1 => fromRegsPortxREG_FILE_22xx31x, B2 => n5289, ZN
                           => n5299);
   U5926 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_20xx31x, A2 => n5292,
                           B1 => fromRegsPortxREG_FILE_23xx31x, B2 => n5291, ZN
                           => n5298);
   U5927 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_17xx31x, A2 => n5294,
                           B1 => fromRegsPortxREG_FILE_19xx31x, B2 => n5293, ZN
                           => n5297);
   U5928 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_18xx31x, A2 => n5295,
                           ZN => n5296);
   U5929 : NAND4_X1 port map( A1 => n5299, A2 => n5298, A3 => n5297, A4 => 
                           n5296, ZN => n5300);
   U5930 : AOI21_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(23), B2 => n5301
                           , A => n5300, ZN => n5315);
   U5931 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_12xx31x, A2 => n5303,
                           B1 => fromRegsPortxREG_FILE_10xx31x, B2 => n5302, ZN
                           => n5313);
   U5932 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_11xx31x, A2 => n5305,
                           B1 => fromRegsPortxREG_FILE_14xx31x, B2 => n5304, ZN
                           => n5309);
   U5933 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_15xx31x, A2 => n5307,
                           B1 => fromRegsPortxREG_FILE_13xx31x, B2 => n5306, ZN
                           => n5308);
   U5934 : NAND2_X1 port map( A1 => n5309, A2 => n5308, ZN => n5310);
   U5935 : AOI21_X1 port map( B1 => n5311, B2 => fromRegsPortxREG_FILE_16xx31x,
                           A => n5310, ZN => n5312);
   U5936 : OAI211_X1 port map( C1 => n5315, C2 => n5314, A => n5313, B => n5312
                           , ZN => n5317);
   U5937 : NAND2_X1 port map( A1 => n5317, A2 => n5316, ZN => n5337);
   U5938 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_06xx31x, A2 => n5319,
                           B1 => fromRegsPortxREG_FILE_03xx31x, B2 => n5318, ZN
                           => n5328);
   U5939 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_09xx31x, A2 => n5321,
                           B1 => fromRegsPortxREG_FILE_04xx31x, B2 => n5320, ZN
                           => n5327);
   U5940 : AOI22_X1 port map( A1 => fromRegsPortxREG_FILE_05xx31x, A2 => n5323,
                           B1 => fromRegsPortxREG_FILE_07xx31x, B2 => n5322, ZN
                           => n5326);
   U5941 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_08xx31x, A2 => n5324,
                           ZN => n5325);
   U5942 : NAND4_X1 port map( A1 => n5328, A2 => n5327, A3 => n5326, A4 => 
                           n5325, ZN => n5335);
   U5943 : NAND2_X1 port map( A1 => n5329, A2 => fromRegsPortxREG_FILE_02xx31x,
                           ZN => n5332);
   U5944 : NAND2_X1 port map( A1 => fromRegsPortxREG_FILE_01xx31x, A2 => n5330,
                           ZN => n5331);
   U5945 : NAND2_X1 port map( A1 => n5332, A2 => n5331, ZN => n5333);
   U5946 : AOI21_X1 port map( B1 => n5335, B2 => n5334, A => n5333, ZN => n5336
                           );
   U5947 : NAND2_X1 port map( A1 => n5337, A2 => n5336, ZN => n7388);
   U5948 : XOR2_X1 port map( A => n7551, B => n7388, Z => n5389);
   U5949 : AOI22_X1 port map( A1 => n5339, A2 => fromRegsPortxREG_FILE_30xx31x,
                           B1 => n5338, B2 => fromRegsPortxREG_FILE_23xx31x, ZN
                           => n5349);
   U5950 : AOI22_X1 port map( A1 => n5341, A2 => fromRegsPortxREG_FILE_11xx31x,
                           B1 => n5340, B2 => fromRegsPortxREG_FILE_09xx31x, ZN
                           => n5348);
   U5951 : AOI22_X1 port map( A1 => n5343, A2 => fromRegsPortxREG_FILE_07xx31x,
                           B1 => n5342, B2 => fromRegsPortxREG_FILE_21xx31x, ZN
                           => n5347);
   U5952 : AOI22_X1 port map( A1 => n5345, A2 => fromRegsPortxREG_FILE_16xx31x,
                           B1 => n5344, B2 => fromRegsPortxREG_FILE_15xx31x, ZN
                           => n5346);
   U5953 : AND4_X1 port map( A1 => n5349, A2 => n5348, A3 => n5347, A4 => n5346
                           , ZN => n5388);
   U5954 : AOI22_X1 port map( A1 => n5351, A2 => fromRegsPortxREG_FILE_29xx31x,
                           B1 => n5350, B2 => fromRegsPortxREG_FILE_17xx31x, ZN
                           => n5361);
   U5955 : AOI22_X1 port map( A1 => n5353, A2 => fromRegsPortxREG_FILE_27xx31x,
                           B1 => n5352, B2 => fromRegsPortxREG_FILE_22xx31x, ZN
                           => n5360);
   U5956 : AOI22_X1 port map( A1 => n5355, A2 => fromRegsPortxREG_FILE_03xx31x,
                           B1 => n5354, B2 => fromRegsPortxREG_FILE_20xx31x, ZN
                           => n5359);
   U5957 : AOI22_X1 port map( A1 => n5357, A2 => fromRegsPortxREG_FILE_04xx31x,
                           B1 => n5356, B2 => fromRegsPortxREG_FILE_12xx31x, ZN
                           => n5358);
   U5958 : AND4_X1 port map( A1 => n5361, A2 => n5360, A3 => n5359, A4 => n5358
                           , ZN => n5387);
   U5959 : AOI22_X1 port map( A1 => n5363, A2 => fromRegsPortxREG_FILE_25xx31x,
                           B1 => n5362, B2 => fromRegsPortxREG_FILE_06xx31x, ZN
                           => n5373);
   U5960 : AOI22_X1 port map( A1 => n5365, A2 => fromRegsPortxREG_FILE_26xx31x,
                           B1 => n5364, B2 => fromRegsPortxREG_FILE_18xx31x, ZN
                           => n5372);
   U5961 : AOI22_X1 port map( A1 => n5367, A2 => fromRegsPortxREG_FILE_19xx31x,
                           B1 => n5366, B2 => fromRegsPortxREG_FILE_13xx31x, ZN
                           => n5371);
   U5962 : AOI22_X1 port map( A1 => n5369, A2 => fromRegsPortxREG_FILE_10xx31x,
                           B1 => n5368, B2 => fromRegsPortxREG_FILE_14xx31x, ZN
                           => n5370);
   U5963 : AND4_X1 port map( A1 => n5373, A2 => n5372, A3 => n5371, A4 => n5370
                           , ZN => n5386);
   U5964 : AOI22_X1 port map( A1 => n5375, A2 => fromRegsPortxREG_FILE_02xx31x,
                           B1 => n5374, B2 => fromRegsPortxREG_FILE_05xx31x, ZN
                           => n5384);
   U5965 : AOI22_X1 port map( A1 => n5377, A2 => fromRegsPortxREG_FILE_28xx31x,
                           B1 => n5376, B2 => fromRegsPortxREG_FILE_24xx31x, ZN
                           => n5383);
   U5966 : NAND2_X1 port map( A1 => n5378, A2 => fromRegsPortxREG_FILE_08xx31x,
                           ZN => n5382);
   U5967 : AOI22_X1 port map( A1 => n5380, A2 => fromRegsPortxREG_FILE_01xx31x,
                           B1 => n5379, B2 => fromRegsPortxREG_FILE_31xx31x, ZN
                           => n5381);
   U5968 : AND4_X1 port map( A1 => n5384, A2 => n5383, A3 => n5382, A4 => n5381
                           , ZN => n5385);
   U5969 : NAND4_X1 port map( A1 => n5388, A2 => n5387, A3 => n5386, A4 => 
                           n5385, ZN => n7413);
   U5970 : XOR2_X1 port map( A => n5389, B => n7413, Z => n5390);
   U5971 : XOR2_X1 port map( A => DP_OP_679J14_122_3096xn2, B => n5390, Z => 
                           n5395);
   U5972 : OR4_X1 port map( A1 => DP_OP_679J14_122_3096xn88, A2 => 
                           DP_OP_679J14_122_3096xn87, A3 => 
                           DP_OP_679J14_122_3096xn71, A4 => 
                           DP_OP_679J14_122_3096xn69, ZN => n5391);
   U5973 : OR4_X1 port map( A1 => DP_OP_679J14_122_3096xn91, A2 => 
                           DP_OP_679J14_122_3096xn90, A3 => 
                           DP_OP_679J14_122_3096xn89, A4 => n5391, ZN => n5392)
                           ;
   U5974 : OR4_X1 port map( A1 => DP_OP_679J14_122_3096xn94, A2 => 
                           DP_OP_679J14_122_3096xn93, A3 => 
                           DP_OP_679J14_122_3096xn92, A4 => n5392, ZN => n5393)
                           ;
   U5975 : OR4_X1 port map( A1 => DP_OP_679J14_122_3096xn97, A2 => 
                           DP_OP_679J14_122_3096xn96, A3 => 
                           DP_OP_679J14_122_3096xn95, A4 => n5393, ZN => n5394)
                           ;
   U5976 : OR4_X1 port map( A1 => n5395, A2 => DP_OP_679J14_122_3096xn99, A3 =>
                           DP_OP_679J14_122_3096xn98, A4 => n5394, ZN => n5401)
                           ;
   U5977 : OR4_X1 port map( A1 => DP_OP_679J14_122_3096xn74, A2 => 
                           DP_OP_679J14_122_3096xn73, A3 => 
                           DP_OP_679J14_122_3096xn72, A4 => 
                           DP_OP_679J14_122_3096xn70, ZN => n5396);
   U5978 : OR4_X1 port map( A1 => DP_OP_679J14_122_3096xn77, A2 => 
                           DP_OP_679J14_122_3096xn76, A3 => 
                           DP_OP_679J14_122_3096xn75, A4 => n5396, ZN => n5397)
                           ;
   U5979 : OR4_X1 port map( A1 => DP_OP_679J14_122_3096xn80, A2 => 
                           DP_OP_679J14_122_3096xn79, A3 => 
                           DP_OP_679J14_122_3096xn78, A4 => n5397, ZN => n5398)
                           ;
   U5980 : OR4_X1 port map( A1 => DP_OP_679J14_122_3096xn83, A2 => 
                           DP_OP_679J14_122_3096xn82, A3 => 
                           DP_OP_679J14_122_3096xn81, A4 => n5398, ZN => n5399)
                           ;
   U5981 : OR4_X1 port map( A1 => DP_OP_679J14_122_3096xn86, A2 => 
                           DP_OP_679J14_122_3096xn85, A3 => 
                           DP_OP_679J14_122_3096xn84, A4 => n5399, ZN => n5400)
                           ;
   U5982 : NOR2_X1 port map( A1 => n5401, A2 => n5400, ZN => n5629);
   U5983 : INV_X1 port map( A => n7413, ZN => n7435);
   U5984 : NOR2_X1 port map( A1 => n7487, A2 => ashr_25xAx30x, ZN => n7328);
   U5985 : NOR2_X1 port map( A1 => n7481, A2 => ashr_25xAx25x, ZN => n7074);
   U5986 : OAI22_X1 port map( A1 => n7477, A2 => ashr_25xAx21x, B1 => n7476, B2
                           => ashr_25xAx20x, ZN => n5425);
   U5987 : AOI22_X1 port map( A1 => n7476, A2 => ashr_25xAx20x, B1 => n7475, B2
                           => ashr_25xAx19x, ZN => n5424);
   U5988 : INV_X1 port map( A => ashr_25xAx15x, ZN => n6766);
   U5989 : AOI22_X1 port map( A1 => n6766, A2 => n6739, B1 => intadd_27xAx3x, 
                           B2 => n6693, ZN => n5417);
   U5990 : NAND2_X1 port map( A1 => n7466, A2 => ashr_25xAx10x, ZN => n6501);
   U5991 : INV_X1 port map( A => ashr_25xAx9x, ZN => n6481);
   U5992 : NOR2_X1 port map( A1 => n6481, A2 => n6480, ZN => n6478);
   U5993 : NOR2_X1 port map( A1 => n7464, A2 => ashr_25xAx8x, ZN => n6444);
   U5994 : INV_X1 port map( A => ashr_25xAx7x, ZN => n6399);
   U5995 : INV_X1 port map( A => ashr_25xAx6x, ZN => n6330);
   U5996 : AOI22_X1 port map( A1 => n6399, A2 => n6377, B1 => n6330, B2 => 
                           n6326, ZN => n5409);
   U5997 : INV_X1 port map( A => ashr_25xAx5x, ZN => n6048);
   U5998 : NAND2_X1 port map( A1 => n6048, A2 => n5402, ZN => n6302);
   U5999 : NAND2_X1 port map( A1 => n7192, A2 => ashr_25xAx4x, ZN => n6239);
   U6000 : CLKBUF_X1 port map( A => n7402, Z => n5711);
   U6001 : NOR2_X1 port map( A1 => intadd_29xAx0x, A2 => n5711, ZN => n6067);
   U6002 : NOR2_X1 port map( A1 => n7268, A2 => ashr_25xAx0x, ZN => n5685);
   U6003 : NOR2_X1 port map( A1 => n7304, A2 => ashr_25xAx1x, ZN => n6064);
   U6004 : OAI22_X1 port map( A1 => n5685, A2 => n6064, B1 => intadd_29xAx1x, 
                           B2 => n7309, ZN => n5403);
   U6005 : NAND2_X1 port map( A1 => intadd_29xAx1x, A2 => n7309, ZN => n6106);
   U6006 : NAND2_X1 port map( A1 => intadd_29xAx2x, A2 => n7207, ZN => n6161);
   U6007 : OAI211_X1 port map( C1 => n6067, C2 => n5403, A => n6106, B => n6161
                           , ZN => n5404);
   U6008 : OAI211_X1 port map( C1 => intadd_29xAx2x, C2 => n7207, A => n6239, B
                           => n5404, ZN => n5405);
   U6009 : OAI211_X1 port map( C1 => n7192, C2 => ashr_25xAx4x, A => n6302, B 
                           => n5405, ZN => n5406);
   U6010 : NAND2_X1 port map( A1 => n7461, A2 => ashr_25xAx5x, ZN => n6291);
   U6011 : OAI211_X1 port map( C1 => n6330, C2 => n6326, A => n5406, B => n6291
                           , ZN => n5408);
   U6012 : INV_X1 port map( A => ashr_25xAx8x, ZN => n6419);
   U6013 : NOR2_X1 port map( A1 => n6419, A2 => n6421, ZN => n6445);
   U6014 : NOR2_X1 port map( A1 => n6399, A2 => n6377, ZN => n5407);
   U6015 : AOI211_X1 port map( C1 => n5409, C2 => n5408, A => n6445, B => n5407
                           , ZN => n5410);
   U6016 : AOI211_X1 port map( C1 => n6481, C2 => n6480, A => n6444, B => n5410
                           , ZN => n5411);
   U6017 : OAI22_X1 port map( A1 => n6478, A2 => n5411, B1 => n7466, B2 => 
                           ashr_25xAx10x, ZN => n5412);
   U6018 : AOI22_X1 port map( A1 => intadd_27xAx0x, A2 => n6553, B1 => n6501, 
                           B2 => n5412, ZN => n5414);
   U6019 : OAI22_X1 port map( A1 => intadd_27xAx0x, A2 => n6553, B1 => 
                           intadd_27xAx1x, B2 => n6626, ZN => n5413);
   U6020 : NAND2_X1 port map( A1 => intadd_27xAx1x, A2 => n6626, ZN => n6613);
   U6021 : NAND2_X1 port map( A1 => intadd_27xAx2x, A2 => n6669, ZN => n6657);
   U6022 : OAI211_X1 port map( C1 => n5414, C2 => n5413, A => n6613, B => n6657
                           , ZN => n5415);
   U6023 : NAND2_X1 port map( A1 => n7469, A2 => ashr_25xAx13x, ZN => n6656);
   U6024 : OAI211_X1 port map( C1 => intadd_27xAx3x, C2 => n6693, A => n5415, B
                           => n6656, ZN => n5416);
   U6025 : AOI22_X1 port map( A1 => n7471, A2 => ashr_25xAx15x, B1 => n5417, B2
                           => n5416, ZN => n5418);
   U6026 : NAND2_X1 port map( A1 => n7472, A2 => ashr_25xAx16x, ZN => n6778);
   U6027 : NOR2_X1 port map( A1 => n7473, A2 => ashr_25xAx17x, ZN => n6802);
   U6028 : NOR2_X1 port map( A1 => n7472, A2 => ashr_25xAx16x, ZN => n6779);
   U6029 : AOI211_X1 port map( C1 => n5418, C2 => n6778, A => n6802, B => n6779
                           , ZN => n5420);
   U6030 : OAI22_X1 port map( A1 => intadd_26xAx0x, A2 => n6806, B1 => 
                           intadd_26xAx1x, B2 => n6861, ZN => n5419);
   U6031 : NAND2_X1 port map( A1 => intadd_26xAx1x, A2 => n6861, ZN => n6855);
   U6032 : NAND2_X1 port map( A1 => intadd_26xAx2x, A2 => n6888, ZN => n6887);
   U6033 : OAI211_X1 port map( C1 => n5420, C2 => n5419, A => n6855, B => n6887
                           , ZN => n5423);
   U6034 : OAI22_X1 port map( A1 => intadd_26xAx4x, A2 => n5720, B1 => 
                           intadd_26xAx5x, B2 => n6958, ZN => n5421);
   U6035 : AOI21_X1 port map( B1 => n7479, B2 => ashr_25xAx23x, A => n5421, ZN 
                           => n5422);
   U6036 : OAI221_X1 port map( B1 => n5425, B2 => n5424, C1 => n5425, C2 => 
                           n5423, A => n5422, ZN => n5427);
   U6037 : NOR2_X1 port map( A1 => n7479, A2 => ashr_25xAx23x, ZN => n6997);
   U6038 : NOR2_X1 port map( A1 => n7478, A2 => ashr_25xAx22x, ZN => n6974);
   U6039 : OAI22_X1 port map( A1 => intadd_26xAx6x, A2 => n7009, B1 => n6997, 
                           B2 => n6974, ZN => n5426);
   U6040 : AOI22_X1 port map( A1 => n7480, A2 => ashr_25xAx24x, B1 => n5427, B2
                           => n5426, ZN => n5428);
   U6041 : AOI211_X1 port map( C1 => intadd_26xAx7x, C2 => n7053, A => n7074, B
                           => n5428, ZN => n5433);
   U6042 : INV_X1 port map( A => ashr_25xAx27x, ZN => n7184);
   U6043 : INV_X1 port map( A => ashr_25xAx26x, ZN => n7160);
   U6044 : AOI22_X1 port map( A1 => n7184, A2 => n7183, B1 => n7160, B2 => 
                           n7120, ZN => n5432);
   U6045 : INV_X1 port map( A => ashr_25xAx25x, ZN => n7129);
   U6046 : OAI22_X1 port map( A1 => n7160, A2 => n7120, B1 => n7129, B2 => 
                           n7097, ZN => n5431);
   U6047 : NAND2_X1 port map( A1 => n7485, A2 => ashr_25xAx29x, ZN => n5429);
   U6048 : NAND2_X1 port map( A1 => n7483, A2 => ashr_25xAx27x, ZN => n7181);
   U6049 : OAI211_X1 port map( C1 => intadd_28xAx0x, C2 => n7242, A => n5429, B
                           => n7181, ZN => n5430);
   U6050 : AOI221_X1 port map( B1 => n5433, B2 => n5432, C1 => n5431, C2 => 
                           n5432, A => n5430, ZN => n5434);
   U6051 : AOI211_X1 port map( C1 => intadd_28xAx1x, C2 => n7252, A => n7328, B
                           => n5434, ZN => n5436);
   U6052 : OAI211_X1 port map( C1 => intadd_28xAx1x, C2 => n7252, A => 
                           intadd_28xAx0x, B => n7242, ZN => n5435);
   U6053 : AOI22_X1 port map( A1 => n7487, A2 => ashr_25xAx30x, B1 => n5436, B2
                           => n5435, ZN => n5439);
   U6054 : INV_X1 port map( A => n7388, ZN => n7489);
   U6055 : NAND2_X1 port map( A1 => n7489, A2 => n7413, ZN => n5437);
   U6056 : AOI22_X1 port map( A1 => n7435, A2 => n7388, B1 => n5439, B2 => 
                           n5437, ZN => n5634);
   U6057 : NAND2_X1 port map( A1 => n7435, A2 => n7388, ZN => n5438);
   U6058 : AOI22_X1 port map( A1 => n5439, A2 => n5438, B1 => n7489, B2 => 
                           n7413, ZN => n5633);
   U6059 : AOI221_X1 port map( B1 => fromMemoryPortxLOADEDDATAx(13), B2 => 
                           n5634, C1 => n6670, C2 => n5633, A => n6716, ZN => 
                           n5440);
   U6060 : AOI21_X1 port map( B1 => n5955, B2 => n5629, A => n5440, ZN => n5441
                           );
   U6061 : CLKBUF_X1 port map( A => n5658, Z => n5620);
   U6062 : INV_X2 port map( A => n5620, ZN => n5746);
   U6063 : NAND2_X1 port map( A1 => IF_ISAxpcReg_signal_2_port, A2 => 
                           IF_ISAxpcReg_signal_3_port, ZN => n5616);
   U6064 : INV_X1 port map( A => n5616, ZN => n5612);
   U6065 : NAND2_X1 port map( A1 => n5612, A2 => IF_ISAxpcReg_signal_4_port, ZN
                           => n5611);
   U6066 : INV_X1 port map( A => n5611, ZN => n5605);
   U6067 : NAND2_X1 port map( A1 => n5605, A2 => IF_ISAxpcReg_signal_5_port, ZN
                           => n5604);
   U6068 : NOR2_X1 port map( A1 => n5604, A2 => n7543, ZN => n5599);
   U6069 : NAND2_X1 port map( A1 => n5599, A2 => IF_ISAxpcReg_signal_7_port, ZN
                           => n5592);
   U6070 : NOR2_X1 port map( A1 => n5592, A2 => n7544, ZN => n5585);
   U6071 : NAND2_X1 port map( A1 => n5585, A2 => IF_ISAxpcReg_signal_9_port, ZN
                           => n5578);
   U6072 : NOR2_X1 port map( A1 => n5578, A2 => n7545, ZN => n5571);
   U6073 : NAND2_X1 port map( A1 => n5571, A2 => IF_ISAxpcReg_signal_11_port, 
                           ZN => n5564);
   U6074 : INV_X1 port map( A => n5564, ZN => n5442);
   U6075 : AND2_X1 port map( A1 => n5442, A2 => IF_ISAxpcReg_signal_12_port, ZN
                           => n5559);
   U6076 : NAND2_X1 port map( A1 => n5559, A2 => IF_ISAxpcReg_signal_13_port, 
                           ZN => n5554);
   U6077 : INV_X1 port map( A => n5554, ZN => n5548);
   U6078 : NAND2_X1 port map( A1 => n5548, A2 => IF_ISAxpcReg_signal_14_port, 
                           ZN => n5547);
   U6079 : INV_X1 port map( A => n5547, ZN => n5542);
   U6080 : NAND2_X1 port map( A1 => n5542, A2 => IF_ISAxpcReg_signal_15_port, 
                           ZN => n5541);
   U6081 : INV_X1 port map( A => n5541, ZN => n5537);
   U6082 : NAND2_X1 port map( A1 => n5537, A2 => IF_ISAxpcReg_signal_16_port, 
                           ZN => n5536);
   U6083 : INV_X1 port map( A => n5536, ZN => n5530);
   U6084 : NAND2_X1 port map( A1 => n5530, A2 => IF_ISAxpcReg_signal_17_port, 
                           ZN => n5529);
   U6085 : INV_X1 port map( A => n5529, ZN => n5523);
   U6086 : NAND2_X1 port map( A1 => n5523, A2 => IF_ISAxpcReg_signal_18_port, 
                           ZN => n5522);
   U6087 : INV_X1 port map( A => n5522, ZN => n5516);
   U6088 : NAND2_X1 port map( A1 => n5516, A2 => IF_ISAxpcReg_signal_19_port, 
                           ZN => n5515);
   U6089 : INV_X1 port map( A => n5515, ZN => n5510);
   U6090 : NAND2_X1 port map( A1 => n5510, A2 => IF_ISAxpcReg_signal_20_port, 
                           ZN => n5509);
   U6091 : INV_X1 port map( A => n5509, ZN => n5503);
   U6092 : NAND2_X1 port map( A1 => n5503, A2 => IF_ISAxpcReg_signal_21_port, 
                           ZN => n5502);
   U6093 : INV_X1 port map( A => n5502, ZN => n5496);
   U6094 : NAND2_X1 port map( A1 => n5496, A2 => IF_ISAxpcReg_signal_22_port, 
                           ZN => n5495);
   U6095 : INV_X1 port map( A => n5495, ZN => n5490);
   U6096 : NAND2_X1 port map( A1 => n5490, A2 => IF_ISAxpcReg_signal_23_port, 
                           ZN => n5489);
   U6097 : INV_X1 port map( A => n5489, ZN => n5484);
   U6098 : NAND2_X1 port map( A1 => n5484, A2 => IF_ISAxpcReg_signal_24_port, 
                           ZN => n5483);
   U6099 : INV_X1 port map( A => n5483, ZN => n5476);
   U6100 : NAND2_X1 port map( A1 => n5476, A2 => IF_ISAxpcReg_signal_25_port, 
                           ZN => n5475);
   U6101 : INV_X1 port map( A => n5475, ZN => n5468);
   U6102 : NAND2_X1 port map( A1 => n5468, A2 => IF_ISAxpcReg_signal_26_port, 
                           ZN => n5467);
   U6103 : INV_X1 port map( A => n5467, ZN => n5462);
   U6104 : NAND2_X1 port map( A1 => n5462, A2 => IF_ISAxpcReg_signal_27_port, 
                           ZN => n5461);
   U6105 : INV_X1 port map( A => n5461, ZN => n5456);
   U6106 : NAND2_X1 port map( A1 => n5456, A2 => IF_ISAxpcReg_signal_28_port, 
                           ZN => n5455);
   U6107 : INV_X1 port map( A => n5455, ZN => n5450);
   U6108 : NAND2_X1 port map( A1 => n5450, A2 => IF_ISAxpcReg_signal_29_port, 
                           ZN => n5449);
   U6109 : INV_X1 port map( A => n5449, ZN => n5655);
   U6110 : XOR2_X1 port map( A => n5655, B => IF_ISAxpcReg_signal_30_port, Z =>
                           n7361);
   U6111 : AOI22_X1 port map( A1 => n5746, A2 => n7361, B1 => intadd_25xSUMx28x
                           , B2 => n5620, ZN => n5928);
   U6112 : NOR2_X1 port map( A1 => IF_ISAxsection_2_port, A2 => n7538, ZN => 
                           n7458);
   U6113 : NAND2_X1 port map( A1 => IF_ISAxsection_2_port, A2 => n7538, ZN => 
                           n5961);
   U6114 : INV_X1 port map( A => n5961, ZN => n5646);
   U6115 : NOR2_X1 port map( A1 => n7458, A2 => n5646, ZN => n7453);
   U6116 : OR2_X1 port map( A1 => n5740, A2 => fromMemoryPortxLOADEDDATAx(6), 
                           ZN => n5747);
   U6117 : AOI21_X1 port map( B1 => n7453, B2 => n5747, A => rst, ZN => n5608);
   U6118 : CLKBUF_X1 port map( A => n5608, Z => n5660);
   U6119 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(12), A2 => n5443
                           , ZN => n5666);
   U6120 : INV_X1 port map( A => n5666, ZN => n5627);
   U6121 : NAND2_X1 port map( A1 => n5746, A2 => n5444, ZN => n5743);
   U6122 : CLKBUF_X1 port map( A => n5743, Z => n5586);
   U6123 : INV_X1 port map( A => n5586, ZN => n5657);
   U6124 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx28x, B1 => n7361
                           , B2 => n5586, ZN => n5931);
   U6125 : INV_X1 port map( A => n5931, ZN => n5445);
   U6126 : AOI22_X1 port map( A1 => n7361, A2 => n5660, B1 => n5627, B2 => 
                           n5445, ZN => n5448);
   U6127 : NAND2_X1 port map( A1 => n5827, A2 => n7535, ZN => n5958);
   U6128 : NOR3_X1 port map( A1 => n5748, A2 => n5739, A3 => n5958, ZN => n5568
                           );
   U6129 : CLKBUF_X1 port map( A => n5568, Z => n5663);
   U6130 : NOR3_X1 port map( A1 => n5936, A2 => n5748, A3 => n5740, ZN => n5662
                           );
   U6131 : INV_X1 port map( A => intadd_28xSUMx2x, ZN => n5446);
   U6132 : AOI22_X1 port map( A1 => intadd_25xSUMx28x, A2 => n5663, B1 => n5662
                           , B2 => n5446, ZN => n5447);
   U6133 : OAI211_X1 port map( C1 => n5625, C2 => n5928, A => n5448, B => n5447
                           , ZN => n7558);
   U6134 : OAI21_X1 port map( B1 => n5450, B2 => IF_ISAxpcReg_signal_29_port, A
                           => n5449, ZN => n5927);
   U6135 : INV_X1 port map( A => n5927, ZN => n7296);
   U6136 : AOI22_X1 port map( A1 => n5746, A2 => n7296, B1 => intadd_25xSUMx27x
                           , B2 => n5658, ZN => n5923);
   U6137 : INV_X1 port map( A => n5586, ZN => n5744);
   U6138 : AOI22_X1 port map( A1 => n5744, A2 => intadd_25xSUMx27x, B1 => n7296
                           , B2 => n5586, ZN => n5926);
   U6139 : INV_X1 port map( A => n5926, ZN => n5451);
   U6140 : AOI22_X1 port map( A1 => n7296, A2 => n5660, B1 => n5627, B2 => 
                           n5451, ZN => n5454);
   U6141 : INV_X1 port map( A => n5662, ZN => n5580);
   U6142 : INV_X1 port map( A => n5580, ZN => n5622);
   U6143 : INV_X1 port map( A => intadd_28xSUMx1x, ZN => n5452);
   U6144 : AOI22_X1 port map( A1 => intadd_25xSUMx27x, A2 => n5663, B1 => n5622
                           , B2 => n5452, ZN => n5453);
   U6145 : OAI211_X1 port map( C1 => n5625, C2 => n5923, A => n5454, B => n5453
                           , ZN => n7559);
   U6146 : OAI21_X1 port map( B1 => n5456, B2 => IF_ISAxpcReg_signal_28_port, A
                           => n5455, ZN => n5922);
   U6147 : INV_X1 port map( A => n5922, ZN => n7248);
   U6148 : AOI22_X1 port map( A1 => n5746, A2 => n7248, B1 => intadd_25xSUMx26x
                           , B2 => n5658, ZN => n5917);
   U6149 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx26x, B1 => n7248
                           , B2 => n5743, ZN => n5918);
   U6150 : INV_X1 port map( A => n5918, ZN => n5457);
   U6151 : AOI22_X1 port map( A1 => n7248, A2 => n5660, B1 => n5627, B2 => 
                           n5457, ZN => n5460);
   U6152 : INV_X1 port map( A => intadd_28xSUMx0x, ZN => n5458);
   U6153 : AOI22_X1 port map( A1 => intadd_25xSUMx26x, A2 => n5663, B1 => n5662
                           , B2 => n5458, ZN => n5459);
   U6154 : OAI211_X1 port map( C1 => n5625, C2 => n5917, A => n5460, B => n5459
                           , ZN => n7560);
   U6155 : OAI21_X1 port map( B1 => n5462, B2 => IF_ISAxpcReg_signal_27_port, A
                           => n5461, ZN => n5915);
   U6156 : INV_X1 port map( A => n5915, ZN => n7204);
   U6157 : AOI22_X1 port map( A1 => n5744, A2 => intadd_25xSUMx25x, B1 => n7204
                           , B2 => n5586, ZN => n5914);
   U6158 : INV_X1 port map( A => intadd_25xSUMx25x, ZN => n7185);
   U6159 : AOI22_X1 port map( A1 => n5746, A2 => n5915, B1 => n7185, B2 => 
                           n5658, ZN => n5910);
   U6160 : AOI22_X1 port map( A1 => n7204, A2 => n5660, B1 => n5910, B2 => 
                           n5659, ZN => n5466);
   U6161 : NOR2_X1 port map( A1 => n7129, A2 => add_x_26xBx25x, ZN => n6002);
   U6162 : AOI21_X1 port map( B1 => n7129, B2 => add_x_26xBx25x, A => n6002, ZN
                           => n5479);
   U6163 : NOR2_X1 port map( A1 => n5479, A2 => intadd_26xn1, ZN => n5463);
   U6164 : AOI21_X1 port map( B1 => ashr_25xAx25x, B2 => add_x_26xBx25x, A => 
                           n5463, ZN => n5471);
   U6165 : INV_X1 port map( A => n5464, ZN => n5916);
   U6166 : OAI22_X1 port map( A1 => ashr_25xAx27x, A2 => add_x_26xBx27x, B1 => 
                           n7168, B2 => n7184, ZN => n7182);
   U6167 : XNOR2_X1 port map( A => n5916, B => n7182, ZN => n5912);
   U6168 : AOI22_X1 port map( A1 => intadd_25xSUMx25x, A2 => n5663, B1 => n5622
                           , B2 => n5912, ZN => n5465);
   U6169 : OAI211_X1 port map( C1 => n5914, C2 => n5666, A => n5466, B => n5465
                           , ZN => n7561);
   U6170 : OAI21_X1 port map( B1 => n5468, B2 => IF_ISAxpcReg_signal_26_port, A
                           => n5467, ZN => n7117);
   U6171 : INV_X1 port map( A => n7117, ZN => n5470);
   U6172 : AOI22_X1 port map( A1 => n5746, A2 => n5470, B1 => intadd_25xSUMx24x
                           , B2 => n5658, ZN => n5904);
   U6173 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx24x, B1 => n5470
                           , B2 => n5586, ZN => n5905);
   U6174 : INV_X1 port map( A => n5905, ZN => n5469);
   U6175 : AOI22_X1 port map( A1 => n5470, A2 => n5660, B1 => n5627, B2 => 
                           n5469, ZN => n5474);
   U6176 : FA_X1 port map( A => n7160, B => n7126, CI => n5471, CO => n5464, S 
                           => n5906);
   U6177 : INV_X1 port map( A => n5906, ZN => n5472);
   U6178 : AOI22_X1 port map( A1 => intadd_25xSUMx24x, A2 => n5663, B1 => n5662
                           , B2 => n5472, ZN => n5473);
   U6179 : OAI211_X1 port map( C1 => n5625, C2 => n5904, A => n5474, B => n5473
                           , ZN => n7562);
   U6180 : OAI21_X1 port map( B1 => n5476, B2 => IF_ISAxpcReg_signal_25_port, A
                           => n5475, ZN => n7079);
   U6181 : INV_X1 port map( A => n7079, ZN => n5478);
   U6182 : AOI22_X1 port map( A1 => n5746, A2 => n5478, B1 => intadd_25xSUMx23x
                           , B2 => n5620, ZN => n5898);
   U6183 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx23x, B1 => n5478
                           , B2 => n5743, ZN => n5899);
   U6184 : INV_X1 port map( A => n5899, ZN => n5477);
   U6185 : AOI22_X1 port map( A1 => n5478, A2 => n5660, B1 => n5627, B2 => 
                           n5477, ZN => n5482);
   U6186 : XNOR2_X1 port map( A => n5479, B => intadd_26xn1, ZN => n5900);
   U6187 : INV_X1 port map( A => n5900, ZN => n5480);
   U6188 : AOI22_X1 port map( A1 => intadd_25xSUMx23x, A2 => n5663, B1 => n5480
                           , B2 => n5662, ZN => n5481);
   U6189 : OAI211_X1 port map( C1 => n5625, C2 => n5898, A => n5482, B => n5481
                           , ZN => n7563);
   U6190 : OAI21_X1 port map( B1 => n5484, B2 => IF_ISAxpcReg_signal_24_port, A
                           => n5483, ZN => n5897);
   U6191 : INV_X1 port map( A => n5897, ZN => n7054);
   U6192 : AOI22_X1 port map( A1 => n5746, A2 => n7054, B1 => intadd_25xSUMx22x
                           , B2 => n5658, ZN => n5892);
   U6193 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx22x, B1 => n7054
                           , B2 => n5743, ZN => n5893);
   U6194 : INV_X1 port map( A => n5893, ZN => n5485);
   U6195 : AOI22_X1 port map( A1 => n7054, A2 => n5660, B1 => n5627, B2 => 
                           n5485, ZN => n5488);
   U6196 : INV_X1 port map( A => intadd_26xSUMx7x, ZN => n5486);
   U6197 : AOI22_X1 port map( A1 => intadd_25xSUMx22x, A2 => n5663, B1 => n5622
                           , B2 => n5486, ZN => n5487);
   U6198 : OAI211_X1 port map( C1 => n5625, C2 => n5892, A => n5488, B => n5487
                           , ZN => n7564);
   U6199 : OAI21_X1 port map( B1 => n5490, B2 => IF_ISAxpcReg_signal_23_port, A
                           => n5489, ZN => n5891);
   U6200 : INV_X1 port map( A => n5891, ZN => n6996);
   U6201 : AOI22_X1 port map( A1 => n5746, A2 => n6996, B1 => intadd_25xSUMx21x
                           , B2 => n5658, ZN => n5887);
   U6202 : AOI22_X1 port map( A1 => n5744, A2 => intadd_25xSUMx21x, B1 => n6996
                           , B2 => n5743, ZN => n5890);
   U6203 : INV_X1 port map( A => n5890, ZN => n5491);
   U6204 : AOI22_X1 port map( A1 => n6996, A2 => n5660, B1 => n5627, B2 => 
                           n5491, ZN => n5494);
   U6205 : INV_X1 port map( A => intadd_26xSUMx6x, ZN => n5492);
   U6206 : AOI22_X1 port map( A1 => intadd_25xSUMx21x, A2 => n5663, B1 => n5622
                           , B2 => n5492, ZN => n5493);
   U6207 : OAI211_X1 port map( C1 => n5625, C2 => n5887, A => n5494, B => n5493
                           , ZN => n7565);
   U6208 : OAI21_X1 port map( B1 => n5496, B2 => IF_ISAxpcReg_signal_22_port, A
                           => n5495, ZN => n6983);
   U6209 : INV_X1 port map( A => n6983, ZN => n5498);
   U6210 : AOI22_X1 port map( A1 => n5746, A2 => n5498, B1 => intadd_25xSUMx20x
                           , B2 => n5658, ZN => n5882);
   U6211 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx20x, B1 => n5498
                           , B2 => n5743, ZN => n5883);
   U6212 : INV_X1 port map( A => n5883, ZN => n5497);
   U6213 : AOI22_X1 port map( A1 => n5498, A2 => n5660, B1 => n5627, B2 => 
                           n5497, ZN => n5501);
   U6214 : INV_X1 port map( A => intadd_26xSUMx5x, ZN => n5499);
   U6215 : AOI22_X1 port map( A1 => intadd_25xSUMx20x, A2 => n5663, B1 => n5622
                           , B2 => n5499, ZN => n5500);
   U6216 : OAI211_X1 port map( C1 => n5625, C2 => n5882, A => n5501, B => n5500
                           , ZN => n7566);
   U6217 : OAI21_X1 port map( B1 => n5503, B2 => IF_ISAxpcReg_signal_21_port, A
                           => n5502, ZN => n5881);
   U6218 : INV_X1 port map( A => n5881, ZN => n5505);
   U6219 : AOI22_X1 port map( A1 => n5746, A2 => n5505, B1 => intadd_25xSUMx19x
                           , B2 => n5658, ZN => n5876);
   U6220 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx19x, B1 => n5505
                           , B2 => n5743, ZN => n5877);
   U6221 : INV_X1 port map( A => n5877, ZN => n5504);
   U6222 : AOI22_X1 port map( A1 => n5505, A2 => n5660, B1 => n5627, B2 => 
                           n5504, ZN => n5508);
   U6223 : INV_X1 port map( A => intadd_26xSUMx4x, ZN => n5506);
   U6224 : AOI22_X1 port map( A1 => intadd_25xSUMx19x, A2 => n5663, B1 => n5622
                           , B2 => n5506, ZN => n5507);
   U6225 : OAI211_X1 port map( C1 => n5625, C2 => n5876, A => n5508, B => n5507
                           , ZN => n7567);
   U6226 : OAI21_X1 port map( B1 => n5510, B2 => IF_ISAxpcReg_signal_20_port, A
                           => n5509, ZN => n5875);
   U6227 : INV_X1 port map( A => n5875, ZN => n6926);
   U6228 : AOI22_X1 port map( A1 => n5746, A2 => n6926, B1 => intadd_25xSUMx18x
                           , B2 => n5658, ZN => n5870);
   U6229 : AOI22_X1 port map( A1 => n5744, A2 => intadd_25xSUMx18x, B1 => n6926
                           , B2 => n5743, ZN => n5871);
   U6230 : INV_X1 port map( A => n5871, ZN => n5511);
   U6231 : AOI22_X1 port map( A1 => n6926, A2 => n5660, B1 => n5627, B2 => 
                           n5511, ZN => n5514);
   U6232 : INV_X1 port map( A => intadd_26xSUMx3x, ZN => n5512);
   U6233 : AOI22_X1 port map( A1 => intadd_25xSUMx18x, A2 => n5663, B1 => n5622
                           , B2 => n5512, ZN => n5513);
   U6234 : OAI211_X1 port map( C1 => n5625, C2 => n5870, A => n5514, B => n5513
                           , ZN => n7568);
   U6235 : OAI21_X1 port map( B1 => n5516, B2 => IF_ISAxpcReg_signal_19_port, A
                           => n5515, ZN => n6893);
   U6236 : INV_X1 port map( A => n6893, ZN => n5518);
   U6237 : AOI22_X1 port map( A1 => n5746, A2 => n5518, B1 => intadd_25xSUMx17x
                           , B2 => n5658, ZN => n5864);
   U6238 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx17x, B1 => n5518
                           , B2 => n5743, ZN => n5866);
   U6239 : INV_X1 port map( A => n5866, ZN => n5517);
   U6240 : AOI22_X1 port map( A1 => n5518, A2 => n5660, B1 => n5627, B2 => 
                           n5517, ZN => n5521);
   U6241 : INV_X1 port map( A => intadd_26xSUMx2x, ZN => n5519);
   U6242 : AOI22_X1 port map( A1 => intadd_25xSUMx17x, A2 => n5568, B1 => n5622
                           , B2 => n5519, ZN => n5520);
   U6243 : OAI211_X1 port map( C1 => n5625, C2 => n5864, A => n5521, B => n5520
                           , ZN => n7569);
   U6244 : OAI21_X1 port map( B1 => n5523, B2 => IF_ISAxpcReg_signal_18_port, A
                           => n5522, ZN => n6859);
   U6245 : INV_X1 port map( A => n6859, ZN => n5525);
   U6246 : AOI22_X1 port map( A1 => n5746, A2 => n5525, B1 => intadd_25xSUMx16x
                           , B2 => n5658, ZN => n5860);
   U6247 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx16x, B1 => n5525
                           , B2 => n5743, ZN => n5863);
   U6248 : INV_X1 port map( A => n5863, ZN => n5524);
   U6249 : AOI22_X1 port map( A1 => n5525, A2 => n5660, B1 => n5627, B2 => 
                           n5524, ZN => n5528);
   U6250 : INV_X1 port map( A => intadd_26xSUMx1x, ZN => n5526);
   U6251 : AOI22_X1 port map( A1 => intadd_25xSUMx16x, A2 => n5568, B1 => n5622
                           , B2 => n5526, ZN => n5527);
   U6252 : OAI211_X1 port map( C1 => n5625, C2 => n5860, A => n5528, B => n5527
                           , ZN => n7570);
   U6253 : OAI21_X1 port map( B1 => n5530, B2 => IF_ISAxpcReg_signal_17_port, A
                           => n5529, ZN => n6805);
   U6254 : INV_X1 port map( A => n6805, ZN => n5532);
   U6255 : AOI22_X1 port map( A1 => n5746, A2 => n5532, B1 => intadd_25xSUMx15x
                           , B2 => n5658, ZN => n5856);
   U6256 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx15x, B1 => n5532
                           , B2 => n5743, ZN => n5859);
   U6257 : INV_X1 port map( A => n5859, ZN => n5531);
   U6258 : AOI22_X1 port map( A1 => n5532, A2 => n5660, B1 => n5627, B2 => 
                           n5531, ZN => n5535);
   U6259 : INV_X1 port map( A => intadd_26xSUMx0x, ZN => n5533);
   U6260 : AOI22_X1 port map( A1 => intadd_25xSUMx15x, A2 => n5663, B1 => n5622
                           , B2 => n5533, ZN => n5534);
   U6261 : OAI211_X1 port map( C1 => n5625, C2 => n5856, A => n5535, B => n5534
                           , ZN => n7571);
   U6262 : OAI21_X1 port map( B1 => n5537, B2 => IF_ISAxpcReg_signal_16_port, A
                           => n5536, ZN => n5854);
   U6263 : INV_X1 port map( A => n5854, ZN => n6776);
   U6264 : AOI22_X1 port map( A1 => n5746, A2 => n6776, B1 => intadd_25xSUMx14x
                           , B2 => n5658, ZN => n5849);
   U6265 : INV_X1 port map( A => ashr_25xAx16x, ZN => n6774);
   U6266 : AOI22_X1 port map( A1 => n6774, A2 => n6783, B1 => add_x_26xBx16x, 
                           B2 => ashr_25xAx16x, ZN => n6775);
   U6267 : AOI22_X1 port map( A1 => n6766, A2 => add_x_26xBx15x, B1 => n6743, 
                           B2 => ashr_25xAx15x, ZN => n6744);
   U6268 : OAI22_X1 port map( A1 => n6766, A2 => n6743, B1 => n6744, B2 => 
                           intadd_27xn1, ZN => n5855);
   U6269 : XOR2_X1 port map( A => n6775, B => n5855, Z => n5848);
   U6270 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx14x, B1 => n6776
                           , B2 => n5743, ZN => n5850);
   U6271 : INV_X1 port map( A => n5850, ZN => n5538);
   U6272 : AOI22_X1 port map( A1 => n5848, A2 => n5622, B1 => n5627, B2 => 
                           n5538, ZN => n5540);
   U6273 : AOI22_X1 port map( A1 => n6776, A2 => n5660, B1 => intadd_25xSUMx14x
                           , B2 => n5663, ZN => n5539);
   U6274 : OAI211_X1 port map( C1 => n5625, C2 => n5849, A => n5540, B => n5539
                           , ZN => n7572);
   U6275 : OAI21_X1 port map( B1 => n5542, B2 => IF_ISAxpcReg_signal_15_port, A
                           => n5541, ZN => n6742);
   U6276 : INV_X1 port map( A => n6742, ZN => n5544);
   U6277 : AOI22_X1 port map( A1 => n5746, A2 => n5544, B1 => intadd_25xSUMx13x
                           , B2 => n5658, ZN => n5843);
   U6278 : XOR2_X1 port map( A => n6744, B => intadd_27xn1, Z => n5842);
   U6279 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx13x, B1 => n5544
                           , B2 => n5743, ZN => n5844);
   U6280 : INV_X1 port map( A => n5844, ZN => n5543);
   U6281 : AOI22_X1 port map( A1 => n5842, A2 => n5622, B1 => n5627, B2 => 
                           n5543, ZN => n5546);
   U6282 : AOI22_X1 port map( A1 => n5544, A2 => n5608, B1 => intadd_25xSUMx13x
                           , B2 => n5663, ZN => n5545);
   U6283 : OAI211_X1 port map( C1 => n5625, C2 => n5843, A => n5546, B => n5545
                           , ZN => n7573);
   U6284 : OAI21_X1 port map( B1 => n5548, B2 => IF_ISAxpcReg_signal_14_port, A
                           => n5547, ZN => n6687);
   U6285 : INV_X1 port map( A => n6687, ZN => n5550);
   U6286 : AOI22_X1 port map( A1 => n5746, A2 => n5550, B1 => intadd_25xSUMx12x
                           , B2 => n5658, ZN => n5838);
   U6287 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx12x, B1 => n5550
                           , B2 => n5586, ZN => n5841);
   U6288 : INV_X1 port map( A => n5841, ZN => n5549);
   U6289 : AOI22_X1 port map( A1 => n5550, A2 => n5608, B1 => n5627, B2 => 
                           n5549, ZN => n5553);
   U6290 : INV_X1 port map( A => intadd_27xSUMx3x, ZN => n5551);
   U6291 : AOI22_X1 port map( A1 => intadd_25xSUMx12x, A2 => n5568, B1 => n5622
                           , B2 => n5551, ZN => n5552);
   U6292 : OAI211_X1 port map( C1 => n5625, C2 => n5838, A => n5553, B => n5552
                           , ZN => n7574);
   U6293 : OAI21_X1 port map( B1 => n5559, B2 => IF_ISAxpcReg_signal_13_port, A
                           => n5554, ZN => n5837);
   U6294 : INV_X1 port map( A => n5837, ZN => n6635);
   U6295 : AOI22_X1 port map( A1 => n5746, A2 => n6635, B1 => intadd_25xSUMx11x
                           , B2 => n5620, ZN => n5832);
   U6296 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx11x, B1 => n6635
                           , B2 => n5586, ZN => n5833);
   U6297 : INV_X1 port map( A => n5833, ZN => n5555);
   U6298 : AOI22_X1 port map( A1 => n6635, A2 => n5608, B1 => n5627, B2 => 
                           n5555, ZN => n5558);
   U6299 : INV_X1 port map( A => intadd_27xSUMx2x, ZN => n5556);
   U6300 : AOI22_X1 port map( A1 => intadd_25xSUMx11x, A2 => n5568, B1 => n5622
                           , B2 => n5556, ZN => n5557);
   U6301 : OAI211_X1 port map( C1 => n5625, C2 => n5832, A => n5558, B => n5557
                           , ZN => n7575);
   U6302 : AOI21_X1 port map( B1 => n5564, B2 => n7547, A => n5559, ZN => n6612
                           );
   U6303 : AOI22_X1 port map( A1 => n5746, A2 => n6612, B1 => intadd_25xSUMx10x
                           , B2 => n5658, ZN => n5825);
   U6304 : INV_X1 port map( A => intadd_25xSUMx10x, ZN => n6611);
   U6305 : INV_X1 port map( A => n6612, ZN => n5560);
   U6306 : AOI22_X1 port map( A1 => n5657, A2 => n6611, B1 => n5560, B2 => 
                           n5743, ZN => n5823);
   U6307 : AOI22_X1 port map( A1 => n6612, A2 => n5608, B1 => n5627, B2 => 
                           n5823, ZN => n5563);
   U6308 : INV_X1 port map( A => intadd_27xSUMx1x, ZN => n5561);
   U6309 : AOI22_X1 port map( A1 => intadd_25xSUMx10x, A2 => n5568, B1 => n5622
                           , B2 => n5561, ZN => n5562);
   U6310 : OAI211_X1 port map( C1 => n5625, C2 => n5825, A => n5563, B => n5562
                           , ZN => n7576);
   U6311 : OAI21_X1 port map( B1 => n5571, B2 => IF_ISAxpcReg_signal_11_port, A
                           => n5564, ZN => n6572);
   U6312 : INV_X1 port map( A => n6572, ZN => n5566);
   U6313 : AOI22_X1 port map( A1 => n5746, A2 => n5566, B1 => intadd_25xSUMx9x,
                           B2 => n5658, ZN => n5817);
   U6314 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx9x, B1 => n5566,
                           B2 => n5743, ZN => n5818);
   U6315 : INV_X1 port map( A => n5818, ZN => n5565);
   U6316 : AOI22_X1 port map( A1 => n5566, A2 => n5608, B1 => n5627, B2 => 
                           n5565, ZN => n5570);
   U6317 : INV_X1 port map( A => intadd_27xSUMx0x, ZN => n5567);
   U6318 : AOI22_X1 port map( A1 => intadd_25xSUMx9x, A2 => n5568, B1 => n5622,
                           B2 => n5567, ZN => n5569);
   U6319 : OAI211_X1 port map( C1 => n5625, C2 => n5817, A => n5570, B => n5569
                           , ZN => n7577);
   U6320 : AOI21_X1 port map( B1 => n5578, B2 => n7545, A => n5571, ZN => n6507
                           );
   U6321 : AOI22_X1 port map( A1 => n5746, A2 => n6507, B1 => intadd_25xSUMx8x,
                           B2 => n5658, ZN => n5809);
   U6322 : OAI22_X1 port map( A1 => ashr_25xAx9x, A2 => n6476, B1 => 
                           add_x_26xBx9x, B2 => n6481, ZN => n6479);
   U6323 : NOR2_X1 port map( A1 => n6419, A2 => n5587, ZN => n6439);
   U6324 : NOR2_X1 port map( A1 => ashr_25xAx4x, A2 => ashr_25xSHx4x, ZN => 
                           n5572);
   U6325 : NAND2_X1 port map( A1 => ashr_25xAx4x, A2 => ashr_25xSHx4x, ZN => 
                           n6241);
   U6326 : OAI21_X1 port map( B1 => n5572, B2 => intadd_29xn1, A => n6241, ZN 
                           => n5606);
   U6327 : INV_X1 port map( A => n5606, ZN => n5573);
   U6328 : AOI22_X1 port map( A1 => n6048, A2 => add_x_26xBx5x, B1 => n6283, B2
                           => ashr_25xAx5x, ZN => n5607);
   U6329 : INV_X1 port map( A => n5607, ZN => n6272);
   U6330 : AOI22_X1 port map( A1 => n6048, A2 => n6283, B1 => n5573, B2 => 
                           n6272, ZN => n5601);
   U6331 : OAI22_X1 port map( A1 => add_x_26xBx8x, A2 => ashr_25xAx8x, B1 => 
                           n6439, B2 => n5588, ZN => n5579);
   U6332 : AOI22_X1 port map( A1 => n6481, A2 => n6476, B1 => n6479, B2 => 
                           n5579, ZN => n5816);
   U6333 : INV_X1 port map( A => ashr_25xAx10x, ZN => n6528);
   U6334 : NOR2_X1 port map( A1 => n5814, A2 => n6528, ZN => n6540);
   U6335 : AOI21_X1 port map( B1 => n5814, B2 => n6528, A => n6540, ZN => n5574
                           );
   U6336 : INV_X1 port map( A => n5574, ZN => n6512);
   U6337 : XOR2_X1 port map( A => n5816, B => n6512, Z => n5808);
   U6338 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx8x, B1 => n6507,
                           B2 => n5743, ZN => n5813);
   U6339 : OAI22_X1 port map( A1 => n5808, A2 => n5580, B1 => n5666, B2 => 
                           n5813, ZN => n5575);
   U6340 : INV_X1 port map( A => n5575, ZN => n5577);
   U6341 : AOI22_X1 port map( A1 => intadd_25xSUMx8x, A2 => n5663, B1 => n6507,
                           B2 => n5660, ZN => n5576);
   U6342 : OAI211_X1 port map( C1 => n5625, C2 => n5809, A => n5577, B => n5576
                           , ZN => n7578);
   U6343 : OAI21_X1 port map( B1 => n5585, B2 => IF_ISAxpcReg_signal_9_port, A 
                           => n5578, ZN => n6472);
   U6344 : INV_X1 port map( A => n6472, ZN => n5582);
   U6345 : AOI22_X1 port map( A1 => n5746, A2 => n5582, B1 => intadd_25xSUMx7x,
                           B2 => n5658, ZN => n5802);
   U6346 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx7x, B1 => n5582,
                           B2 => n5743, ZN => n5801);
   U6347 : XOR2_X1 port map( A => n6479, B => n5579, Z => n5803);
   U6348 : OAI22_X1 port map( A1 => n5666, A2 => n5801, B1 => n5580, B2 => 
                           n5803, ZN => n5581);
   U6349 : INV_X1 port map( A => n5581, ZN => n5584);
   U6350 : AOI22_X1 port map( A1 => n5582, A2 => n5608, B1 => intadd_25xSUMx7x,
                           B2 => n5663, ZN => n5583);
   U6351 : OAI211_X1 port map( C1 => n5625, C2 => n5802, A => n5584, B => n5583
                           , ZN => n7579);
   U6352 : AOI21_X1 port map( B1 => n5592, B2 => n7544, A => n5585, ZN => n6438
                           );
   U6353 : AOI22_X1 port map( A1 => n5746, A2 => n6438, B1 => intadd_25xSUMx6x,
                           B2 => n5658, ZN => n5795);
   U6354 : AOI22_X1 port map( A1 => n5657, A2 => intadd_25xSUMx6x, B1 => n6438,
                           B2 => n5586, ZN => n5800);
   U6355 : INV_X1 port map( A => n5800, ZN => n5589);
   U6356 : AOI22_X1 port map( A1 => n6419, A2 => add_x_26xBx8x, B1 => n5587, B2
                           => ashr_25xAx8x, ZN => n6448);
   U6357 : XNOR2_X1 port map( A => n5588, B => n6448, ZN => n5794);
   U6358 : AOI22_X1 port map( A1 => n5627, A2 => n5589, B1 => n5622, B2 => 
                           n5794, ZN => n5591);
   U6359 : AOI22_X1 port map( A1 => intadd_25xSUMx6x, A2 => n5663, B1 => n6438,
                           B2 => n5660, ZN => n5590);
   U6360 : OAI211_X1 port map( C1 => n5625, C2 => n5795, A => n5591, B => n5590
                           , ZN => n7580);
   U6361 : OR2_X1 port map( A1 => n5599, A2 => IF_ISAxpcReg_signal_7_port, ZN 
                           => n5593);
   U6362 : AND2_X1 port map( A1 => n5593, A2 => n5592, ZN => n5595);
   U6363 : AOI22_X1 port map( A1 => n5744, A2 => intadd_25xSUMx5x, B1 => n5595,
                           B2 => n5743, ZN => n5790);
   U6364 : INV_X1 port map( A => n5595, ZN => n6393);
   U6365 : INV_X1 port map( A => intadd_25xSUMx5x, ZN => n5594);
   U6366 : AOI22_X1 port map( A1 => n5746, A2 => n6393, B1 => n5594, B2 => 
                           n5658, ZN => n5788);
   U6367 : AOI22_X1 port map( A1 => n5595, A2 => n5608, B1 => n5788, B2 => 
                           n5659, ZN => n5598);
   U6368 : FA_X1 port map( A => ashr_25xAx7x, B => add_x_26xBx7x, CI => n5596, 
                           CO => n5588, S => n5792);
   U6369 : AOI22_X1 port map( A1 => n5792, A2 => n5622, B1 => intadd_25xSUMx5x,
                           B2 => n5663, ZN => n5597);
   U6370 : OAI211_X1 port map( C1 => n5790, C2 => n5666, A => n5598, B => n5597
                           , ZN => n7581);
   U6371 : AOI21_X1 port map( B1 => n5604, B2 => n7543, A => n5599, ZN => n6335
                           );
   U6372 : AOI22_X1 port map( A1 => n5746, A2 => n6335, B1 => intadd_25xSUMx4x,
                           B2 => n5658, ZN => n5781);
   U6373 : AOI22_X1 port map( A1 => n5744, A2 => intadd_25xSUMx4x, B1 => n6335,
                           B2 => n5743, ZN => n5786);
   U6374 : INV_X1 port map( A => n5786, ZN => n5600);
   U6375 : AOI22_X1 port map( A1 => n6335, A2 => n5608, B1 => n5627, B2 => 
                           n5600, ZN => n5603);
   U6376 : FA_X1 port map( A => ashr_25xAx6x, B => add_x_26xBx6x, CI => n5601, 
                           CO => n5596, S => n5782);
   U6377 : AOI22_X1 port map( A1 => intadd_25xSUMx4x, A2 => n5663, B1 => n5782,
                           B2 => n5622, ZN => n5602);
   U6378 : OAI211_X1 port map( C1 => n5625, C2 => n5781, A => n5603, B => n5602
                           , ZN => n7582);
   U6379 : OAI21_X1 port map( B1 => n5605, B2 => IF_ISAxpcReg_signal_5_port, A 
                           => n5604, ZN => n5780);
   U6380 : INV_X1 port map( A => n5780, ZN => n6282);
   U6381 : AOI22_X1 port map( A1 => n5744, A2 => intadd_25xSUMx3x, B1 => n6282,
                           B2 => n5743, ZN => n5779);
   U6382 : INV_X1 port map( A => intadd_25xSUMx3x, ZN => n6290);
   U6383 : AOI22_X1 port map( A1 => n5746, A2 => n5780, B1 => n6290, B2 => 
                           n5658, ZN => n5776);
   U6384 : XNOR2_X1 port map( A => n5607, B => n5606, ZN => n5777);
   U6385 : AOI22_X1 port map( A1 => n5776, A2 => n5659, B1 => n5622, B2 => 
                           n5777, ZN => n5610);
   U6386 : AOI22_X1 port map( A1 => n6282, A2 => n5608, B1 => intadd_25xSUMx3x,
                           B2 => n5663, ZN => n5609);
   U6387 : OAI211_X1 port map( C1 => n5779, C2 => n5666, A => n5610, B => n5609
                           , ZN => n7583);
   U6388 : OAI21_X1 port map( B1 => n5612, B2 => IF_ISAxpcReg_signal_4_port, A 
                           => n5611, ZN => n6240);
   U6389 : INV_X1 port map( A => n6240, ZN => n5769);
   U6390 : AOI22_X1 port map( A1 => n5746, A2 => n5769, B1 => intadd_25xSUMx2x,
                           B2 => n5658, ZN => n5771);
   U6391 : INV_X1 port map( A => intadd_25xSUMx2x, ZN => n6260);
   U6392 : AOI22_X1 port map( A1 => n5744, A2 => n6260, B1 => n6240, B2 => 
                           n5743, ZN => n5770);
   U6393 : OAI21_X1 port map( B1 => ashr_25xSHx4x, B2 => ashr_25xAx4x, A => 
                           n6241, ZN => n6259);
   U6394 : XNOR2_X1 port map( A => intadd_29xn1, B => n6259, ZN => n5775);
   U6395 : INV_X1 port map( A => n5775, ZN => n5613);
   U6396 : AOI22_X1 port map( A1 => n5627, A2 => n5770, B1 => n5622, B2 => 
                           n5613, ZN => n5615);
   U6397 : AOI22_X1 port map( A1 => intadd_25xSUMx2x, A2 => n5663, B1 => n5769,
                           B2 => n5660, ZN => n5614);
   U6398 : OAI211_X1 port map( C1 => n5625, C2 => n5771, A => n5615, B => n5614
                           , ZN => n7584);
   U6399 : OAI21_X1 port map( B1 => IF_ISAxpcReg_signal_2_port, B2 => 
                           IF_ISAxpcReg_signal_3_port, A => n5616, ZN => n6189)
                           ;
   U6400 : INV_X1 port map( A => n6189, ZN => n5763);
   U6401 : AOI22_X1 port map( A1 => n5746, A2 => n5763, B1 => intadd_25xSUMx1x,
                           B2 => n5620, ZN => n5765);
   U6402 : INV_X1 port map( A => intadd_25xSUMx1x, ZN => n6215);
   U6403 : AOI22_X1 port map( A1 => n5744, A2 => n6215, B1 => n6189, B2 => 
                           n5743, ZN => n5764);
   U6404 : AOI22_X1 port map( A1 => n5763, A2 => n5660, B1 => n5764, B2 => 
                           n5627, ZN => n5619);
   U6405 : INV_X1 port map( A => intadd_29xSUMx2x, ZN => n5617);
   U6406 : AOI22_X1 port map( A1 => intadd_25xSUMx1x, A2 => n5663, B1 => n5662,
                           B2 => n5617, ZN => n5618);
   U6407 : OAI211_X1 port map( C1 => n5625, C2 => n5765, A => n5619, B => n5618
                           , ZN => n7585);
   U6408 : INV_X1 port map( A => intadd_25xSUMx0x, ZN => n6094);
   U6409 : AOI22_X1 port map( A1 => n5744, A2 => n6094, B1 => 
                           IF_ISAxpcReg_signal_2_port, B2 => n5743, ZN => n5758
                           );
   U6410 : AOI22_X1 port map( A1 => n5746, A2 => n7546, B1 => n5620, B2 => 
                           intadd_25xSUMx0x, ZN => n5759);
   U6411 : INV_X1 port map( A => intadd_29xSUMx1x, ZN => n5621);
   U6412 : AOI22_X1 port map( A1 => intadd_25xSUMx0x, A2 => n5663, B1 => n5622,
                           B2 => n5621, ZN => n5624);
   U6413 : NAND2_X1 port map( A1 => n5660, A2 => n7546, ZN => n5623);
   U6414 : OAI211_X1 port map( C1 => n5759, C2 => n5625, A => n5624, B => n5623
                           , ZN => n5626);
   U6415 : AOI21_X1 port map( B1 => n5758, B2 => n5627, A => n5626, ZN => n5628
                           );
   U6416 : INV_X1 port map( A => n5628, ZN => n7586);
   U6417 : NOR2_X1 port map( A1 => intadd_29xBx0x, A2 => n7542, ZN => 
                           intadd_25xCI);
   U6418 : INV_X1 port map( A => n5629, ZN => n5635);
   U6419 : INV_X1 port map( A => n5630, ZN => n5631);
   U6420 : INV_X1 port map( A => n5692, ZN => n5727);
   U6421 : NAND3_X1 port map( A1 => n5632, A2 => n5631, A3 => n5727, ZN => 
                           n6017);
   U6422 : OR2_X1 port map( A1 => n5719, A2 => n5692, ZN => n6015);
   U6423 : OAI22_X1 port map( A1 => n5634, A2 => n6017, B1 => n5633, B2 => 
                           n6015, ZN => n6019);
   U6424 : AOI21_X1 port map( B1 => n5635, B2 => n5680, A => n6019, ZN => n5640
                           );
   U6425 : NAND3_X1 port map( A1 => n5640, A2 => n5637, A3 => n5636, ZN => 
                           n5638);
   U6426 : OAI21_X1 port map( B1 => n5640, B2 => n5639, A => n5638, ZN => n5648
                           );
   U6427 : INV_X1 port map( A => n5648, ZN => n5641);
   U6428 : AOI22_X1 port map( A1 => n7458, A2 => IF_ISAxsection_0_port, B1 => 
                           n5642, B2 => n5641, ZN => n5668);
   U6429 : INV_X1 port map( A => n5668, ZN => n5644);
   U6430 : INV_X2 port map( A => n7416, ZN => n7418);
   U6431 : AOI21_X1 port map( B1 => n7418, B2 => n7542, A => intadd_25xCI, ZN 
                           => n6068);
   U6432 : INV_X1 port map( A => n6068, ZN => n5643);
   U6433 : AOI21_X1 port map( B1 => n7458, B2 => IF_ISAxsection_0_port, A => 
                           n7118, ZN => n5647);
   U6434 : NAND3_X1 port map( A1 => n5642, A2 => n7457, A3 => n5647, ZN => 
                           n5669);
   U6435 : OAI22_X1 port map( A1 => n5644, A2 => n5643, B1 => n5669, B2 => 
                           intadd_29xSUMx0x, ZN => n5645);
   U6436 : AND2_X1 port map( A1 => IF_ISAxsection_0_port, A2 => 
                           fromMemoryPort_sync_port, ZN => n7455);
   U6437 : NAND2_X1 port map( A1 => n5646, A2 => n7455, ZN => n7526);
   U6438 : NAND2_X1 port map( A1 => n5645, A2 => n7526, ZN => n5650);
   U6439 : NAND2_X1 port map( A1 => IF_ISAxsection_0_port, A2 => n5646, ZN => 
                           n6044);
   U6440 : NOR2_X1 port map( A1 => rst, A2 => n6044, ZN => n6597);
   U6441 : NAND2_X1 port map( A1 => fromMemoryPort_sync_port, A2 => n6597, ZN 
                           => n7531);
   U6442 : OAI211_X1 port map( C1 => n5648, C2 => n7457, A => n5647, B => n7531
                           , ZN => n5667);
   U6443 : NAND2_X1 port map( A1 => n5667, A2 => IF_ISAxN2460, ZN => n5649);
   U6444 : AOI21_X1 port map( B1 => n5650, B2 => n5649, A => rst, ZN => 
                           IF_ISAxN10904);
   U6445 : NAND2_X1 port map( A1 => n5651, A2 => fromMemoryPortxLOADEDDATAx(31)
                           , ZN => n5652);
   U6446 : NAND2_X1 port map( A1 => n5653, A2 => n5652, ZN => n7379);
   U6447 : INV_X1 port map( A => n7379, ZN => n7392);
   U6448 : AOI22_X1 port map( A1 => n7379, A2 => n7548, B1 => 
                           IF_ISAxpcReg_signal_31_port, B2 => n7392, ZN => 
                           n5654);
   U6449 : XNOR2_X1 port map( A => intadd_25xn1, B => n5654, ZN => n5942);
   U6450 : NAND2_X1 port map( A1 => n5655, A2 => IF_ISAxpcReg_signal_30_port, 
                           ZN => n5656);
   U6451 : XOR2_X1 port map( A => IF_ISAxpcReg_signal_31_port, B => n5656, Z =>
                           n5946);
   U6452 : INV_X1 port map( A => n5946, ZN => n7438);
   U6453 : AOI22_X1 port map( A1 => n5657, A2 => n5942, B1 => n7438, B2 => 
                           n5743, ZN => n5945);
   U6454 : INV_X1 port map( A => n5942, ZN => n7383);
   U6455 : AOI22_X1 port map( A1 => n5746, A2 => n5946, B1 => n7383, B2 => 
                           n5658, ZN => n5940);
   U6456 : AOI22_X1 port map( A1 => n7438, A2 => n5660, B1 => n5940, B2 => 
                           n5659, ZN => n5665);
   U6457 : NAND2_X1 port map( A1 => n7435, A2 => n7379, ZN => n6013);
   U6458 : OAI21_X1 port map( B1 => n7435, B2 => n7379, A => n6013, ZN => n5661
                           );
   U6459 : XNOR2_X1 port map( A => n5661, B => intadd_28xn1, ZN => n5949);
   U6460 : AOI22_X1 port map( A1 => n5942, A2 => n5663, B1 => n5949, B2 => 
                           n5662, ZN => n5664);
   U6461 : OAI211_X1 port map( C1 => n5945, C2 => n5666, A => n5665, B => n5664
                           , ZN => n7557);
   U6462 : OAI21_X1 port map( B1 => n5668, B2 => n5667, A => IF_ISAxN2459, ZN 
                           => n5673);
   U6463 : NAND2_X1 port map( A1 => n7414, A2 => ashr_25xAx0x, ZN => n6250);
   U6464 : INV_X2 port map( A => n7130, ZN => n7414);
   U6465 : NOR2_X1 port map( A1 => ashr_25xAx0x, A2 => n7414, ZN => n5972);
   U6466 : INV_X1 port map( A => n5972, ZN => n5966);
   U6467 : AOI21_X1 port map( B1 => n6250, B2 => n5966, A => n5669, ZN => n5670
                           );
   U6468 : INV_X1 port map( A => n5670, ZN => n5672);
   U6469 : NOR2_X1 port map( A1 => n7526, A2 => IF_ISAxN2459, ZN => n5671);
   U6470 : AOI211_X1 port map( C1 => n5673, C2 => n5672, A => rst, B => n5671, 
                           ZN => n7552);
   U6471 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => intadd_28xAx2x, ZN
                           => DP_OP_719J14_125_1055xn164);
   U6472 : AOI21_X1 port map( B1 => n5674, B2 => n7364, A => intadd_28xAx1x, ZN
                           => DP_OP_719J14_125_1055xn163);
   U6473 : AOI21_X1 port map( B1 => n5675, B2 => n5678, A => intadd_28xAx0x, ZN
                           => DP_OP_719J14_125_1055xn162);
   U6474 : AOI21_X1 port map( B1 => n5675, B2 => n7364, A => n7184, ZN => 
                           DP_OP_719J14_125_1055xn161);
   U6475 : AOI21_X1 port map( B1 => n5675, B2 => n7364, A => n7160, ZN => 
                           DP_OP_719J14_125_1055xn160);
   U6476 : AOI21_X1 port map( B1 => n5675, B2 => n5678, A => n7129, ZN => 
                           DP_OP_719J14_125_1055xn159);
   U6477 : AOI21_X1 port map( B1 => n5675, B2 => n7364, A => intadd_26xAx7x, ZN
                           => DP_OP_719J14_125_1055xn158);
   U6478 : AOI21_X1 port map( B1 => n5675, B2 => n7364, A => intadd_26xAx6x, ZN
                           => DP_OP_719J14_125_1055xn157);
   U6479 : AOI21_X1 port map( B1 => n5675, B2 => n5678, A => intadd_26xAx5x, ZN
                           => DP_OP_719J14_125_1055xn156);
   U6480 : AOI21_X1 port map( B1 => n5675, B2 => n7364, A => intadd_26xAx4x, ZN
                           => DP_OP_719J14_125_1055xn155);
   U6481 : AOI21_X1 port map( B1 => n5675, B2 => n5677, A => intadd_26xAx3x, ZN
                           => DP_OP_719J14_125_1055xn154);
   U6482 : AOI21_X1 port map( B1 => n5679, B2 => n5677, A => intadd_26xAx2x, ZN
                           => DP_OP_719J14_125_1055xn153);
   U6483 : AOI21_X1 port map( B1 => n5675, B2 => n5677, A => intadd_26xAx1x, ZN
                           => DP_OP_719J14_125_1055xn152);
   U6484 : AOI21_X1 port map( B1 => n5679, B2 => n5677, A => intadd_26xAx0x, ZN
                           => DP_OP_719J14_125_1055xn151);
   U6485 : AOI21_X1 port map( B1 => n5675, B2 => n5677, A => n6774, ZN => 
                           DP_OP_719J14_125_1055xn150);
   U6486 : AOI21_X1 port map( B1 => n5675, B2 => n5676, A => n6766, ZN => 
                           DP_OP_719J14_125_1055xn149);
   U6487 : AOI21_X1 port map( B1 => n5679, B2 => n5677, A => intadd_27xAx3x, ZN
                           => DP_OP_719J14_125_1055xn148);
   U6488 : AOI21_X1 port map( B1 => n5679, B2 => n5676, A => intadd_27xAx2x, ZN
                           => DP_OP_719J14_125_1055xn147);
   U6489 : AOI21_X1 port map( B1 => n5679, B2 => n5677, A => intadd_27xAx1x, ZN
                           => DP_OP_719J14_125_1055xn146);
   U6490 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => intadd_27xAx0x, ZN
                           => DP_OP_719J14_125_1055xn145);
   U6491 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => n6528, ZN => 
                           DP_OP_719J14_125_1055xn144);
   U6492 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => n6481, ZN => 
                           DP_OP_719J14_125_1055xn143);
   U6493 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => n6419, ZN => 
                           DP_OP_719J14_125_1055xn142);
   U6494 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => n6399, ZN => 
                           DP_OP_719J14_125_1055xn141);
   U6495 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => n6330, ZN => 
                           DP_OP_719J14_125_1055xn140);
   U6496 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => n6048, ZN => 
                           DP_OP_719J14_125_1055xn139);
   U6497 : INV_X1 port map( A => ashr_25xAx4x, ZN => n6251);
   U6498 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => n6251, ZN => 
                           DP_OP_719J14_125_1055xn138);
   U6499 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => intadd_29xAx2x, ZN
                           => DP_OP_719J14_125_1055xn137);
   U6500 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => intadd_29xAx1x, ZN
                           => DP_OP_719J14_125_1055xn136);
   U6501 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => intadd_29xAx0x, ZN
                           => DP_OP_719J14_125_1055xn135);
   U6502 : INV_X1 port map( A => ashr_25xAx0x, ZN => n6026);
   U6503 : AOI21_X1 port map( B1 => n5679, B2 => n5678, A => n6026, ZN => 
                           DP_OP_719J14_125_1055xn134);
   U6504 : NOR2_X1 port map( A1 => n5680, A2 => n5693, ZN => n5682);
   U6505 : NOR2_X1 port map( A1 => n5682, A2 => n5681, ZN => n7159);
   U6506 : INV_X2 port map( A => n7399, ZN => n7209);
   U6507 : AOI22_X1 port map( A1 => n7209, A2 => intadd_26xAx4x, B1 => 
                           intadd_26xAx5x, B2 => n7086, ZN => n6196);
   U6508 : OAI22_X1 port map( A1 => n7086, A2 => intadd_26xAx6x, B1 => 
                           intadd_26xAx7x, B2 => n7209, ZN => n6199);
   U6509 : AOI22_X1 port map( A1 => n7304, A2 => n6196, B1 => n6199, B2 => 
                           n7402, ZN => n6066);
   U6510 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx27x, B1 => 
                           ashr_25xAx28x, B2 => n7399, ZN => n6195);
   U6511 : OAI22_X1 port map( A1 => n7267, A2 => n7129, B1 => n7160, B2 => 
                           n7209, ZN => n6198);
   U6512 : INV_X1 port map( A => n6198, ZN => n5683);
   U6513 : MUX2_X1 port map( A => n6195, B => n5683, S => n7304, Z => n6065);
   U6514 : AOI22_X1 port map( A1 => n6941, A2 => n6066, B1 => n6065, B2 => 
                           n6900, ZN => n6642);
   U6515 : NOR2_X1 port map( A1 => n7376, A2 => n6900, ZN => n6365);
   U6516 : INV_X2 port map( A => n7402, ZN => n7404);
   U6517 : NAND2_X1 port map( A1 => n7209, A2 => n7413, ZN => n6219);
   U6518 : OAI22_X1 port map( A1 => n7267, A2 => ashr_25xAx29x, B1 => 
                           ashr_25xAx30x, B2 => n7209, ZN => n6194);
   U6519 : OR2_X1 port map( A1 => n5711, A2 => n6194, ZN => n5712);
   U6520 : OAI21_X1 port map( B1 => n7404, B2 => n6219, A => n5712, ZN => n6645
                           );
   U6521 : AOI22_X1 port map( A1 => n7376, A2 => n6642, B1 => n6365, B2 => 
                           n6645, ZN => n6309);
   U6522 : NAND2_X1 port map( A1 => n5690, A2 => n6020, ZN => n5684);
   U6523 : NOR2_X1 port map( A1 => n5689, A2 => n5684, ZN => n6346);
   U6524 : AND2_X1 port map( A1 => n6346, A2 => n7192, ZN => n7046);
   U6525 : INV_X1 port map( A => n7046, ZN => n7427);
   U6526 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx5x, B1 => 
                           ashr_25xAx4x, B2 => n7399, ZN => n6374);
   U6527 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx3x, B1 => 
                           ashr_25xAx2x, B2 => n7399, ZN => n6177);
   U6528 : AOI22_X1 port map( A1 => n7404, A2 => n6374, B1 => n6177, B2 => 
                           n7402, ZN => n6465);
   U6529 : INV_X1 port map( A => n5685, ZN => n5967);
   U6530 : OAI21_X1 port map( B1 => n7399, B2 => ashr_25xAx1x, A => n5967, ZN 
                           => n6176);
   U6531 : NOR2_X1 port map( A1 => n5711, A2 => n6176, ZN => n6467);
   U6532 : AOI22_X1 port map( A1 => n7311, A2 => n6465, B1 => n6467, B2 => 
                           n7309, ZN => n6643);
   U6533 : NOR2_X1 port map( A1 => n5689, A2 => n5692, ZN => n5725);
   U6534 : NOR2_X1 port map( A1 => n7192, A2 => n5710, ZN => n5686);
   U6535 : AND2_X1 port map( A1 => n5725, A2 => n5686, ZN => n7348);
   U6536 : NAND2_X1 port map( A1 => n7376, A2 => n7348, ZN => n7004);
   U6537 : OAI22_X1 port map( A1 => n6309, A2 => n7427, B1 => n6643, B2 => 
                           n7004, ZN => n5736);
   U6538 : INV_X1 port map( A => intadd_25xBx0x, ZN => n6962);
   U6539 : AOI22_X1 port map( A1 => n7414, A2 => intadd_26xAx4x, B1 => 
                           intadd_26xAx5x, B2 => n7412, ZN => n6203);
   U6540 : CLKBUF_X1 port map( A => n7412, Z => n7130);
   U6541 : OAI22_X1 port map( A1 => n7130, A2 => intadd_26xAx6x, B1 => 
                           intadd_26xAx7x, B2 => n7414, ZN => n6206);
   U6542 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6203, B1 => n6206, 
                           B2 => n7259, ZN => n6482);
   U6543 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx27x, B1 => 
                           ashr_25xAx28x, B2 => n7412, ZN => n6202);
   U6544 : OAI22_X1 port map( A1 => n7130, A2 => n7129, B1 => n7160, B2 => 
                           n7414, ZN => n6205);
   U6545 : INV_X1 port map( A => n6205, ZN => n5687);
   U6546 : MUX2_X1 port map( A => n6202, B => n5687, S => intadd_29xBx0x, Z => 
                           n6074);
   U6547 : AOI22_X1 port map( A1 => n6962, A2 => n6482, B1 => n6074, B2 => 
                           n6456, ZN => n6637);
   U6548 : NOR2_X1 port map( A1 => intadd_29xBx2x, A2 => n6456, ZN => n6417);
   U6549 : NOR2_X1 port map( A1 => n7130, A2 => n7435, ZN => n6207);
   U6550 : CLKBUF_X1 port map( A => n7259, Z => n7231);
   U6551 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx29x, B1 => 
                           ashr_25xAx30x, B2 => n7412, ZN => n6201);
   U6552 : NOR2_X1 port map( A1 => n7231, A2 => n6201, ZN => n5691);
   U6553 : AOI21_X1 port map( B1 => n6207, B2 => n7231, A => n5691, ZN => n7286
                           );
   U6554 : INV_X1 port map( A => n7286, ZN => n5688);
   U6555 : AOI22_X1 port map( A1 => n7236, A2 => n6637, B1 => n6417, B2 => 
                           n5688, ZN => n6279);
   U6556 : NOR2_X1 port map( A1 => n5715, A2 => n5689, ZN => n5728);
   U6557 : NAND2_X1 port map( A1 => n5690, A2 => n5728, ZN => n6072);
   U6558 : NOR2_X1 port map( A1 => ashr_25xSHx4x, A2 => n6072, ZN => n7166);
   U6559 : INV_X1 port map( A => n7166, ZN => n7220);
   U6560 : NOR2_X1 port map( A1 => intadd_29xBx0x, A2 => n7435, ZN => n6343);
   U6561 : NOR2_X1 port map( A1 => n6343, A2 => n5691, ZN => n6046);
   U6562 : NAND2_X1 port map( A1 => n7413, A2 => n6811, ZN => n6246);
   U6563 : OAI21_X1 port map( B1 => n6046, B2 => n6456, A => n6246, ZN => n6634
                           );
   U6564 : AOI22_X1 port map( A1 => n7236, A2 => n6637, B1 => n6634, B2 => 
                           ashr_25xSHx3x, ZN => n6278);
   U6565 : NOR3_X1 port map( A1 => n5699, A2 => n5692, A3 => n5698, ZN => n5709
                           );
   U6566 : NAND2_X1 port map( A1 => n6022, A2 => n5709, ZN => n6047);
   U6567 : INV_X1 port map( A => n6047, ZN => n6247);
   U6568 : OAI21_X1 port map( B1 => n7331, B2 => n7413, A => n6247, ZN => n7329
                           );
   U6569 : AOI21_X1 port map( B1 => n7331, B2 => n6278, A => n7329, ZN => n5707
                           );
   U6570 : INV_X1 port map( A => intadd_25xSUMx19x, ZN => n5696);
   U6571 : NAND2_X1 port map( A1 => n5694, A2 => n5693, ZN => n7384);
   U6572 : NAND2_X1 port map( A1 => intadd_26xAx4x, A2 => add_x_26xBx21x, ZN =>
                           n5695);
   U6573 : NOR3_X1 port map( A1 => n5697, A2 => n5699, A3 => n5715, ZN => n7127
                           );
   U6574 : CLKBUF_X1 port map( A => n7127, Z => n7410);
   U6575 : INV_X1 port map( A => n7410, ZN => n7316);
   U6576 : OAI22_X1 port map( A1 => n5696, A2 => n7384, B1 => n5695, B2 => 
                           n7316, ZN => n5706);
   U6577 : NOR3_X1 port map( A1 => n5698, A2 => n5716, A3 => n5710, ZN => n5968
                           );
   U6578 : INV_X1 port map( A => n5968, ZN => n7398);
   U6579 : NOR3_X1 port map( A1 => n5699, A2 => n5698, A3 => n5697, ZN => n5700
                           );
   U6580 : AND2_X1 port map( A1 => n6020, A2 => n5700, ZN => n7327);
   U6581 : CLKBUF_X1 port map( A => n7327, Z => n7073);
   U6582 : INV_X1 port map( A => n7073, ZN => n7397);
   U6583 : AOI211_X1 port map( C1 => n7398, C2 => n7397, A => ashr_25xAx21x, B 
                           => n7477, ZN => n5705);
   U6584 : NOR2_X1 port map( A1 => n5702, A2 => n5701, ZN => n5703);
   U6585 : NOR2_X1 port map( A1 => n5703, A2 => n7251, ZN => n7227);
   U6586 : OAI22_X1 port map( A1 => intadd_26xBx4x, A2 => n7227, B1 => n7118, 
                           B2 => n5881, ZN => n5704);
   U6587 : NOR4_X1 port map( A1 => n5707, A2 => n5706, A3 => n5705, A4 => n5704
                           , ZN => n5734);
   U6588 : NOR2_X1 port map( A1 => ashr_25xSHx4x, A2 => n5715, ZN => n5708);
   U6589 : AND2_X1 port map( A1 => n5725, A2 => n5708, ZN => n7420);
   U6590 : AND2_X1 port map( A1 => n7420, A2 => ashr_25xSHx3x, ZN => n7431);
   U6591 : AOI22_X1 port map( A1 => n7333, A2 => intadd_27xAx2x, B1 => 
                           intadd_27xAx1x, B2 => n7412, ZN => n6724);
   U6592 : AOI22_X1 port map( A1 => n7333, A2 => intadd_27xAx0x, B1 => n6528, 
                           B2 => n7412, ZN => n6558);
   U6593 : AOI22_X1 port map( A1 => n7418, A2 => n6724, B1 => n6558, B2 => 
                           n7259, ZN => n6812);
   U6594 : AOI22_X1 port map( A1 => n7414, A2 => n6481, B1 => n6419, B2 => 
                           n7412, ZN => n6557);
   U6595 : AOI22_X1 port map( A1 => n7414, A2 => n6399, B1 => n6330, B2 => 
                           n7412, ZN => n6367);
   U6596 : AOI22_X1 port map( A1 => n7418, A2 => n6557, B1 => n6367, B2 => 
                           n7259, ZN => n6458);
   U6597 : AOI22_X1 port map( A1 => n6962, A2 => n6812, B1 => n6458, B2 => 
                           n6456, ZN => n6647);
   U6598 : INV_X1 port map( A => n5709, ZN => n7385);
   U6599 : NOR2_X1 port map( A1 => n7385, A2 => n5710, ZN => n6325);
   U6600 : INV_X1 port map( A => n6325, ZN => n6386);
   U6601 : INV_X1 port map( A => n7353, ZN => n7190);
   U6602 : NAND2_X1 port map( A1 => n7413, A2 => n5711, ZN => n6676);
   U6603 : NAND2_X1 port map( A1 => n6676, A2 => n5712, ZN => n6651);
   U6604 : AND2_X1 port map( A1 => n7376, A2 => n6642, ZN => n5714);
   U6605 : NOR2_X1 port map( A1 => n7435, A2 => n7376, ZN => n6520);
   U6606 : NAND2_X1 port map( A1 => n6520, A2 => n6900, ZN => n6350);
   U6607 : INV_X1 port map( A => n6350, ZN => n5713);
   U6608 : AOI211_X1 port map( C1 => n6365, C2 => n6651, A => n5714, B => n5713
                           , ZN => n6289);
   U6609 : INV_X1 port map( A => n7420, ZN => n7343);
   U6610 : NOR2_X1 port map( A1 => ashr_25xSHx3x, A2 => n7343, ZN => n7018);
   U6611 : AOI22_X1 port map( A1 => n7333, A2 => intadd_26xAx4x, B1 => 
                           intadd_26xAx3x, B2 => n7412, ZN => n7015);
   U6612 : AOI22_X1 port map( A1 => n7333, A2 => intadd_26xAx2x, B1 => 
                           intadd_26xAx1x, B2 => n7412, ZN => n6895);
   U6613 : AOI22_X1 port map( A1 => n7418, A2 => n7015, B1 => n6895, B2 => 
                           n7416, ZN => n7093);
   U6614 : AOI22_X1 port map( A1 => n7333, A2 => intadd_26xAx0x, B1 => n6774, 
                           B2 => n7412, ZN => n6894);
   U6615 : AOI22_X1 port map( A1 => n7333, A2 => n6766, B1 => intadd_27xAx3x, 
                           B2 => n7412, ZN => n6725);
   U6616 : AOI22_X1 port map( A1 => n7418, A2 => n6894, B1 => n6725, B2 => 
                           n7416, ZN => n6813);
   U6617 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n7093, B1 => n6813, 
                           B2 => n6456, ZN => n7263);
   U6618 : INV_X1 port map( A => n7320, ZN => n7386);
   U6619 : INV_X1 port map( A => n7410, ZN => n7255);
   U6620 : INV_X1 port map( A => n5716, ZN => n5717);
   U6621 : NAND2_X1 port map( A1 => n6020, A2 => n5717, ZN => n5718);
   U6622 : NOR2_X1 port map( A1 => n5719, A2 => n5718, ZN => n7253);
   U6623 : AOI221_X1 port map( B1 => n7327, B2 => n7477, C1 => n7253, C2 => 
                           n5720, A => n7251, ZN => n5721);
   U6624 : OAI221_X1 port map( B1 => intadd_26xBx4x, B2 => n7386, C1 => 
                           add_x_26xBx21x, C2 => n7255, A => n5721, ZN => n5722
                           );
   U6625 : AOI22_X1 port map( A1 => n7018, A2 => n7263, B1 => ashr_25xAx21x, B2
                           => n5722, ZN => n5723);
   U6626 : OAI221_X1 port map( B1 => n7190, B2 => n7192, C1 => n7190, C2 => 
                           n6289, A => n5723, ZN => n5732);
   U6627 : INV_X1 port map( A => n7309, ZN => n6941);
   U6628 : INV_X1 port map( A => n7267, ZN => n7268);
   U6629 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx13x, B1 => 
                           ashr_25xAx12x, B2 => n7086, ZN => n6730);
   U6630 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx11x, B1 => 
                           ashr_25xAx10x, B2 => n7086, ZN => n6566);
   U6631 : AOI22_X1 port map( A1 => n7404, A2 => n6730, B1 => n6566, B2 => 
                           n7402, ZN => n6822);
   U6632 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx9x, B1 => 
                           ashr_25xAx8x, B2 => n7086, ZN => n6565);
   U6633 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx7x, B1 => 
                           ashr_25xAx6x, B2 => n7086, ZN => n6375);
   U6634 : AOI22_X1 port map( A1 => n7404, A2 => n6565, B1 => n6375, B2 => 
                           n7402, ZN => n6466);
   U6635 : AOI22_X1 port map( A1 => n6941, A2 => n6822, B1 => n6466, B2 => 
                           n6900, ZN => n6644);
   U6636 : AND2_X1 port map( A1 => n6020, A2 => n7192, ZN => n5724);
   U6637 : AND2_X1 port map( A1 => n5725, A2 => n5724, ZN => n7409);
   U6638 : AND2_X1 port map( A1 => n7409, A2 => n7207, ZN => n7394);
   U6639 : INV_X1 port map( A => n7394, ZN => n7314);
   U6640 : AND2_X1 port map( A1 => n7409, A2 => n7376, ZN => n7307);
   U6641 : AOI22_X1 port map( A1 => n7268, A2 => intadd_26xAx4x, B1 => 
                           intadd_26xAx3x, B2 => n7086, ZN => n6998);
   U6642 : AOI22_X1 port map( A1 => n7268, A2 => intadd_26xAx2x, B1 => 
                           intadd_26xAx1x, B2 => n7399, ZN => n6899);
   U6643 : AOI22_X1 port map( A1 => n7404, A2 => n6998, B1 => n6899, B2 => 
                           n7402, ZN => n7088);
   U6644 : AOI22_X1 port map( A1 => n7268, A2 => intadd_26xAx0x, B1 => n6774, 
                           B2 => n7399, ZN => n6898);
   U6645 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx15x, B1 => 
                           ashr_25xAx14x, B2 => n7086, ZN => n6731);
   U6646 : INV_X1 port map( A => n6731, ZN => n5726);
   U6647 : AOI22_X1 port map( A1 => n7404, A2 => n6898, B1 => n5726, B2 => 
                           n7402, ZN => n6821);
   U6648 : AOI22_X1 port map( A1 => n6941, A2 => n7088, B1 => n6821, B2 => 
                           n7309, ZN => n7271);
   U6649 : AND2_X1 port map( A1 => n5728, A2 => n5727, ZN => n5729);
   U6650 : AND2_X1 port map( A1 => n5729, A2 => ashr_25xSHx4x, ZN => n7352);
   U6651 : NAND2_X1 port map( A1 => n7236, A2 => n7352, ZN => n6929);
   U6652 : INV_X1 port map( A => n6929, ZN => n7000);
   U6653 : AOI22_X1 port map( A1 => n7414, A2 => n6048, B1 => n6251, B2 => 
                           n7412, ZN => n6366);
   U6654 : AOI22_X1 port map( A1 => n7414, A2 => intadd_29xAx2x, B1 => 
                           intadd_29xAx1x, B2 => n7412, ZN => n6160);
   U6655 : AOI22_X1 port map( A1 => n7418, A2 => n6366, B1 => n6160, B2 => 
                           n7259, ZN => n6457);
   U6656 : AOI21_X1 port map( B1 => n7414, B2 => intadd_29xAx0x, A => n5972, ZN
                           => n6159);
   U6657 : NAND2_X1 port map( A1 => n7418, A2 => n6159, ZN => n6459);
   U6658 : AOI22_X1 port map( A1 => n6962, A2 => n6457, B1 => n6459, B2 => 
                           n6456, ZN => n6646);
   U6659 : AOI22_X1 port map( A1 => n7307, A2 => n7271, B1 => n7000, B2 => 
                           n6646, ZN => n5730);
   U6660 : OAI21_X1 port map( B1 => n6644, B2 => n7314, A => n5730, ZN => n5731
                           );
   U6661 : AOI211_X1 port map( C1 => n7431, C2 => n6647, A => n5732, B => n5731
                           , ZN => n5733);
   U6662 : OAI211_X1 port map( C1 => n6279, C2 => n7220, A => n5734, B => n5733
                           , ZN => n5735);
   U6663 : AOI211_X1 port map( C1 => DP_OP_719J14_125_1055xn90, C2 => n7159, A 
                           => n5736, B => n5735, ZN => n5738);
   U6664 : NAND2_X1 port map( A1 => n7520, A2 => n6044, ZN => n6717);
   U6665 : INV_X1 port map( A => n6717, ZN => n7029);
   U6666 : INV_X1 port map( A => n7029, ZN => n7533);
   U6667 : INV_X1 port map( A => n6597, ZN => n7439);
   U6668 : OAI22_X1 port map( A1 => n5738, A2 => n7533, B1 => n5737, B2 => 
                           n7439, ZN => IF_ISAxN10958);
   U6669 : NAND2_X1 port map( A1 => ashr_25xAx0x, A2 => n7130, ZN => 
                           intadd_29xCI);
   U6670 : OR4_X1 port map( A1 => IF_ISAxsection_2_port, A2 => n5749, A3 => 
                           n5748, A4 => n5739, ZN => n5787);
   U6671 : INV_X1 port map( A => n5787, ZN => n5943);
   U6672 : NOR4_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(2), A2 => n6361, 
                           A3 => n5749, A4 => n5740, ZN => n5742);
   U6673 : AND2_X1 port map( A1 => n5742, A2 => n5741, ZN => n5941);
   U6674 : INV_X1 port map( A => n5941, ZN => n5865);
   U6675 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(12), A2 => n5742
                           , ZN => n5930);
   U6676 : OAI22_X1 port map( A1 => n5746, A2 => n5865, B1 => n5930, B2 => 
                           n5743, ZN => n5752);
   U6677 : OAI211_X1 port map( C1 => n5744, C2 => n5930, A => n5755, B => n7535
                           , ZN => n5745);
   U6678 : AOI21_X1 port map( B1 => n5746, B2 => n5941, A => n5745, ZN => n5750
                           );
   U6679 : NOR3_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(2), A2 => 
                           fromMemoryPortxLOADEDDATAx(4), A3 => n5747, ZN => 
                           n5939);
   U6680 : NOR4_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(3), A2 => 
                           IF_ISAxsection_2_port, A3 => n5749, A4 => n5748, ZN 
                           => n5754);
   U6681 : NOR2_X2 port map( A1 => n5939, A2 => n5754, ZN => n5932);
   U6682 : OAI22_X1 port map( A1 => n5750, A2 => n7542, B1 => intadd_29xSUMx0x,
                           B2 => n5932, ZN => n5751);
   U6683 : AOI221_X1 port map( B1 => n5943, B2 => n6068, C1 => n5752, C2 => 
                           n6068, A => n5751, ZN => n5753);
   U6684 : NAND2_X1 port map( A1 => n7458, A2 => n7523, ZN => n5756);
   U6685 : OAI22_X1 port map( A1 => n5753, A2 => n5952, B1 => n7542, B2 => 
                           n5756, ZN => n7626);
   U6686 : NAND2_X1 port map( A1 => n5827, A2 => n5754, ZN => n5831);
   U6687 : NOR2_X1 port map( A1 => n5936, A2 => n5930, ZN => n5824);
   U6688 : AND2_X1 port map( A1 => n5755, A2 => n7535, ZN => n5757);
   U6689 : OAI21_X1 port map( B1 => n5936, B2 => n5757, A => n5756, ZN => n5822
                           );
   U6690 : AOI22_X1 port map( A1 => n5824, A2 => n5758, B1 => n7546, B2 => 
                           n5822, ZN => n5762);
   U6691 : INV_X1 port map( A => n5939, ZN => n5826);
   U6692 : OAI22_X1 port map( A1 => intadd_29xSUMx1x, A2 => n5826, B1 => n5865,
                           B2 => n5759, ZN => n5760);
   U6693 : OAI221_X1 port map( B1 => n5760, B2 => n5943, C1 => n5760, C2 => 
                           intadd_25xSUMx0x, A => n5827, ZN => n5761);
   U6694 : OAI211_X1 port map( C1 => intadd_29xSUMx1x, C2 => n5831, A => n5762,
                           B => n5761, ZN => n7625);
   U6695 : AOI22_X1 port map( A1 => n5764, A2 => n5824, B1 => n5763, B2 => 
                           n5822, ZN => n5768);
   U6696 : INV_X1 port map( A => n5941, ZN => n5929);
   U6697 : OAI22_X1 port map( A1 => intadd_29xSUMx2x, A2 => n5826, B1 => n5929,
                           B2 => n5765, ZN => n5766);
   U6698 : OAI221_X1 port map( B1 => n5766, B2 => n5943, C1 => n5766, C2 => 
                           intadd_25xSUMx1x, A => n5827, ZN => n5767);
   U6699 : OAI211_X1 port map( C1 => intadd_29xSUMx2x, C2 => n5831, A => n5768,
                           B => n5767, ZN => n7624);
   U6700 : AOI22_X1 port map( A1 => n5770, A2 => n5824, B1 => n5769, B2 => 
                           n5822, ZN => n5774);
   U6701 : OAI22_X1 port map( A1 => n5775, A2 => n5826, B1 => n5865, B2 => 
                           n5771, ZN => n5772);
   U6702 : OAI221_X1 port map( B1 => n5772, B2 => n5943, C1 => n5772, C2 => 
                           intadd_25xSUMx2x, A => n5827, ZN => n5773);
   U6703 : OAI211_X1 port map( C1 => n5775, C2 => n5831, A => n5774, B => n5773
                           , ZN => n7623);
   U6704 : INV_X1 port map( A => n5822, ZN => n5947);
   U6705 : INV_X1 port map( A => n5824, ZN => n5944);
   U6706 : INV_X1 port map( A => n5932, ZN => n5911);
   U6707 : AOI222_X1 port map( A1 => n5777, A2 => n5911, B1 => n5941, B2 => 
                           n5776, C1 => n5943, C2 => intadd_25xSUMx3x, ZN => 
                           n5778);
   U6708 : OAI222_X1 port map( A1 => n5780, A2 => n5947, B1 => n5944, B2 => 
                           n5779, C1 => n5952, C2 => n5778, ZN => n7622);
   U6709 : INV_X1 port map( A => n5831, ZN => n5950);
   U6710 : AOI22_X1 port map( A1 => n5782, A2 => n5950, B1 => n6335, B2 => 
                           n5822, ZN => n5785);
   U6711 : INV_X1 port map( A => intadd_25xSUMx4x, ZN => n6318);
   U6712 : OAI22_X1 port map( A1 => n5787, A2 => n6318, B1 => n5865, B2 => 
                           n5781, ZN => n5783);
   U6713 : OAI221_X1 port map( B1 => n5783, B2 => n5939, C1 => n5783, C2 => 
                           n5782, A => n5827, ZN => n5784);
   U6714 : OAI211_X1 port map( C1 => n5786, C2 => n5944, A => n5785, B => n5784
                           , ZN => n7621);
   U6715 : INV_X1 port map( A => n5787, ZN => n5935);
   U6716 : AOI22_X1 port map( A1 => n5935, A2 => intadd_25xSUMx5x, B1 => n5941,
                           B2 => n5788, ZN => n5789);
   U6717 : OAI21_X1 port map( B1 => n5790, B2 => n5930, A => n5789, ZN => n5791
                           );
   U6718 : AOI21_X1 port map( B1 => n5792, B2 => n5911, A => n5791, ZN => n5793
                           );
   U6719 : OAI22_X1 port map( A1 => n5947, A2 => n6393, B1 => n5793, B2 => 
                           n5952, ZN => n7620);
   U6720 : AOI22_X1 port map( A1 => n5950, A2 => n5794, B1 => n6438, B2 => 
                           n5822, ZN => n5799);
   U6721 : INV_X1 port map( A => n5794, ZN => n5796);
   U6722 : OAI22_X1 port map( A1 => n5796, A2 => n5826, B1 => n5865, B2 => 
                           n5795, ZN => n5797);
   U6723 : OAI221_X1 port map( B1 => n5797, B2 => n5943, C1 => n5797, C2 => 
                           intadd_25xSUMx6x, A => n5827, ZN => n5798);
   U6724 : OAI211_X1 port map( C1 => n5800, C2 => n5944, A => n5799, B => n5798
                           , ZN => n7619);
   U6725 : NOR2_X1 port map( A1 => n5801, A2 => n5930, ZN => n5805);
   U6726 : OAI22_X1 port map( A1 => n5932, A2 => n5803, B1 => n5865, B2 => 
                           n5802, ZN => n5804);
   U6727 : AOI211_X1 port map( C1 => intadd_25xSUMx7x, C2 => n5935, A => n5805,
                           B => n5804, ZN => n5806);
   U6728 : OAI22_X1 port map( A1 => n5947, A2 => n6472, B1 => n5806, B2 => 
                           n5952, ZN => n7618);
   U6729 : INV_X1 port map( A => n5808, ZN => n5807);
   U6730 : AOI22_X1 port map( A1 => n5807, A2 => n5950, B1 => n6507, B2 => 
                           n5822, ZN => n5812);
   U6731 : OAI22_X1 port map( A1 => n5929, A2 => n5809, B1 => n5826, B2 => 
                           n5808, ZN => n5810);
   U6732 : OAI221_X1 port map( B1 => n5810, B2 => n5943, C1 => n5810, C2 => 
                           intadd_25xSUMx8x, A => n5827, ZN => n5811);
   U6733 : OAI211_X1 port map( C1 => n5813, C2 => n5944, A => n5812, B => n5811
                           , ZN => n7617);
   U6734 : NAND2_X1 port map( A1 => n6528, A2 => n5814, ZN => n5815);
   U6735 : AOI21_X1 port map( B1 => n5816, B2 => n5815, A => n6540, ZN => 
                           intadd_27xCI);
   U6736 : NOR2_X1 port map( A1 => n5932, A2 => intadd_27xSUMx0x, ZN => n5820);
   U6737 : OAI22_X1 port map( A1 => n5818, A2 => n5930, B1 => n5865, B2 => 
                           n5817, ZN => n5819);
   U6738 : AOI211_X1 port map( C1 => intadd_25xSUMx9x, C2 => n5943, A => n5820,
                           B => n5819, ZN => n5821);
   U6739 : OAI22_X1 port map( A1 => n5947, A2 => n6572, B1 => n5821, B2 => 
                           n5952, ZN => n7616);
   U6740 : AOI22_X1 port map( A1 => n5824, A2 => n5823, B1 => n6612, B2 => 
                           n5822, ZN => n5830);
   U6741 : OAI22_X1 port map( A1 => intadd_27xSUMx1x, A2 => n5826, B1 => n5865,
                           B2 => n5825, ZN => n5828);
   U6742 : OAI221_X1 port map( B1 => n5828, B2 => n5943, C1 => n5828, C2 => 
                           intadd_25xSUMx10x, A => n5827, ZN => n5829);
   U6743 : OAI211_X1 port map( C1 => intadd_27xSUMx1x, C2 => n5831, A => n5830,
                           B => n5829, ZN => n7615);
   U6744 : NOR2_X1 port map( A1 => n5929, A2 => n5832, ZN => n5835);
   U6745 : OAI22_X1 port map( A1 => n5932, A2 => intadd_27xSUMx2x, B1 => n5833,
                           B2 => n5930, ZN => n5834);
   U6746 : AOI211_X1 port map( C1 => intadd_25xSUMx11x, C2 => n5935, A => n5835
                           , B => n5834, ZN => n5836);
   U6747 : OAI22_X1 port map( A1 => n5947, A2 => n5837, B1 => n5836, B2 => 
                           n5952, ZN => n7614);
   U6748 : OAI22_X1 port map( A1 => n5932, A2 => intadd_27xSUMx3x, B1 => n5865,
                           B2 => n5838, ZN => n5839);
   U6749 : AOI21_X1 port map( B1 => n5943, B2 => intadd_25xSUMx12x, A => n5839,
                           ZN => n5840);
   U6750 : OAI222_X1 port map( A1 => n6687, A2 => n5947, B1 => n5944, B2 => 
                           n5841, C1 => n5952, C2 => n5840, ZN => n7613);
   U6751 : AND2_X1 port map( A1 => n5911, A2 => n5842, ZN => n5846);
   U6752 : OAI22_X1 port map( A1 => n5844, A2 => n5930, B1 => n5865, B2 => 
                           n5843, ZN => n5845);
   U6753 : AOI211_X1 port map( C1 => n5943, C2 => intadd_25xSUMx13x, A => n5846
                           , B => n5845, ZN => n5847);
   U6754 : OAI22_X1 port map( A1 => n5947, A2 => n6742, B1 => n5847, B2 => 
                           n5952, ZN => n7612);
   U6755 : AND2_X1 port map( A1 => n5911, A2 => n5848, ZN => n5852);
   U6756 : OAI22_X1 port map( A1 => n5850, A2 => n5930, B1 => n5865, B2 => 
                           n5849, ZN => n5851);
   U6757 : AOI211_X1 port map( C1 => n5943, C2 => intadd_25xSUMx14x, A => n5852
                           , B => n5851, ZN => n5853);
   U6758 : OAI22_X1 port map( A1 => n5947, A2 => n5854, B1 => n5853, B2 => 
                           n5952, ZN => n7611);
   U6759 : AOI22_X1 port map( A1 => ashr_25xAx16x, A2 => add_x_26xBx16x, B1 => 
                           n6775, B2 => n5855, ZN => intadd_26xCI);
   U6760 : OAI22_X1 port map( A1 => n5932, A2 => intadd_26xSUMx0x, B1 => n5865,
                           B2 => n5856, ZN => n5857);
   U6761 : AOI21_X1 port map( B1 => n5943, B2 => intadd_25xSUMx15x, A => n5857,
                           ZN => n5858);
   U6762 : OAI222_X1 port map( A1 => n6805, A2 => n5947, B1 => n5944, B2 => 
                           n5859, C1 => n5952, C2 => n5858, ZN => n7610);
   U6763 : OAI22_X1 port map( A1 => n5932, A2 => intadd_26xSUMx1x, B1 => n5865,
                           B2 => n5860, ZN => n5861);
   U6764 : AOI21_X1 port map( B1 => n5943, B2 => intadd_25xSUMx16x, A => n5861,
                           ZN => n5862);
   U6765 : OAI222_X1 port map( A1 => n6859, A2 => n5947, B1 => n5944, B2 => 
                           n5863, C1 => n5952, C2 => n5862, ZN => n7609);
   U6766 : NOR2_X1 port map( A1 => n5932, A2 => intadd_26xSUMx2x, ZN => n5868);
   U6767 : OAI22_X1 port map( A1 => n5866, A2 => n5930, B1 => n5865, B2 => 
                           n5864, ZN => n5867);
   U6768 : AOI211_X1 port map( C1 => intadd_25xSUMx17x, C2 => n5935, A => n5868
                           , B => n5867, ZN => n5869);
   U6769 : OAI22_X1 port map( A1 => n5947, A2 => n6893, B1 => n5869, B2 => 
                           n5952, ZN => n7608);
   U6770 : NOR2_X1 port map( A1 => n5932, A2 => intadd_26xSUMx3x, ZN => n5873);
   U6771 : OAI22_X1 port map( A1 => n5871, A2 => n5930, B1 => n5929, B2 => 
                           n5870, ZN => n5872);
   U6772 : AOI211_X1 port map( C1 => intadd_25xSUMx18x, C2 => n5935, A => n5873
                           , B => n5872, ZN => n5874);
   U6773 : OAI22_X1 port map( A1 => n5947, A2 => n5875, B1 => n5874, B2 => 
                           n5936, ZN => n7607);
   U6774 : NOR2_X1 port map( A1 => n5929, A2 => n5876, ZN => n5879);
   U6775 : OAI22_X1 port map( A1 => n5932, A2 => intadd_26xSUMx4x, B1 => n5877,
                           B2 => n5930, ZN => n5878);
   U6776 : AOI211_X1 port map( C1 => intadd_25xSUMx19x, C2 => n5935, A => n5879
                           , B => n5878, ZN => n5880);
   U6777 : OAI22_X1 port map( A1 => n5947, A2 => n5881, B1 => n5880, B2 => 
                           n5936, ZN => n7606);
   U6778 : NOR2_X1 port map( A1 => n5929, A2 => n5882, ZN => n5885);
   U6779 : OAI22_X1 port map( A1 => n5932, A2 => intadd_26xSUMx5x, B1 => n5883,
                           B2 => n5930, ZN => n5884);
   U6780 : AOI211_X1 port map( C1 => intadd_25xSUMx20x, C2 => n5935, A => n5885
                           , B => n5884, ZN => n5886);
   U6781 : OAI22_X1 port map( A1 => n5947, A2 => n6983, B1 => n5886, B2 => 
                           n5936, ZN => n7605);
   U6782 : OAI22_X1 port map( A1 => n5932, A2 => intadd_26xSUMx6x, B1 => n5929,
                           B2 => n5887, ZN => n5888);
   U6783 : AOI21_X1 port map( B1 => n5943, B2 => intadd_25xSUMx21x, A => n5888,
                           ZN => n5889);
   U6784 : OAI222_X1 port map( A1 => n5891, A2 => n5947, B1 => n5944, B2 => 
                           n5890, C1 => n5952, C2 => n5889, ZN => n7604);
   U6785 : NOR2_X1 port map( A1 => n5929, A2 => n5892, ZN => n5895);
   U6786 : OAI22_X1 port map( A1 => n5932, A2 => intadd_26xSUMx7x, B1 => n5893,
                           B2 => n5930, ZN => n5894);
   U6787 : AOI211_X1 port map( C1 => intadd_25xSUMx22x, C2 => n5935, A => n5895
                           , B => n5894, ZN => n5896);
   U6788 : OAI22_X1 port map( A1 => n5947, A2 => n5897, B1 => n5896, B2 => 
                           n5936, ZN => n7603);
   U6789 : NOR2_X1 port map( A1 => n5929, A2 => n5898, ZN => n5902);
   U6790 : OAI22_X1 port map( A1 => n5932, A2 => n5900, B1 => n5899, B2 => 
                           n5930, ZN => n5901);
   U6791 : AOI211_X1 port map( C1 => intadd_25xSUMx23x, C2 => n5935, A => n5902
                           , B => n5901, ZN => n5903);
   U6792 : OAI22_X1 port map( A1 => n5947, A2 => n7079, B1 => n5903, B2 => 
                           n5936, ZN => n7602);
   U6793 : NOR2_X1 port map( A1 => n5929, A2 => n5904, ZN => n5908);
   U6794 : OAI22_X1 port map( A1 => n5932, A2 => n5906, B1 => n5905, B2 => 
                           n5930, ZN => n5907);
   U6795 : AOI211_X1 port map( C1 => intadd_25xSUMx24x, C2 => n5935, A => n5908
                           , B => n5907, ZN => n5909);
   U6796 : OAI22_X1 port map( A1 => n5947, A2 => n7117, B1 => n5909, B2 => 
                           n5936, ZN => n7601);
   U6797 : AOI222_X1 port map( A1 => n5912, A2 => n5911, B1 => n5941, B2 => 
                           n5910, C1 => n5943, C2 => intadd_25xSUMx25x, ZN => 
                           n5913);
   U6798 : OAI222_X1 port map( A1 => n5915, A2 => n5947, B1 => n5944, B2 => 
                           n5914, C1 => n5936, C2 => n5913, ZN => n7600);
   U6799 : OAI22_X1 port map( A1 => n7182, A2 => n5916, B1 => ashr_25xAx27x, B2
                           => add_x_26xBx27x, ZN => intadd_28xCI);
   U6800 : NOR2_X1 port map( A1 => n5929, A2 => n5917, ZN => n5920);
   U6801 : OAI22_X1 port map( A1 => n5932, A2 => intadd_28xSUMx0x, B1 => n5918,
                           B2 => n5930, ZN => n5919);
   U6802 : AOI211_X1 port map( C1 => intadd_25xSUMx26x, C2 => n5935, A => n5920
                           , B => n5919, ZN => n5921);
   U6803 : OAI22_X1 port map( A1 => n5947, A2 => n5922, B1 => n5921, B2 => 
                           n5936, ZN => n7599);
   U6804 : OAI22_X1 port map( A1 => n5932, A2 => intadd_28xSUMx1x, B1 => n5929,
                           B2 => n5923, ZN => n5924);
   U6805 : AOI21_X1 port map( B1 => n5943, B2 => intadd_25xSUMx27x, A => n5924,
                           ZN => n5925);
   U6806 : OAI222_X1 port map( A1 => n5927, A2 => n5947, B1 => n5944, B2 => 
                           n5926, C1 => n5952, C2 => n5925, ZN => n7598);
   U6807 : INV_X1 port map( A => n7361, ZN => n5938);
   U6808 : NOR2_X1 port map( A1 => n5929, A2 => n5928, ZN => n5934);
   U6809 : OAI22_X1 port map( A1 => n5932, A2 => intadd_28xSUMx2x, B1 => n5931,
                           B2 => n5930, ZN => n5933);
   U6810 : AOI211_X1 port map( C1 => intadd_25xSUMx28x, C2 => n5935, A => n5934
                           , B => n5933, ZN => n5937);
   U6811 : OAI22_X1 port map( A1 => n5947, A2 => n5938, B1 => n5937, B2 => 
                           n5936, ZN => n7597);
   U6812 : AOI222_X1 port map( A1 => n5943, A2 => n5942, B1 => n5941, B2 => 
                           n5940, C1 => n5939, C2 => n5949, ZN => n5953);
   U6813 : OAI22_X1 port map( A1 => n5947, A2 => n5946, B1 => n5945, B2 => 
                           n5944, ZN => n5948);
   U6814 : AOI21_X1 port map( B1 => n5950, B2 => n5949, A => n5948, ZN => n5951
                           );
   U6815 : OAI21_X1 port map( B1 => n5953, B2 => n5952, A => n5951, ZN => n7596
                           );
   U6816 : NOR3_X1 port map( A1 => n5955, A2 => n5954, A3 => n5958, ZN => n7594
                           );
   U6817 : AOI211_X1 port map( C1 => fromMemoryPortxLOADEDDATAx(5), C2 => 
                           fromMemoryPortxLOADEDDATAx(14), A => n5958, B => 
                           fromMemoryPortxLOADEDDATAx(13), ZN => n5956);
   U6818 : AND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(12), A2 => n5956,
                           ZN => n7593);
   U6819 : NOR2_X1 port map( A1 => n7538, A2 => n7535, ZN => n5957);
   U6820 : AOI21_X1 port map( B1 => n5957, B2 => n7520, A => n5956, ZN => n7592
                           );
   U6821 : INV_X1 port map( A => n5958, ZN => n5960);
   U6822 : NAND2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(5), A2 => n5960,
                           ZN => n5959);
   U6823 : INV_X1 port map( A => n5959, ZN => n7595);
   U6824 : NOR2_X1 port map( A1 => n7209, A2 => n5959, ZN => n7591);
   U6825 : NOR2_X1 port map( A1 => n7192, A2 => n5959, ZN => n7590);
   U6826 : NOR2_X1 port map( A1 => n7311, A2 => n5959, ZN => n7589);
   U6827 : NOR2_X1 port map( A1 => n7376, A2 => n5959, ZN => n7588);
   U6828 : NOR2_X1 port map( A1 => n7304, A2 => n5959, ZN => n7587);
   U6829 : NOR2_X1 port map( A1 => rst, A2 => IF_ISAxsection_0_port, ZN => 
                           n7556);
   U6830 : INV_X1 port map( A => n7556, ZN => n7553);
   U6831 : NAND2_X1 port map( A1 => IF_ISAxsection_0_port, A2 => n5960, ZN => 
                           n5962);
   U6832 : OAI22_X1 port map( A1 => n7452, A2 => n5962, B1 => n5961, B2 => 
                           n7553, ZN => n7555);
   U6833 : INV_X1 port map( A => n7458, ZN => n5964);
   U6834 : OAI22_X1 port map( A1 => n5964, A2 => n7553, B1 => n5963, B2 => 
                           n5962, ZN => n7554);
   U6835 : INV_X1 port map( A => n7253, ZN => n7389);
   U6836 : INV_X1 port map( A => n7073, ZN => n7115);
   U6837 : OAI221_X1 port map( B1 => n7209, B2 => n7389, C1 => n7399, C2 => 
                           n7115, A => n7387, ZN => n5965);
   U6838 : AOI221_X1 port map( B1 => n7410, B2 => n7414, C1 => n7320, C2 => 
                           n7130, A => n5965, ZN => n6025);
   U6839 : INV_X1 port map( A => n7384, ZN => n7276);
   U6840 : OAI22_X1 port map( A1 => n5967, A2 => n7115, B1 => n5966, B2 => 
                           n7316, ZN => n5971);
   U6841 : CLKBUF_X1 port map( A => n5968, Z => n7322);
   U6842 : AOI22_X1 port map( A1 => n7251, A2 => n7130, B1 => n7322, B2 => 
                           n7086, ZN => n5969);
   U6843 : OAI211_X1 port map( C1 => n7118, C2 => n7549, A => n5969, B => n6044
                           , ZN => n5970);
   U6844 : AOI211_X1 port map( C1 => IF_ISAxN2459, C2 => n7276, A => n5971, B 
                           => n5970, ZN => n6024);
   U6845 : NOR2_X1 port map( A1 => intadd_28xBx1x, A2 => ashr_25xAx29x, ZN => 
                           n7257);
   U6846 : AOI22_X1 port map( A1 => n7184, A2 => add_x_26xBx27x, B1 => n7160, 
                           B2 => add_x_26xBx26x, ZN => n6008);
   U6847 : NOR2_X1 port map( A1 => n7080, A2 => ashr_25xAx25x, ZN => n7076);
   U6848 : OAI22_X1 port map( A1 => intadd_26xAx6x, A2 => add_x_26xBx23x, B1 =>
                           intadd_26xAx2x, B2 => add_x_26xBx19x, ZN => n5998);
   U6849 : NOR2_X1 port map( A1 => intadd_26xBx0x, A2 => ashr_25xAx17x, ZN => 
                           n6808);
   U6850 : NOR2_X1 port map( A1 => n6774, A2 => add_x_26xBx16x, ZN => n5993);
   U6851 : NAND2_X1 port map( A1 => n6048, A2 => add_x_26xBx5x, ZN => n5978);
   U6852 : NOR2_X1 port map( A1 => intadd_29xBx2x, A2 => ashr_25xAx3x, ZN => 
                           n6175);
   U6853 : NOR2_X1 port map( A1 => intadd_29xAx2x, A2 => ashr_25xSHx3x, ZN => 
                           n6174);
   U6854 : NOR2_X1 port map( A1 => intadd_29xBx1x, A2 => ashr_25xAx2x, ZN => 
                           n6136);
   U6855 : NAND2_X1 port map( A1 => ashr_25xAx1x, A2 => n7418, ZN => n6070);
   U6856 : AOI22_X1 port map( A1 => n7231, A2 => intadd_29xAx0x, B1 => n6070, 
                           B2 => n5972, ZN => n5973);
   U6857 : INV_X1 port map( A => n5973, ZN => n5974);
   U6858 : OAI22_X1 port map( A1 => n6136, A2 => n5974, B1 => intadd_29xAx1x, 
                           B2 => intadd_25xBx0x, ZN => n5975);
   U6859 : OAI22_X1 port map( A1 => n7331, A2 => ashr_25xAx4x, B1 => n6174, B2 
                           => n5975, ZN => n5976);
   U6860 : OAI22_X1 port map( A1 => n6175, A2 => n5976, B1 => n6251, B2 => 
                           ashr_25xSHx4x, ZN => n5977);
   U6861 : AOI22_X1 port map( A1 => ashr_25xAx5x, A2 => n6283, B1 => n5978, B2 
                           => n5977, ZN => n5979);
   U6862 : NAND2_X1 port map( A1 => ashr_25xAx6x, A2 => n6332, ZN => n6329);
   U6863 : AOI22_X1 port map( A1 => n6330, A2 => add_x_26xBx6x, B1 => n5979, B2
                           => n6329, ZN => n5981);
   U6864 : NAND2_X1 port map( A1 => n6399, A2 => add_x_26xBx7x, ZN => n6406);
   U6865 : OAI22_X1 port map( A1 => n6528, A2 => add_x_26xBx10x, B1 => n6481, 
                           B2 => add_x_26xBx9x, ZN => n5985);
   U6866 : OAI22_X1 port map( A1 => n6399, A2 => add_x_26xBx7x, B1 => n6419, B2
                           => add_x_26xBx8x, ZN => n5980);
   U6867 : AOI211_X1 port map( C1 => n5981, C2 => n6406, A => n5985, B => n5980
                           , ZN => n5991);
   U6868 : OAI22_X1 port map( A1 => n6766, A2 => add_x_26xBx15x, B1 => 
                           intadd_27xAx0x, B2 => add_x_26xBx11x, ZN => n5983);
   U6869 : OAI22_X1 port map( A1 => intadd_27xAx3x, A2 => add_x_26xBx14x, B1 =>
                           intadd_27xAx1x, B2 => add_x_26xBx12x, ZN => n5982);
   U6870 : AOI211_X1 port map( C1 => intadd_27xBx2x, C2 => ashr_25xAx13x, A => 
                           n5983, B => n5982, ZN => n5990);
   U6871 : AOI22_X1 port map( A1 => n6481, A2 => add_x_26xBx9x, B1 => n6419, B2
                           => add_x_26xBx8x, ZN => n5986);
   U6872 : AOI22_X1 port map( A1 => intadd_27xAx0x, A2 => add_x_26xBx11x, B1 =>
                           n6528, B2 => add_x_26xBx10x, ZN => n5984);
   U6873 : OAI21_X1 port map( B1 => n5986, B2 => n5985, A => n5984, ZN => n5989
                           );
   U6874 : NAND2_X1 port map( A1 => n6766, A2 => add_x_26xBx15x, ZN => n5987);
   U6875 : NAND2_X1 port map( A1 => intadd_27xAx3x, A2 => add_x_26xBx14x, ZN =>
                           n6689);
   U6876 : NAND2_X1 port map( A1 => intadd_27xAx2x, A2 => add_x_26xBx13x, ZN =>
                           n6649);
   U6877 : NAND2_X1 port map( A1 => intadd_27xAx1x, A2 => add_x_26xBx12x, ZN =>
                           n6610);
   U6878 : NAND4_X1 port map( A1 => n5987, A2 => n6689, A3 => n6649, A4 => 
                           n6610, ZN => n5988);
   U6879 : AOI221_X1 port map( B1 => n5991, B2 => n5990, C1 => n5989, C2 => 
                           n5990, A => n5988, ZN => n5992);
   U6880 : OAI22_X1 port map( A1 => n6783, A2 => ashr_25xAx16x, B1 => n5993, B2
                           => n5992, ZN => n5996);
   U6881 : AOI22_X1 port map( A1 => intadd_26xBx3x, A2 => ashr_25xAx20x, B1 => 
                           intadd_26xBx1x, B2 => ashr_25xAx18x, ZN => n5995);
   U6882 : AOI22_X1 port map( A1 => intadd_26xBx5x, A2 => ashr_25xAx22x, B1 => 
                           intadd_26xBx4x, B2 => ashr_25xAx21x, ZN => n5994);
   U6883 : OAI211_X1 port map( C1 => n6808, C2 => n5996, A => n5995, B => n5994
                           , ZN => n5997);
   U6884 : AOI211_X1 port map( C1 => intadd_26xBx0x, C2 => ashr_25xAx17x, A => 
                           n5998, B => n5997, ZN => n6001);
   U6885 : NOR2_X1 port map( A1 => intadd_26xBx7x, A2 => ashr_25xAx24x, ZN => 
                           n7051);
   U6886 : NOR2_X1 port map( A1 => intadd_26xBx6x, A2 => ashr_25xAx23x, ZN => 
                           n7006);
   U6887 : NOR2_X1 port map( A1 => intadd_26xBx3x, A2 => ashr_25xAx20x, ZN => 
                           n6918);
   U6888 : NOR2_X1 port map( A1 => intadd_26xBx2x, A2 => ashr_25xAx19x, ZN => 
                           n6885);
   U6889 : AOI211_X1 port map( C1 => intadd_26xAx1x, C2 => add_x_26xBx18x, A =>
                           n6918, B => n6885, ZN => n5999);
   U6890 : NAND2_X1 port map( A1 => intadd_26xAx5x, A2 => add_x_26xBx22x, ZN =>
                           n6975);
   U6891 : OAI211_X1 port map( C1 => intadd_26xBx4x, C2 => ashr_25xAx21x, A => 
                           n5999, B => n6975, ZN => n6000);
   U6892 : NOR4_X1 port map( A1 => n6001, A2 => n7051, A3 => n7006, A4 => n6000
                           , ZN => n6003);
   U6893 : AOI211_X1 port map( C1 => intadd_26xBx7x, C2 => ashr_25xAx24x, A => 
                           n6003, B => n6002, ZN => n6004);
   U6894 : OAI22_X1 port map( A1 => n7076, A2 => n6004, B1 => n7160, B2 => 
                           add_x_26xBx26x, ZN => n6007);
   U6895 : NOR2_X1 port map( A1 => n7184, A2 => add_x_26xBx27x, ZN => n6006);
   U6896 : OAI22_X1 port map( A1 => intadd_28xAx1x, A2 => add_x_26xBx29x, B1 =>
                           intadd_28xAx0x, B2 => add_x_26xBx28x, ZN => n6005);
   U6897 : AOI211_X1 port map( C1 => n6008, C2 => n6007, A => n6006, B => n6005
                           , ZN => n6009);
   U6898 : AOI211_X1 port map( C1 => intadd_28xAx0x, C2 => add_x_26xBx28x, A =>
                           n7257, B => n6009, ZN => n6010);
   U6899 : NAND2_X1 port map( A1 => intadd_28xAx2x, A2 => add_x_26xBx30x, ZN =>
                           n7317);
   U6900 : AOI22_X1 port map( A1 => n6010, A2 => n7317, B1 => intadd_28xBx2x, 
                           B2 => ashr_25xAx30x, ZN => n6014);
   U6901 : NAND2_X1 port map( A1 => n7413, A2 => n7392, ZN => n6011);
   U6902 : INV_X1 port map( A => n6013, ZN => n7411);
   U6903 : AOI21_X1 port map( B1 => n6014, B2 => n6011, A => n7411, ZN => n6018
                           );
   U6904 : INV_X1 port map( A => n6011, ZN => n6012);
   U6905 : AOI21_X1 port map( B1 => n6014, B2 => n6013, A => n6012, ZN => n6016
                           );
   U6906 : OAI22_X1 port map( A1 => n6018, A2 => n6017, B1 => n6016, B2 => 
                           n6015, ZN => n6021);
   U6907 : AOI22_X1 port map( A1 => n6022, A2 => n6021, B1 => n6020, B2 => 
                           n6019, ZN => n6023);
   U6908 : OAI211_X1 port map( C1 => n6026, C2 => n6025, A => n6024, B => n6023
                           , ZN => n6043);
   U6909 : CLKBUF_X1 port map( A => n7159, Z => n7368);
   U6910 : NAND2_X1 port map( A1 => n7376, A2 => n6900, ZN => n7406);
   U6911 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx4x, B1 => 
                           ashr_25xAx5x, B2 => n7086, ZN => n6122);
   U6912 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx6x, B1 => 
                           ashr_25xAx7x, B2 => n7399, ZN => n6117);
   U6913 : AOI22_X1 port map( A1 => n7304, A2 => n6122, B1 => n6117, B2 => 
                           n7402, ZN => n6229);
   U6914 : NOR2_X1 port map( A1 => intadd_29xAx0x, A2 => n7209, ZN => n6148);
   U6915 : AOI22_X1 port map( A1 => n7209, A2 => intadd_29xAx1x, B1 => 
                           intadd_29xAx2x, B2 => n7399, ZN => n6124);
   U6916 : NAND3_X1 port map( A1 => n7304, A2 => n7209, A3 => ashr_25xAx0x, ZN 
                           => n6430);
   U6917 : INV_X1 port map( A => n6430, ZN => n6245);
   U6918 : AOI221_X1 port map( B1 => n6148, B2 => n7304, C1 => n6124, C2 => 
                           n5711, A => n6245, ZN => n6027);
   U6919 : INV_X1 port map( A => n6110, ZN => n7311);
   U6920 : NAND2_X1 port map( A1 => n7311, A2 => n7376, ZN => n7269);
   U6921 : INV_X1 port map( A => n7269, ZN => n7400);
   U6922 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx8x, B1 => 
                           ashr_25xAx9x, B2 => n7086, ZN => n6116);
   U6923 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx10x, B1 => 
                           ashr_25xAx11x, B2 => n7267, ZN => n6119);
   U6924 : AOI22_X1 port map( A1 => n7304, A2 => n6116, B1 => n6119, B2 => 
                           n5711, ZN => n6230);
   U6925 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx12x, B1 => 
                           ashr_25xAx13x, B2 => n7267, ZN => n6118);
   U6926 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx14x, B1 => 
                           ashr_25xAx15x, B2 => n7267, ZN => n6121);
   U6927 : AOI22_X1 port map( A1 => n7304, A2 => n6118, B1 => n6121, B2 => 
                           n7402, ZN => n6228);
   U6928 : AOI22_X1 port map( A1 => n7311, A2 => n6230, B1 => n6228, B2 => 
                           n6900, ZN => n6411);
   U6929 : AOI22_X1 port map( A1 => n6027, A2 => n7400, B1 => n7207, B2 => 
                           n6411, ZN => n6028);
   U6930 : AND2_X1 port map( A1 => n6325, A2 => n7192, ZN => n6653);
   U6931 : INV_X1 port map( A => n6653, ZN => n6494);
   U6932 : NAND2_X1 port map( A1 => n7427, A2 => n6494, ZN => n6683);
   U6933 : OAI211_X1 port map( C1 => n7406, C2 => n6229, A => n6028, B => n6683
                           , ZN => n6039);
   U6934 : NAND2_X1 port map( A1 => intadd_29xBx2x, A2 => intadd_29xBx1x, ZN =>
                           n7415);
   U6935 : NOR3_X1 port map( A1 => n7231, A2 => n6250, A3 => n7415, ZN => n6788
                           );
   U6936 : NOR2_X1 port map( A1 => n7269, A2 => n6430, ZN => n6787);
   U6937 : AOI22_X1 port map( A1 => n7420, A2 => n6788, B1 => n7409, B2 => 
                           n6787, ZN => n6038);
   U6938 : INV_X1 port map( A => n6346, ZN => n6387);
   U6939 : NOR2_X1 port map( A1 => n7192, A2 => n6387, ZN => n6715);
   U6940 : AND2_X1 port map( A1 => n6325, A2 => n7349, ZN => n6678);
   U6941 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx16x, B1 => 
                           ashr_25xAx17x, B2 => n7267, ZN => n6120);
   U6942 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx18x, B1 => 
                           ashr_25xAx19x, B2 => n7086, ZN => n6113);
   U6943 : AOI22_X1 port map( A1 => n7304, A2 => n6120, B1 => n6113, B2 => 
                           n7402, ZN => n6227);
   U6944 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx20x, B1 => 
                           ashr_25xAx21x, B2 => n7267, ZN => n6112);
   U6945 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx22x, B1 => 
                           ashr_25xAx23x, B2 => n7086, ZN => n6115);
   U6946 : AOI22_X1 port map( A1 => n7304, A2 => n6112, B1 => n6115, B2 => 
                           n5711, ZN => n6237);
   U6947 : AOI22_X1 port map( A1 => n7311, A2 => n6227, B1 => n6237, B2 => 
                           n6900, ZN => n6410);
   U6948 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx24x, B1 => 
                           ashr_25xAx25x, B2 => n7267, ZN => n6114);
   U6949 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx26x, B1 => 
                           ashr_25xAx27x, B2 => n7086, ZN => n6109);
   U6950 : AOI22_X1 port map( A1 => n7304, A2 => n6114, B1 => n6109, B2 => 
                           n7402, ZN => n6238);
   U6951 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx28x, B1 => 
                           ashr_25xAx29x, B2 => n7267, ZN => n6108);
   U6952 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx30x, B1 => n7413, B2
                           => n7267, ZN => n6111);
   U6953 : AOI22_X1 port map( A1 => n7304, A2 => n6108, B1 => n6111, B2 => 
                           n5711, ZN => n6592);
   U6954 : AOI22_X1 port map( A1 => n7311, A2 => n6238, B1 => n6592, B2 => 
                           n7309, ZN => n7049);
   U6955 : AOI22_X1 port map( A1 => n7376, A2 => n6410, B1 => n7049, B2 => 
                           n7207, ZN => n6786);
   U6956 : OAI21_X1 port map( B1 => n6715, B2 => n6678, A => n6786, ZN => n6037
                           );
   U6957 : AOI22_X1 port map( A1 => n7414, A2 => intadd_26xAx7x, B1 => n7129, 
                           B2 => n7130, ZN => n6129);
   U6958 : AOI22_X1 port map( A1 => n7414, A2 => n7160, B1 => n7184, B2 => 
                           n7130, ZN => n6338);
   U6959 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6129, B1 => n6338, 
                           B2 => n7259, ZN => n6252);
   U6960 : AOI22_X1 port map( A1 => n7414, A2 => intadd_28xAx0x, B1 => 
                           intadd_28xAx1x, B2 => n7130, ZN => n6337);
   U6961 : AOI22_X1 port map( A1 => n7414, A2 => intadd_28xAx2x, B1 => n7435, 
                           B2 => n7130, ZN => n6131);
   U6962 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6337, B1 => n6131, 
                           B2 => n7259, ZN => n7245);
   U6963 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6252, B1 => n7245, 
                           B2 => n6456, ZN => n7042);
   U6964 : NAND2_X1 port map( A1 => n7042, A2 => ashr_25xSHx3x, ZN => n6030);
   U6965 : AOI22_X1 port map( A1 => n7414, A2 => n6774, B1 => intadd_26xAx0x, 
                           B2 => n7130, ZN => n6100);
   U6966 : AOI22_X1 port map( A1 => n7414, A2 => intadd_26xAx1x, B1 => 
                           intadd_26xAx2x, B2 => n7130, ZN => n6128);
   U6967 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6100, B1 => n6128, 
                           B2 => n7231, ZN => n6232);
   U6968 : AOI22_X1 port map( A1 => n7414, A2 => intadd_26xAx3x, B1 => 
                           intadd_26xAx4x, B2 => n7130, ZN => n6127);
   U6969 : AOI22_X1 port map( A1 => n7414, A2 => intadd_26xAx5x, B1 => 
                           intadd_26xAx6x, B2 => n7130, ZN => n6130);
   U6970 : AOI22_X1 port map( A1 => n7418, A2 => n6127, B1 => n6130, B2 => 
                           n7231, ZN => n6253);
   U6971 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6232, B1 => n6253, 
                           B2 => n6456, ZN => n6423);
   U6972 : NAND2_X1 port map( A1 => n6423, A2 => intadd_29xBx2x, ZN => n6029);
   U6973 : AND2_X1 port map( A1 => n6030, A2 => n6029, ZN => n6789);
   U6974 : INV_X1 port map( A => n6789, ZN => n6035);
   U6975 : NAND2_X1 port map( A1 => n6072, A2 => n6047, ZN => n6058);
   U6976 : INV_X1 port map( A => n7415, ZN => n7341);
   U6977 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx2x, B1 => 
                           ashr_25xAx3x, B2 => n7130, ZN => n6102);
   U6978 : OAI22_X1 port map( A1 => n7414, A2 => n6070, B1 => n7418, B2 => 
                           n6102, ZN => n6031);
   U6979 : AOI22_X1 port map( A1 => n7414, A2 => n6419, B1 => n6481, B2 => 
                           n7412, ZN => n6096);
   U6980 : AOI22_X1 port map( A1 => n7414, A2 => n6528, B1 => intadd_27xAx0x, 
                           B2 => n7412, ZN => n6099);
   U6981 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6096, B1 => n6099, 
                           B2 => n7231, ZN => n6236);
   U6982 : AOI22_X1 port map( A1 => n7414, A2 => intadd_27xAx1x, B1 => 
                           intadd_27xAx2x, B2 => n7130, ZN => n6098);
   U6983 : AOI22_X1 port map( A1 => n7414, A2 => intadd_27xAx3x, B1 => n6766, 
                           B2 => n7130, ZN => n6101);
   U6984 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6098, B1 => n6101, 
                           B2 => n7259, ZN => n6233);
   U6985 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6236, B1 => n6233, 
                           B2 => n6456, ZN => n6422);
   U6986 : AOI22_X1 port map( A1 => n7341, A2 => n6031, B1 => n6422, B2 => 
                           ashr_25xSHx3x, ZN => n6033);
   U6987 : NOR2_X1 port map( A1 => intadd_29xBx1x, A2 => ashr_25xSHx3x, ZN => 
                           n7422);
   U6988 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx4x, B1 => 
                           ashr_25xAx5x, B2 => n7130, ZN => n6103);
   U6989 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx6x, B1 => 
                           ashr_25xAx7x, B2 => n7130, ZN => n6095);
   U6990 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6103, B1 => n6095, 
                           B2 => n7416, ZN => n6234);
   U6991 : AOI211_X1 port map( C1 => n7422, C2 => n6234, A => n6788, B => 
                           ashr_25xSHx4x, ZN => n6032);
   U6992 : NAND2_X1 port map( A1 => n6033, A2 => n6032, ZN => n6034);
   U6993 : OAI211_X1 port map( C1 => n6035, C2 => n7331, A => n6058, B => n6034
                           , ZN => n6036);
   U6994 : NAND4_X1 port map( A1 => n6039, A2 => n6038, A3 => n6037, A4 => 
                           n6036, ZN => n6040);
   U6995 : AOI21_X1 port map( B1 => DP_OP_719J14_125_1055xn69, B2 => n7368, A 
                           => n6040, ZN => n6041);
   U6996 : INV_X1 port map( A => n6041, ZN => n6042);
   U6997 : OAI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(0), A2 => n6044,
                           B1 => n6043, B2 => n6042, ZN => n6045);
   U6998 : NOR2_X1 port map( A1 => rst, A2 => n6045, ZN => IF_ISAxN10936);
   U6999 : OAI22_X1 port map( A1 => n7404, A2 => n7389, B1 => n7418, B2 => 
                           n7386, ZN => n6084);
   U7000 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6074, B1 => n6046, 
                           B2 => n6456, ZN => n6461);
   U7001 : AOI22_X1 port map( A1 => n7414, A2 => intadd_26xAx0x, B1 => 
                           intadd_26xAx1x, B2 => n7412, ZN => n6167);
   U7002 : AOI22_X1 port map( A1 => n7414, A2 => intadd_26xAx2x, B1 => 
                           intadd_26xAx3x, B2 => n7412, ZN => n6204);
   U7003 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6167, B1 => n6204, 
                           B2 => n7231, ZN => n6483);
   U7004 : OAI221_X1 port map( B1 => intadd_29xBx1x, B2 => n6482, C1 => 
                           intadd_25xBx0x, C2 => n6483, A => n7236, ZN => n6075
                           );
   U7005 : OAI21_X1 port map( B1 => n6461, B2 => intadd_29xBx2x, A => n6075, ZN
                           => n6827);
   U7006 : INV_X1 port map( A => n6827, ZN => n6055);
   U7007 : NOR2_X1 port map( A1 => n6047, A2 => n7331, ZN => n6734);
   U7008 : AOI22_X1 port map( A1 => n7209, A2 => n6048, B1 => n6330, B2 => 
                           n7086, ZN => n6184);
   U7009 : AOI22_X1 port map( A1 => n7209, A2 => n6399, B1 => n6419, B2 => 
                           n7267, ZN => n6179);
   U7010 : AOI22_X1 port map( A1 => n7304, A2 => n6184, B1 => n6179, B2 => 
                           n5711, ZN => n6286);
   U7011 : INV_X1 port map( A => n7406, ZN => n7275);
   U7012 : AOI22_X1 port map( A1 => n7209, A2 => n6481, B1 => n6528, B2 => 
                           n7086, ZN => n6178);
   U7013 : AOI22_X1 port map( A1 => n7209, A2 => intadd_27xAx0x, B1 => 
                           intadd_27xAx1x, B2 => n7086, ZN => n6181);
   U7014 : AOI22_X1 port map( A1 => n7304, A2 => n6178, B1 => n6181, B2 => 
                           n5711, ZN => n6287);
   U7015 : AOI22_X1 port map( A1 => n7209, A2 => intadd_27xAx2x, B1 => 
                           intadd_27xAx3x, B2 => n7086, ZN => n6180);
   U7016 : AOI22_X1 port map( A1 => n7209, A2 => n6766, B1 => n6774, B2 => 
                           n7086, ZN => n6183);
   U7017 : AOI22_X1 port map( A1 => n7304, A2 => n6180, B1 => n6183, B2 => 
                           n5711, ZN => n6285);
   U7018 : AOI22_X1 port map( A1 => n7311, A2 => n6287, B1 => n6285, B2 => 
                           n7309, ZN => n6455);
   U7019 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx3x, B1 => 
                           ashr_25xAx4x, B2 => n7399, ZN => n6185);
   U7020 : INV_X1 port map( A => n6185, ZN => n6052);
   U7021 : NOR2_X1 port map( A1 => ashr_25xAx1x, A2 => n7086, ZN => n6050);
   U7022 : NOR2_X1 port map( A1 => n7209, A2 => ashr_25xAx2x, ZN => n6049);
   U7023 : NOR2_X1 port map( A1 => n6050, A2 => n6049, ZN => n6051);
   U7024 : MUX2_X1 port map( A => n6052, B => n6051, S => n7304, Z => n6053);
   U7025 : OAI22_X1 port map( A1 => n7376, A2 => n6455, B1 => n6053, B2 => 
                           n7269, ZN => n6054);
   U7026 : AOI211_X1 port map( C1 => n6286, C2 => n7275, A => n7349, B => n6054
                           , ZN => n6087);
   U7027 : AOI222_X1 port map( A1 => DP_OP_719J14_125_1055xn70, A2 => n7368, B1
                           => n6055, B2 => n6734, C1 => n6325, C2 => n6087, ZN 
                           => n6056);
   U7028 : INV_X1 port map( A => n6056, ZN => n6083);
   U7029 : AOI22_X1 port map( A1 => n7414, A2 => intadd_29xAx0x, B1 => 
                           intadd_29xAx1x, B2 => n7412, ZN => n6057);
   U7030 : AOI22_X1 port map( A1 => n7414, A2 => intadd_29xAx2x, B1 => n6251, 
                           B2 => n7412, ZN => n6164);
   U7031 : AOI221_X1 port map( B1 => n6057, B2 => n7418, C1 => n6164, C2 => 
                           n7259, A => n7415, ZN => n6061);
   U7032 : NAND2_X1 port map( A1 => n7331, A2 => n6058, ZN => n6720);
   U7033 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx9x, B1 => 
                           ashr_25xAx10x, B2 => n7412, ZN => n6169);
   U7034 : INV_X1 port map( A => n6169, ZN => n6059);
   U7035 : AOI22_X1 port map( A1 => n7414, A2 => intadd_27xAx0x, B1 => 
                           intadd_27xAx1x, B2 => n7412, ZN => n6166);
   U7036 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6059, B1 => n6166, 
                           B2 => n7416, ZN => n6277);
   U7037 : AOI22_X1 port map( A1 => n7414, A2 => intadd_27xAx2x, B1 => 
                           intadd_27xAx3x, B2 => n7412, ZN => n6165);
   U7038 : AOI22_X1 port map( A1 => n7414, A2 => n6766, B1 => n6774, B2 => 
                           n7412, ZN => n6168);
   U7039 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6165, B1 => n6168, 
                           B2 => n7231, ZN => n6274);
   U7040 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6277, B1 => n6274, 
                           B2 => n6456, ZN => n6484);
   U7041 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx5x, B1 => 
                           ashr_25xAx6x, B2 => n7412, ZN => n6162);
   U7042 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx7x, B1 => 
                           ashr_25xAx8x, B2 => n7412, ZN => n6170);
   U7043 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6162, B1 => n6170, 
                           B2 => n7416, ZN => n6275);
   U7044 : INV_X1 port map( A => n7422, ZN => n7132);
   U7045 : OAI22_X1 port map( A1 => n7236, A2 => n6484, B1 => n6275, B2 => 
                           n7132, ZN => n6060);
   U7046 : NOR3_X1 port map( A1 => n6061, A2 => n6720, A3 => n6060, ZN => n6063
                           );
   U7047 : OAI22_X1 port map( A1 => n7418, A2 => n7387, B1 => n7118, B2 => 
                           n7542, ZN => n6062);
   U7048 : AOI211_X1 port map( C1 => n7327, C2 => n6064, A => n6063, B => n6062
                           , ZN => n6081);
   U7049 : NAND2_X1 port map( A1 => n7311, A2 => n6065, ZN => n6085);
   U7050 : OAI21_X1 port map( B1 => n7311, B2 => n6651, A => n6085, ZN => n6469
                           );
   U7051 : AOI22_X1 port map( A1 => n7209, A2 => intadd_26xAx0x, B1 => 
                           intadd_26xAx1x, B2 => n7267, ZN => n6182);
   U7052 : AOI22_X1 port map( A1 => n7209, A2 => intadd_26xAx2x, B1 => 
                           intadd_26xAx3x, B2 => n7086, ZN => n6197);
   U7053 : AOI22_X1 port map( A1 => n7304, A2 => n6182, B1 => n6197, B2 => 
                           n5711, ZN => n6284);
   U7054 : AOI22_X1 port map( A1 => n7311, A2 => n6284, B1 => n6066, B2 => 
                           n6900, ZN => n6454);
   U7055 : NOR2_X1 port map( A1 => n6454, A2 => n7207, ZN => n6086);
   U7056 : AOI21_X1 port map( B1 => n7207, B2 => n6469, A => n6086, ZN => n6815
                           );
   U7057 : NAND2_X1 port map( A1 => intadd_29xAx0x, A2 => n7231, ZN => n6071);
   U7058 : AOI22_X1 port map( A1 => n6068, A2 => n7276, B1 => n6067, B2 => 
                           n7327, ZN => n6069);
   U7059 : OAI221_X1 port map( B1 => n7316, B2 => n6071, C1 => n7255, C2 => 
                           n6070, A => n6069, ZN => n6079);
   U7060 : INV_X1 port map( A => n6072, ZN => n6073);
   U7061 : AND2_X1 port map( A1 => ashr_25xSHx4x, A2 => n6073, ZN => n6598);
   U7062 : INV_X1 port map( A => n6598, ZN => n6463);
   U7063 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6074, B1 => n7286, 
                           B2 => n6456, ZN => n6462);
   U7064 : OAI21_X1 port map( B1 => n7236, B2 => n6462, A => n6075, ZN => n6819
                           );
   U7065 : NOR2_X1 port map( A1 => n7415, A2 => n6459, ZN => n6828);
   U7066 : NAND2_X1 port map( A1 => n7400, A2 => n6467, ZN => n6820);
   U7067 : INV_X1 port map( A => n6820, ZN => n6076);
   U7068 : AOI22_X1 port map( A1 => n7420, A2 => n6828, B1 => n7409, B2 => 
                           n6076, ZN => n6077);
   U7069 : OAI21_X1 port map( B1 => n6463, B2 => n6819, A => n6077, ZN => n6078
                           );
   U7070 : AOI211_X1 port map( C1 => n6678, C2 => n6815, A => n6079, B => n6078
                           , ZN => n6080);
   U7071 : OAI211_X1 port map( C1 => n7304, C2 => n7398, A => n6081, B => n6080
                           , ZN => n6082);
   U7072 : AOI211_X1 port map( C1 => ashr_25xAx1x, C2 => n6084, A => n6083, B 
                           => n6082, ZN => n6090);
   U7073 : NOR2_X1 port map( A1 => n7387, A2 => n7533, ZN => n6547);
   U7074 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(1), A2 => n6597,
                           B1 => n6547, B2 => ashr_25xAx1x, ZN => n6089);
   U7075 : NAND2_X1 port map( A1 => n6715, A2 => n7029, ZN => n6632);
   U7076 : INV_X1 port map( A => n6632, ZN => n6453);
   U7077 : OAI21_X1 port map( B1 => n7311, B2 => n6645, A => n6085, ZN => n7083
                           );
   U7078 : AOI21_X1 port map( B1 => n7207, B2 => n7083, A => n6086, ZN => n6829
                           );
   U7079 : NOR2_X1 port map( A1 => n6387, A2 => n7533, ZN => n6305);
   U7080 : AOI22_X1 port map( A1 => n6453, A2 => n6829, B1 => n6305, B2 => 
                           n6087, ZN => n6088);
   U7081 : OAI211_X1 port map( C1 => n6090, C2 => n7533, A => n6089, B => n6088
                           , ZN => IF_ISAxN10938);
   U7082 : INV_X1 port map( A => n7118, ZN => n7447);
   U7083 : AOI22_X1 port map( A1 => n7251, A2 => n6811, B1 => n7447, B2 => 
                           n7546, ZN => n6093);
   U7084 : OAI22_X1 port map( A1 => intadd_29xBx1x, A2 => n7386, B1 => n7311, 
                           B2 => n7389, ZN => n6091);
   U7085 : OAI21_X1 port map( B1 => n7251, B2 => n6091, A => ashr_25xAx2x, ZN 
                           => n6092);
   U7086 : OAI211_X1 port map( C1 => n7384, C2 => n6094, A => n6093, B => n6092
                           , ZN => n6156);
   U7087 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn71, A2 => n7368, ZN 
                           => n6154);
   U7088 : INV_X1 port map( A => n6095, ZN => n6097);
   U7089 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6097, B1 => n6096, 
                           B2 => n7259, ZN => n6314);
   U7090 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6099, B1 => n6098, 
                           B2 => n7416, ZN => n6313);
   U7091 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6101, B1 => n6100, 
                           B2 => n7231, ZN => n6312);
   U7092 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6313, B1 => n6312, 
                           B2 => n6456, ZN => n6508);
   U7093 : OAI221_X1 port map( B1 => n7418, B2 => n6103, C1 => n7231, C2 => 
                           n6102, A => n7341, ZN => n6104);
   U7094 : OAI21_X1 port map( B1 => n7236, B2 => n6508, A => n6104, ZN => n6105
                           );
   U7095 : AOI211_X1 port map( C1 => n7422, C2 => n6314, A => n6720, B => n6105
                           , ZN => n6143);
   U7096 : NAND2_X1 port map( A1 => n7311, A2 => ashr_25xAx2x, ZN => n6107);
   U7097 : AOI21_X1 port map( B1 => n6107, B2 => n6106, A => n7397, ZN => n6142
                           );
   U7098 : AOI22_X1 port map( A1 => n7404, A2 => n6109, B1 => n6108, B2 => 
                           n7402, ZN => n6681);
   U7099 : NOR2_X1 port map( A1 => n6110, A2 => n6681, ZN => n6145);
   U7100 : NOR2_X1 port map( A1 => n5711, A2 => n6111, ZN => n6672);
   U7101 : NOR2_X1 port map( A1 => n6941, A2 => n6672, ZN => n6146);
   U7102 : NOR2_X1 port map( A1 => n6145, A2 => n6146, ZN => n6500);
   U7103 : AOI22_X1 port map( A1 => n7404, A2 => n6113, B1 => n6112, B2 => 
                           n7402, ZN => n6319);
   U7104 : AOI22_X1 port map( A1 => n7404, A2 => n6115, B1 => n6114, B2 => 
                           n7402, ZN => n6682);
   U7105 : AOI22_X1 port map( A1 => n6941, A2 => n6319, B1 => n6682, B2 => 
                           n6900, ZN => n6525);
   U7106 : NOR2_X1 port map( A1 => n6525, A2 => n7207, ZN => n6147);
   U7107 : AOI21_X1 port map( B1 => n6500, B2 => n7207, A => n6147, ZN => n6858
                           );
   U7108 : INV_X1 port map( A => n6715, ZN => n6729);
   U7109 : AOI22_X1 port map( A1 => n7304, A2 => n6117, B1 => n6116, B2 => 
                           n5711, ZN => n6321);
   U7110 : AOI22_X1 port map( A1 => n7304, A2 => n6119, B1 => n6118, B2 => 
                           n7402, ZN => n6322);
   U7111 : AOI22_X1 port map( A1 => n7304, A2 => n6121, B1 => n6120, B2 => 
                           n7402, ZN => n6320);
   U7112 : AOI22_X1 port map( A1 => n6941, A2 => n6322, B1 => n6320, B2 => 
                           n6900, ZN => n6523);
   U7113 : INV_X1 port map( A => n6122, ZN => n6123);
   U7114 : AOI221_X1 port map( B1 => n6124, B2 => n7304, C1 => n6123, C2 => 
                           n5711, A => n7269, ZN => n6125);
   U7115 : AOI211_X1 port map( C1 => n7207, C2 => n6523, A => n6125, B => n7349
                           , ZN => n6126);
   U7116 : OAI21_X1 port map( B1 => n7406, B2 => n6321, A => n6126, ZN => n6144
                           );
   U7117 : OAI22_X1 port map( A1 => n6858, A2 => n6729, B1 => n6386, B2 => 
                           n6144, ZN => n6141);
   U7118 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx2x, B1 => 
                           ashr_25xAx1x, B2 => n7412, ZN => n6249);
   U7119 : AOI22_X1 port map( A1 => intadd_29xBx0x, A2 => n6249, B1 => n6250, 
                           B2 => n7259, ZN => n6502);
   U7120 : NAND2_X1 port map( A1 => n7341, A2 => n6502, ZN => n6857);
   U7121 : AOI22_X1 port map( A1 => n7418, A2 => n6128, B1 => n6127, B2 => 
                           n7231, ZN => n6311);
   U7122 : AOI22_X1 port map( A1 => n7418, A2 => n6130, B1 => n6129, B2 => 
                           n7231, ZN => n6340);
   U7123 : AOI22_X1 port map( A1 => n6962, A2 => n6311, B1 => n6340, B2 => 
                           n6456, ZN => n6509);
   U7124 : NOR2_X1 port map( A1 => n6509, A2 => ashr_25xSHx3x, ZN => n6134);
   U7125 : NAND2_X1 port map( A1 => n7418, A2 => n6131, ZN => n6711);
   U7126 : AOI221_X1 port map( B1 => n6338, B2 => n7418, C1 => n6337, C2 => 
                           n7416, A => n6811, ZN => n6132);
   U7127 : AOI21_X1 port map( B1 => n6456, B2 => n6711, A => n6132, ZN => n6517
                           );
   U7128 : NOR2_X1 port map( A1 => intadd_29xBx2x, A2 => n6517, ZN => n6135);
   U7129 : NOR2_X1 port map( A1 => n6134, A2 => n6135, ZN => n6843);
   U7130 : INV_X1 port map( A => n6132, ZN => n6133);
   U7131 : NAND2_X1 port map( A1 => n6343, A2 => n6133, ZN => n6526);
   U7132 : AOI21_X1 port map( B1 => n6135, B2 => n6526, A => n6134, ZN => n6863
                           );
   U7133 : OAI221_X1 port map( B1 => n6734, B2 => n6843, C1 => n6734, C2 => 
                           n6598, A => n6863, ZN => n6139);
   U7134 : NOR2_X1 port map( A1 => intadd_29xAx1x, A2 => intadd_25xBx0x, ZN => 
                           n6137);
   U7135 : OAI21_X1 port map( B1 => n6137, B2 => n6136, A => n7127, ZN => n6138
                           );
   U7136 : OAI211_X1 port map( C1 => n7343, C2 => n6857, A => n6139, B => n6138
                           , ZN => n6140);
   U7137 : NOR4_X1 port map( A1 => n6143, A2 => n6142, A3 => n6141, A4 => n6140
                           , ZN => n6153);
   U7138 : INV_X1 port map( A => n6144, ZN => n6151);
   U7139 : AOI21_X1 port map( B1 => n6146, B2 => n6676, A => n6145, ZN => n6519
                           );
   U7140 : AOI21_X1 port map( B1 => n6519, B2 => n7207, A => n6147, ZN => n6841
                           );
   U7141 : INV_X1 port map( A => n6678, ZN => n6580);
   U7142 : INV_X1 port map( A => n7409, ZN => n7206);
   U7143 : AOI21_X1 port map( B1 => n7209, B2 => ashr_25xAx2x, A => n6148, ZN 
                           => n6244);
   U7144 : NAND2_X1 port map( A1 => n7209, A2 => ashr_25xAx0x, ZN => n6149);
   U7145 : AOI22_X1 port map( A1 => n7404, A2 => n6244, B1 => n6149, B2 => 
                           n7402, ZN => n6513);
   U7146 : NAND2_X1 port map( A1 => n7400, A2 => n6513, ZN => n6845);
   U7147 : OAI22_X1 port map( A1 => n6841, A2 => n6580, B1 => n7206, B2 => 
                           n6845, ZN => n6150);
   U7148 : AOI21_X1 port map( B1 => n6346, B2 => n6151, A => n6150, ZN => n6152
                           );
   U7149 : NAND3_X1 port map( A1 => n6154, A2 => n6153, A3 => n6152, ZN => 
                           n6155);
   U7150 : AOI211_X1 port map( C1 => n7322, C2 => n7309, A => n6156, B => n6155
                           , ZN => n6158);
   U7151 : OAI22_X1 port map( A1 => n6158, A2 => n6717, B1 => n6157, B2 => 
                           n7439, ZN => IF_ISAxN10939);
   U7152 : NOR2_X1 port map( A1 => intadd_29xAx2x, A2 => n7207, ZN => n6218);
   U7153 : AOI22_X1 port map( A1 => n7418, A2 => n6160, B1 => n6159, B2 => 
                           n7231, ZN => n6563);
   U7154 : OR2_X1 port map( A1 => n7415, A2 => n6563, ZN => n6906);
   U7155 : OAI22_X1 port map( A1 => n6161, A2 => n7115, B1 => n7343, B2 => 
                           n6906, ZN => n6217);
   U7156 : INV_X1 port map( A => n6162, ZN => n6163);
   U7157 : AOI221_X1 port map( B1 => n6164, B2 => intadd_29xBx0x, C1 => n6163, 
                           C2 => n7259, A => n7415, ZN => n6172);
   U7158 : AOI22_X1 port map( A1 => n7418, A2 => n6166, B1 => n6165, B2 => 
                           n7416, ZN => n6372);
   U7159 : AOI22_X1 port map( A1 => n7418, A2 => n6168, B1 => n6167, B2 => 
                           n7231, ZN => n6369);
   U7160 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6372, B1 => n6369, 
                           B2 => n6456, ZN => n6551);
   U7161 : AOI22_X1 port map( A1 => n7418, A2 => n6170, B1 => n6169, B2 => 
                           n7259, ZN => n6370);
   U7162 : OAI22_X1 port map( A1 => n7236, A2 => n6551, B1 => n6370, B2 => 
                           n7132, ZN => n6171);
   U7163 : NOR3_X1 port map( A1 => n6172, A2 => n6720, A3 => n6171, ZN => n6173
                           );
   U7164 : AOI221_X1 port map( B1 => n6175, B2 => n7410, C1 => n6174, C2 => 
                           n7410, A => n6173, ZN => n6214);
   U7165 : OAI22_X1 port map( A1 => intadd_29xBx2x, A2 => n7386, B1 => n7376, 
                           B2 => n7389, ZN => n6212);
   U7166 : AOI22_X1 port map( A1 => n7404, A2 => n6177, B1 => n6176, B2 => 
                           n7402, ZN => n6564);
   U7167 : NAND2_X1 port map( A1 => n7400, A2 => n6564, ZN => n6884);
   U7168 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn72, A2 => n7159, ZN 
                           => n6193);
   U7169 : AOI22_X1 port map( A1 => n7404, A2 => n6179, B1 => n6178, B2 => 
                           n7402, ZN => n6382);
   U7170 : AOI22_X1 port map( A1 => n7404, A2 => n6181, B1 => n6180, B2 => 
                           n7402, ZN => n6383);
   U7171 : AOI22_X1 port map( A1 => n7404, A2 => n6183, B1 => n6182, B2 => 
                           n7402, ZN => n6381);
   U7172 : AOI22_X1 port map( A1 => n7311, A2 => n6383, B1 => n6381, B2 => 
                           n6900, ZN => n6575);
   U7173 : INV_X1 port map( A => n6184, ZN => n6186);
   U7174 : OAI221_X1 port map( B1 => n7404, B2 => n6186, C1 => n7402, C2 => 
                           n6185, A => n7400, ZN => n6187);
   U7175 : OAI211_X1 port map( C1 => n7376, C2 => n6575, A => n7192, B => n6187
                           , ZN => n6188);
   U7176 : AOI21_X1 port map( B1 => n7275, B2 => n6382, A => n6188, ZN => n6223
                           );
   U7177 : OAI22_X1 port map( A1 => n7376, A2 => n7398, B1 => n7118, B2 => 
                           n6189, ZN => n6191);
   U7178 : NOR2_X1 port map( A1 => n7387, A2 => intadd_29xBx2x, ZN => n6190);
   U7179 : AOI211_X1 port map( C1 => n6325, C2 => n6223, A => n6191, B => n6190
                           , ZN => n6192);
   U7180 : OAI211_X1 port map( C1 => n6884, C2 => n7206, A => n6193, B => n6192
                           , ZN => n6211);
   U7181 : AOI22_X1 port map( A1 => n7404, A2 => n6195, B1 => n6194, B2 => 
                           n7402, ZN => n6574);
   U7182 : AOI21_X1 port map( B1 => n7311, B2 => n6574, A => n7376, ZN => n6222
                           );
   U7183 : AOI22_X1 port map( A1 => n7404, A2 => n6197, B1 => n6196, B2 => 
                           n7402, ZN => n6380);
   U7184 : OAI22_X1 port map( A1 => n7402, A2 => n6199, B1 => n6198, B2 => 
                           n7304, ZN => n6363);
   U7185 : AOI22_X1 port map( A1 => n6941, A2 => n6380, B1 => n6363, B2 => 
                           n7309, ZN => n6576);
   U7186 : NOR2_X1 port map( A1 => n6576, A2 => n7207, ZN => n6220);
   U7187 : AOI221_X1 port map( B1 => n6222, B2 => n7435, C1 => n6222, C2 => 
                           n7311, A => n6220, ZN => n6200);
   U7188 : INV_X1 port map( A => n6200, ZN => n6897);
   U7189 : AOI22_X1 port map( A1 => n7418, A2 => n6202, B1 => n6201, B2 => 
                           n7259, ZN => n6389);
   U7190 : INV_X1 port map( A => n6246, ZN => n6342);
   U7191 : AOI21_X1 port map( B1 => intadd_29xBx1x, B2 => n6389, A => n6342, ZN
                           => n6548);
   U7192 : AOI22_X1 port map( A1 => n7418, A2 => n6204, B1 => n6203, B2 => 
                           n7231, ZN => n6368);
   U7193 : OAI22_X1 port map( A1 => n7231, A2 => n6206, B1 => n6205, B2 => 
                           n7418, ZN => n6388);
   U7194 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6368, B1 => n6388, 
                           B2 => n6456, ZN => n6552);
   U7195 : NOR2_X1 port map( A1 => n6552, A2 => ashr_25xSHx3x, ZN => n6208);
   U7196 : AOI21_X1 port map( B1 => n6548, B2 => ashr_25xSHx3x, A => n6208, ZN 
                           => n6881);
   U7197 : AND2_X1 port map( A1 => n7418, A2 => n6207, ZN => n7396);
   U7198 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6389, B1 => n7396, 
                           B2 => n6456, ZN => n6577);
   U7199 : AOI21_X1 port map( B1 => n6577, B2 => ashr_25xSHx3x, A => n6208, ZN 
                           => n6879);
   U7200 : AOI22_X1 port map( A1 => n6734, A2 => n6881, B1 => n6598, B2 => 
                           n6879, ZN => n6209);
   U7201 : OAI21_X1 port map( B1 => n6580, B2 => n6897, A => n6209, ZN => n6210
                           );
   U7202 : AOI211_X1 port map( C1 => ashr_25xAx3x, C2 => n6212, A => n6211, B 
                           => n6210, ZN => n6213);
   U7203 : OAI211_X1 port map( C1 => n6215, C2 => n7384, A => n6214, B => n6213
                           , ZN => n6216);
   U7204 : AOI211_X1 port map( C1 => n6218, C2 => n7327, A => n6217, B => n6216
                           , ZN => n6226);
   U7205 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(3), A2 => n6597,
                           B1 => n6547, B2 => ashr_25xAx3x, ZN => n6225);
   U7206 : NOR2_X1 port map( A1 => n5711, A2 => n6219, ZN => n6723);
   U7207 : NAND2_X1 port map( A1 => n6723, A2 => n6900, ZN => n6221);
   U7208 : AOI21_X1 port map( B1 => n6222, B2 => n6221, A => n6220, ZN => n6880
                           );
   U7209 : AOI22_X1 port map( A1 => n6453, A2 => n6880, B1 => n6305, B2 => 
                           n6223, ZN => n6224);
   U7210 : OAI211_X1 port map( C1 => n6226, C2 => n7533, A => n6225, B => n6224
                           , ZN => IF_ISAxN10940);
   U7211 : AOI22_X1 port map( A1 => n7311, A2 => n6228, B1 => n6227, B2 => 
                           n6900, ZN => n6595);
   U7212 : OAI22_X1 port map( A1 => n7406, A2 => n6230, B1 => n6229, B2 => 
                           n7269, ZN => n6231);
   U7213 : AOI21_X1 port map( B1 => n7207, B2 => n6595, A => n6231, ZN => n6269
                           );
   U7214 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6233, B1 => n6232, 
                           B2 => n6456, ZN => n6622);
   U7215 : OAI22_X1 port map( A1 => intadd_29xBx2x, A2 => n6622, B1 => n6234, 
                           B2 => n7415, ZN => n6235);
   U7216 : AOI211_X1 port map( C1 => n6236, C2 => n7422, A => n6720, B => n6235
                           , ZN => n6268);
   U7217 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn73, A2 => n7368, ZN 
                           => n6266);
   U7218 : MUX2_X1 port map( A => n6238, B => n6237, S => n7311, Z => n6593);
   U7219 : AOI22_X1 port map( A1 => n6593, A2 => n7376, B1 => n6592, B2 => 
                           n6365, ZN => n6919);
   U7220 : NAND2_X1 port map( A1 => n6919, A2 => n6350, ZN => n6946);
   U7221 : OAI22_X1 port map( A1 => n7118, A2 => n6240, B1 => n7397, B2 => 
                           n6239, ZN => n6243);
   U7222 : OAI22_X1 port map( A1 => n6251, A2 => n7387, B1 => n7386, B2 => 
                           n6241, ZN => n6242);
   U7223 : AOI211_X1 port map( C1 => n6678, C2 => n6946, A => n6243, B => n6242
                           , ZN => n6265);
   U7224 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx4x, B1 => 
                           ashr_25xAx3x, B2 => n7267, ZN => n6310);
   U7225 : AOI22_X1 port map( A1 => n7404, A2 => n6310, B1 => n6244, B2 => 
                           n7402, ZN => n6429);
   U7226 : AOI22_X1 port map( A1 => n7311, A2 => n6429, B1 => n6245, B2 => 
                           n6900, ZN => n6932);
   U7227 : INV_X1 port map( A => n6932, ZN => n6601);
   U7228 : OAI21_X1 port map( B1 => n7245, B2 => n6456, A => n6246, ZN => n6609
                           );
   U7229 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6253, B1 => n6252, 
                           B2 => intadd_25xBx0x, ZN => n6623);
   U7230 : OAI221_X1 port map( B1 => n7236, B2 => n6609, C1 => ashr_25xSHx3x, 
                           C2 => n6623, A => n6247, ZN => n6937);
   U7231 : AOI21_X1 port map( B1 => n7387, B2 => n6937, A => n7331, ZN => n6248
                           );
   U7232 : AOI21_X1 port map( B1 => n7307, B2 => n6601, A => n6248, ZN => n6264
                           );
   U7233 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx4x, B1 => 
                           ashr_25xAx3x, B2 => n7412, ZN => n6324);
   U7234 : MUX2_X1 port map( A => n6249, B => n6324, S => intadd_29xBx0x, Z => 
                           n6415);
   U7235 : OR2_X1 port map( A1 => n7231, A2 => n6250, ZN => n6418);
   U7236 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n6415, B1 => n6418, 
                           B2 => intadd_25xBx0x, ZN => n6607);
   U7237 : OAI221_X1 port map( B1 => n6251, B2 => n7389, C1 => ashr_25xAx4x, C2
                           => n7397, A => n7398, ZN => n6257);
   U7238 : NOR2_X1 port map( A1 => n7245, A2 => n6811, ZN => n6255);
   U7239 : AOI221_X1 port map( B1 => n6253, B2 => intadd_29xBx1x, C1 => n6252, 
                           C2 => intadd_25xBx0x, A => ashr_25xSHx3x, ZN => 
                           n6254);
   U7240 : AOI21_X1 port map( B1 => n6255, B2 => ashr_25xSHx3x, A => n6254, ZN 
                           => n6920);
   U7241 : OAI22_X1 port map( A1 => n6919, A2 => n6729, B1 => n6920, B2 => 
                           n6463, ZN => n6256);
   U7242 : AOI21_X1 port map( B1 => n7349, B2 => n6257, A => n6256, ZN => n6258
                           );
   U7243 : INV_X1 port map( A => n6258, ZN => n6262);
   U7244 : OAI22_X1 port map( A1 => n6260, A2 => n7384, B1 => n6259, B2 => 
                           n7316, ZN => n6261);
   U7245 : AOI211_X1 port map( C1 => n6607, C2 => n7018, A => n6262, B => n6261
                           , ZN => n6263);
   U7246 : NAND4_X1 port map( A1 => n6266, A2 => n6265, A3 => n6264, A4 => 
                           n6263, ZN => n6267);
   U7247 : AOI211_X1 port map( C1 => n6269, C2 => n6683, A => n6268, B => n6267
                           , ZN => n6271);
   U7248 : OAI22_X1 port map( A1 => n6271, A2 => n6717, B1 => n6270, B2 => 
                           n7439, ZN => IF_ISAxN10941);
   U7249 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(5), A2 => n6597,
                           B1 => n6547, B2 => ashr_25xAx5x, ZN => n6308);
   U7250 : INV_X1 port map( A => n6643, ZN => n6273);
   U7251 : AOI22_X1 port map( A1 => n6273, A2 => n7307, B1 => n7410, B2 => 
                           n6272, ZN => n6301);
   U7252 : AOI22_X1 port map( A1 => n6962, A2 => n6274, B1 => n6483, B2 => 
                           intadd_25xBx0x, ZN => n6636);
   U7253 : OAI22_X1 port map( A1 => n7236, A2 => n6636, B1 => n6275, B2 => 
                           n7415, ZN => n6276);
   U7254 : AOI211_X1 port map( C1 => n7422, C2 => n6277, A => n6720, B => n6276
                           , ZN => n6299);
   U7255 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn74, A2 => n7368, ZN 
                           => n6297);
   U7256 : OAI22_X1 port map( A1 => n7461, A2 => n7398, B1 => n6283, B2 => 
                           n7387, ZN => n6281);
   U7257 : INV_X1 port map( A => n6734, ZN => n6938);
   U7258 : OAI22_X1 port map( A1 => n6279, A2 => n6463, B1 => n6278, B2 => 
                           n6938, ZN => n6280);
   U7259 : AOI211_X1 port map( C1 => n6282, C2 => n7447, A => n6281, B => n6280
                           , ZN => n6296);
   U7260 : OAI22_X1 port map( A1 => n7461, A2 => n7389, B1 => n7386, B2 => 
                           n6283, ZN => n6294);
   U7261 : AOI22_X1 port map( A1 => n6941, A2 => n6285, B1 => n6284, B2 => 
                           n7309, ZN => n6640);
   U7262 : AOI22_X1 port map( A1 => n7275, A2 => n6287, B1 => n7400, B2 => 
                           n6286, ZN => n6288);
   U7263 : OAI211_X1 port map( C1 => n7376, C2 => n6640, A => n7192, B => n6288
                           , ZN => n6303);
   U7264 : OAI22_X1 port map( A1 => n6289, A2 => n6580, B1 => n6386, B2 => 
                           n6303, ZN => n6293);
   U7265 : OAI22_X1 port map( A1 => n6291, A2 => n7115, B1 => n6290, B2 => 
                           n7384, ZN => n6292);
   U7266 : AOI211_X1 port map( C1 => ashr_25xAx5x, C2 => n6294, A => n6293, B 
                           => n6292, ZN => n6295);
   U7267 : NAND3_X1 port map( A1 => n6297, A2 => n6296, A3 => n6295, ZN => 
                           n6298);
   U7268 : AOI211_X1 port map( C1 => n7018, C2 => n6646, A => n6299, B => n6298
                           , ZN => n6300);
   U7269 : OAI211_X1 port map( C1 => n6302, C2 => n7397, A => n6301, B => n6300
                           , ZN => n6306);
   U7270 : INV_X1 port map( A => n6303, ZN => n6304);
   U7271 : AOI22_X1 port map( A1 => n7029, A2 => n6306, B1 => n6305, B2 => 
                           n6304, ZN => n6307);
   U7272 : OAI211_X1 port map( C1 => n6309, C2 => n6632, A => n6308, B => n6307
                           , ZN => IF_ISAxN10942);
   U7273 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx6x, B1 => 
                           ashr_25xAx5x, B2 => n7267, ZN => n6428);
   U7274 : AOI22_X1 port map( A1 => n7404, A2 => n6428, B1 => n6310, B2 => 
                           n7402, ZN => n6515);
   U7275 : AOI22_X1 port map( A1 => n6941, A2 => n6515, B1 => n6513, B2 => 
                           n7309, ZN => n6978);
   U7276 : INV_X1 port map( A => n7307, ZN => n6967);
   U7277 : AOI22_X1 port map( A1 => n6962, A2 => n6312, B1 => n6311, B2 => 
                           intadd_25xBx0x, ZN => n6707);
   U7278 : AOI22_X1 port map( A1 => n7341, A2 => n6314, B1 => n7422, B2 => 
                           n6313, ZN => n6315);
   U7279 : OAI21_X1 port map( B1 => intadd_29xBx2x, B2 => n6707, A => n6315, ZN
                           => n6316);
   U7280 : OAI22_X1 port map( A1 => n6978, A2 => n6967, B1 => n6720, B2 => 
                           n6316, ZN => n6360);
   U7281 : NAND2_X1 port map( A1 => n6330, A2 => add_x_26xBx6x, ZN => n6317);
   U7282 : OAI22_X1 port map( A1 => n6318, A2 => n7384, B1 => n6317, B2 => 
                           n7316, ZN => n6359);
   U7283 : AOI22_X1 port map( A1 => n6941, A2 => n6320, B1 => n6319, B2 => 
                           n6900, ZN => n6686);
   U7284 : OAI22_X1 port map( A1 => n7406, A2 => n6322, B1 => n7269, B2 => 
                           n6321, ZN => n6323);
   U7285 : AOI211_X1 port map( C1 => n6686, C2 => n7207, A => n7349, B => n6323
                           , ZN => n6345);
   U7286 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx6x, B1 => 
                           ashr_25xAx5x, B2 => n7412, ZN => n6414);
   U7287 : AOI22_X1 port map( A1 => n7418, A2 => n6414, B1 => n6324, B2 => 
                           n7259, ZN => n6504);
   U7288 : AOI22_X1 port map( A1 => n6962, A2 => n6504, B1 => n6502, B2 => 
                           intadd_25xBx0x, ZN => n6697);
   U7289 : INV_X1 port map( A => n6697, ZN => n6981);
   U7290 : AOI22_X1 port map( A1 => n6325, A2 => n6345, B1 => n7018, B2 => 
                           n6981, ZN => n6328);
   U7291 : OAI221_X1 port map( B1 => n7462, B2 => n6330, C1 => n6326, C2 => 
                           ashr_25xAx6x, A => n7327, ZN => n6327);
   U7292 : OAI211_X1 port map( C1 => n7316, C2 => n6329, A => n6328, B => n6327
                           , ZN => n6358);
   U7293 : AOI221_X1 port map( B1 => n6330, B2 => n7398, C1 => n7389, C2 => 
                           n7398, A => n7462, ZN => n6334);
   U7294 : AOI21_X1 port map( B1 => n7320, B2 => ashr_25xAx6x, A => n7251, ZN 
                           => n6331);
   U7295 : OAI22_X1 port map( A1 => n6332, A2 => n6331, B1 => n6330, B2 => 
                           n7387, ZN => n6333);
   U7296 : AOI211_X1 port map( C1 => n6335, C2 => n7447, A => n6334, B => n6333
                           , ZN => n6354);
   U7297 : INV_X1 port map( A => n6365, ZN => n6568);
   U7298 : INV_X1 port map( A => n6672, ZN => n6336);
   U7299 : OAI221_X1 port map( B1 => n7311, B2 => n6681, C1 => n7309, C2 => 
                           n6682, A => n7376, ZN => n6349);
   U7300 : OAI21_X1 port map( B1 => n6568, B2 => n6336, A => n6349, ZN => n6982
                           );
   U7301 : INV_X1 port map( A => n6711, ZN => n7300);
   U7302 : NAND2_X1 port map( A1 => intadd_29xBx1x, A2 => n7300, ZN => n6341);
   U7303 : AOI22_X1 port map( A1 => n7418, A2 => n6338, B1 => n6337, B2 => 
                           n7259, ZN => n6339);
   U7304 : AOI22_X1 port map( A1 => n6962, A2 => n6340, B1 => n6339, B2 => 
                           intadd_25xBx0x, ZN => n6708);
   U7305 : NAND2_X1 port map( A1 => n7236, A2 => n6708, ZN => n6344);
   U7306 : OAI21_X1 port map( B1 => n7236, B2 => n6341, A => n6344, ZN => n6959
                           );
   U7307 : AOI22_X1 port map( A1 => n6715, A2 => n6982, B1 => n6598, B2 => 
                           n6959, ZN => n6353);
   U7308 : AOI211_X1 port map( C1 => n7300, C2 => intadd_29xBx1x, A => n6343, B
                           => n6342, ZN => n6673);
   U7309 : OAI21_X1 port map( B1 => n7236, B2 => n6673, A => n6344, ZN => n6988
                           );
   U7310 : AOI22_X1 port map( A1 => n6346, A2 => n6345, B1 => n6734, B2 => 
                           n6988, ZN => n6352);
   U7311 : INV_X1 port map( A => n6676, ZN => n6347);
   U7312 : OAI21_X1 port map( B1 => n6672, B2 => n6347, A => n6365, ZN => n6348
                           );
   U7313 : NAND3_X1 port map( A1 => n6350, A2 => n6349, A3 => n6348, ZN => 
                           n6969);
   U7314 : NAND2_X1 port map( A1 => n6678, A2 => n6969, ZN => n6351);
   U7315 : NAND4_X1 port map( A1 => n6354, A2 => n6353, A3 => n6352, A4 => 
                           n6351, ZN => n6355);
   U7316 : AOI21_X1 port map( B1 => DP_OP_719J14_125_1055xn75, B2 => n7159, A 
                           => n6355, ZN => n6356);
   U7317 : INV_X1 port map( A => n6356, ZN => n6357);
   U7318 : NOR4_X1 port map( A1 => n6360, A2 => n6359, A3 => n6358, A4 => n6357
                           , ZN => n6362);
   U7319 : OAI22_X1 port map( A1 => n6362, A2 => n6717, B1 => n6361, B2 => 
                           n7439, ZN => IF_ISAxN10943);
   U7320 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(7), ZN => n7442);
   U7321 : INV_X1 port map( A => n6363, ZN => n6364);
   U7322 : AOI22_X1 port map( A1 => n6941, A2 => n6364, B1 => n6574, B2 => 
                           n6900, ZN => n6750);
   U7323 : NOR2_X1 port map( A1 => n6750, A2 => n7207, ZN => n6373);
   U7324 : AOI21_X1 port map( B1 => n6365, B2 => n6723, A => n6373, ZN => n7011
                           );
   U7325 : AOI22_X1 port map( A1 => n7418, A2 => n6367, B1 => n6366, B2 => 
                           n7259, ZN => n6560);
   U7326 : AOI22_X1 port map( A1 => n6962, A2 => n6560, B1 => n6563, B2 => 
                           intadd_25xBx0x, ZN => n7001);
   U7327 : AOI22_X1 port map( A1 => n6962, A2 => n6369, B1 => n6368, B2 => 
                           n6456, ZN => n6719);
   U7328 : OAI22_X1 port map( A1 => intadd_29xBx2x, A2 => n6719, B1 => n6370, 
                           B2 => n7415, ZN => n6371);
   U7329 : AOI211_X1 port map( C1 => n7422, C2 => n6372, A => n6720, B => n6371
                           , ZN => n6408);
   U7330 : OR2_X1 port map( A1 => n6520, A2 => n6373, ZN => n7019);
   U7331 : AOI22_X1 port map( A1 => n7404, A2 => n6375, B1 => n6374, B2 => 
                           n7402, ZN => n6567);
   U7332 : AOI22_X1 port map( A1 => n6941, A2 => n6567, B1 => n6564, B2 => 
                           n7309, ZN => n7005);
   U7333 : INV_X1 port map( A => n7005, ZN => n7372);
   U7334 : AOI22_X1 port map( A1 => n6678, A2 => n7019, B1 => n7372, B2 => 
                           n7307, ZN => n6405);
   U7335 : NOR2_X1 port map( A1 => n6399, A2 => n7397, ZN => n6379);
   U7336 : AOI221_X1 port map( B1 => n7327, B2 => n6399, C1 => n7253, C2 => 
                           ashr_25xAx7x, A => n7322, ZN => n6376);
   U7337 : INV_X1 port map( A => n6376, ZN => n6378);
   U7338 : MUX2_X1 port map( A => n6379, B => n6378, S => n6377, Z => n6403);
   U7339 : AOI22_X1 port map( A1 => n6941, A2 => n6381, B1 => n6380, B2 => 
                           n7309, ZN => n6748);
   U7340 : AOI22_X1 port map( A1 => n7275, A2 => n6383, B1 => n7400, B2 => 
                           n6382, ZN => n6384);
   U7341 : OAI211_X1 port map( C1 => n7376, C2 => n6748, A => n7192, B => n6384
                           , ZN => n6385);
   U7342 : AOI21_X1 port map( B1 => n6387, B2 => n6386, A => n6385, ZN => n6402
                           );
   U7343 : INV_X1 port map( A => n6388, ZN => n6390);
   U7344 : AOI22_X1 port map( A1 => n6962, A2 => n6390, B1 => n6389, B2 => 
                           n6456, ZN => n6722);
   U7345 : NOR2_X1 port map( A1 => n6722, A2 => ashr_25xSHx3x, ZN => n6391);
   U7346 : AOI21_X1 port map( B1 => n7396, B2 => n6417, A => n6391, ZN => n7008
                           );
   U7347 : NOR2_X1 port map( A1 => n7435, A2 => n7236, ZN => n6633);
   U7348 : NOR2_X1 port map( A1 => n6633, A2 => n6391, ZN => n7012);
   U7349 : OAI22_X1 port map( A1 => n7008, A2 => n6463, B1 => n7012, B2 => 
                           n6938, ZN => n6401);
   U7350 : NOR2_X1 port map( A1 => n7316, A2 => add_x_26xBx7x, ZN => n6392);
   U7351 : AOI211_X1 port map( C1 => n7320, C2 => add_x_26xBx7x, A => n7251, B 
                           => n6392, ZN => n6398);
   U7352 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn76, A2 => n7368, ZN 
                           => n6397);
   U7353 : OAI22_X1 port map( A1 => n7387, A2 => n6394, B1 => n7118, B2 => 
                           n6393, ZN => n6395);
   U7354 : AOI21_X1 port map( B1 => intadd_25xSUMx5x, B2 => n7276, A => n6395, 
                           ZN => n6396);
   U7355 : OAI211_X1 port map( C1 => n6399, C2 => n6398, A => n6397, B => n6396
                           , ZN => n6400);
   U7356 : NOR4_X1 port map( A1 => n6403, A2 => n6402, A3 => n6401, A4 => n6400
                           , ZN => n6404);
   U7357 : OAI211_X1 port map( C1 => n6406, C2 => n7255, A => n6405, B => n6404
                           , ZN => n6407);
   U7358 : AOI211_X1 port map( C1 => n7018, C2 => n7001, A => n6408, B => n6407
                           , ZN => n6409);
   U7359 : OAI222_X1 port map( A1 => n7442, A2 => n7439, B1 => n6632, B2 => 
                           n7011, C1 => n7533, C2 => n6409, ZN => IF_ISAxN10944
                           );
   U7360 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(8), ZN => n7443);
   U7361 : NOR2_X1 port map( A1 => n7049, A2 => n7207, ZN => n6435);
   U7362 : NOR2_X1 port map( A1 => n7427, A2 => n7533, ZN => n6596);
   U7363 : AOI22_X1 port map( A1 => n7376, A2 => n6411, B1 => n6410, B2 => 
                           n7207, ZN => n6437);
   U7364 : AOI22_X1 port map( A1 => n6453, A2 => n6435, B1 => n6596, B2 => 
                           n6437, ZN => n6452);
   U7365 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn77, A2 => n7368, ZN 
                           => n6434);
   U7366 : AOI21_X1 port map( B1 => n7236, B2 => n7042, A => n6633, ZN => n6412
                           );
   U7367 : INV_X1 port map( A => n6412, ZN => n7060);
   U7368 : AND2_X1 port map( A1 => intadd_29xBx2x, A2 => n7042, ZN => n6413);
   U7369 : AOI22_X1 port map( A1 => n6734, A2 => n7060, B1 => n6598, B2 => 
                           n6413, ZN => n6433);
   U7370 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx8x, B1 => 
                           ashr_25xAx7x, B2 => n7412, ZN => n6503);
   U7371 : AOI22_X1 port map( A1 => n7418, A2 => n6503, B1 => n6414, B2 => 
                           n7231, ZN => n6606);
   U7372 : INV_X1 port map( A => n6415, ZN => n6416);
   U7373 : AOI22_X1 port map( A1 => n6962, A2 => n6606, B1 => n6416, B2 => 
                           n6456, ZN => n6765);
   U7374 : INV_X1 port map( A => n6417, ZN => n6562);
   U7375 : OAI22_X1 port map( A1 => n6765, A2 => ashr_25xSHx3x, B1 => n6418, B2
                           => n6562, ZN => n7040);
   U7376 : OAI21_X1 port map( B1 => n6419, B2 => n7389, A => n7398, ZN => n6420
                           );
   U7377 : AND2_X1 port map( A1 => n6421, A2 => n6420, ZN => n6427);
   U7378 : INV_X1 port map( A => n6422, ZN => n6425);
   U7379 : NOR2_X1 port map( A1 => n6423, A2 => intadd_29xBx2x, ZN => n6424);
   U7380 : AOI211_X1 port map( C1 => intadd_29xBx2x, C2 => n6425, A => n6720, B
                           => n6424, ZN => n6426);
   U7381 : AOI211_X1 port map( C1 => n7420, C2 => n7040, A => n6427, B => n6426
                           , ZN => n6432);
   U7382 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx8x, B1 => 
                           ashr_25xAx7x, B2 => n7267, ZN => n6514);
   U7383 : AOI22_X1 port map( A1 => n7404, A2 => n6514, B1 => n6428, B2 => 
                           n7402, ZN => n6600);
   U7384 : AOI22_X1 port map( A1 => n6941, A2 => n6600, B1 => n6429, B2 => 
                           n6900, ZN => n6771);
   U7385 : OAI22_X1 port map( A1 => n6771, A2 => n7207, B1 => n6430, B2 => 
                           n6568, ZN => n7055);
   U7386 : NAND2_X1 port map( A1 => n7409, A2 => n7055, ZN => n6431);
   U7387 : NAND4_X1 port map( A1 => n6434, A2 => n6433, A3 => n6432, A4 => 
                           n6431, ZN => n6450);
   U7388 : NOR2_X1 port map( A1 => n6520, A2 => n6435, ZN => n7034);
   U7389 : INV_X1 port map( A => n7034, ZN => n6436);
   U7390 : AOI22_X1 port map( A1 => n6653, A2 => n6437, B1 => n6678, B2 => 
                           n6436, ZN => n6447);
   U7391 : INV_X1 port map( A => intadd_25xSUMx6x, ZN => n6442);
   U7392 : AOI22_X1 port map( A1 => n7320, A2 => n6439, B1 => n6438, B2 => 
                           n7447, ZN => n6441);
   U7393 : OAI21_X1 port map( B1 => add_x_26xBx8x, B2 => ashr_25xAx8x, A => 
                           n7251, ZN => n6440);
   U7394 : OAI211_X1 port map( C1 => n6442, C2 => n7384, A => n6441, B => n6440
                           , ZN => n6443);
   U7395 : AOI221_X1 port map( B1 => n6445, B2 => n7327, C1 => n6444, C2 => 
                           n7073, A => n6443, ZN => n6446);
   U7396 : OAI211_X1 port map( C1 => n6448, C2 => n7255, A => n6447, B => n6446
                           , ZN => n6449);
   U7397 : OAI21_X1 port map( B1 => n6450, B2 => n6449, A => n7029, ZN => n6451
                           );
   U7398 : OAI211_X1 port map( C1 => n7439, C2 => n7443, A => n6452, B => n6451
                           , ZN => IF_ISAxN10945);
   U7399 : NAND2_X1 port map( A1 => n7376, A2 => n6453, ZN => n6591);
   U7400 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(9), A2 => n6597,
                           B1 => n6547, B2 => ashr_25xAx9x, ZN => n6499);
   U7401 : AOI22_X1 port map( A1 => n7376, A2 => n6455, B1 => n6454, B2 => 
                           n7207, ZN => n6495);
   U7402 : AOI22_X1 port map( A1 => n6962, A2 => n6458, B1 => n6457, B2 => 
                           n6456, ZN => n6814);
   U7403 : INV_X1 port map( A => n6814, ZN => n6460);
   U7404 : OAI22_X1 port map( A1 => n6460, A2 => ashr_25xSHx3x, B1 => n6459, B2
                           => n6562, ZN => n7089);
   U7405 : AOI21_X1 port map( B1 => n7236, B2 => n6461, A => n6633, ZN => n7096
                           );
   U7406 : NAND2_X1 port map( A1 => n7236, A2 => n6462, ZN => n7082);
   U7407 : OAI22_X1 port map( A1 => n7096, A2 => n6938, B1 => n6463, B2 => 
                           n7082, ZN => n6464);
   U7408 : AOI21_X1 port map( B1 => n7420, B2 => n7089, A => n6464, ZN => n6493
                           );
   U7409 : AOI22_X1 port map( A1 => n6941, A2 => n6466, B1 => n6465, B2 => 
                           n6900, ZN => n6818);
   U7410 : INV_X1 port map( A => n6467, ZN => n6468);
   U7411 : OAI22_X1 port map( A1 => n7207, A2 => n6818, B1 => n6468, B2 => 
                           n6568, ZN => n7094);
   U7412 : INV_X1 port map( A => n6469, ZN => n6470);
   U7413 : AOI21_X1 port map( B1 => n6470, B2 => n7376, A => n6520, ZN => n7085
                           );
   U7414 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn78, A2 => n7368, ZN 
                           => n6475);
   U7415 : NAND3_X1 port map( A1 => n6480, A2 => n7253, A3 => ashr_25xAx9x, ZN 
                           => n6471);
   U7416 : OAI21_X1 port map( B1 => n7118, B2 => n6472, A => n6471, ZN => n6473
                           );
   U7417 : AOI21_X1 port map( B1 => n7251, B2 => add_x_26xBx9x, A => n6473, ZN 
                           => n6474);
   U7418 : OAI211_X1 port map( C1 => n7085, C2 => n6580, A => n6475, B => n6474
                           , ZN => n6491);
   U7419 : NOR2_X1 port map( A1 => n6481, A2 => n6476, ZN => n6477);
   U7420 : AOI22_X1 port map( A1 => n6478, A2 => n7073, B1 => n6477, B2 => 
                           n7320, ZN => n6489);
   U7421 : AOI22_X1 port map( A1 => intadd_25xSUMx7x, A2 => n7276, B1 => n6479,
                           B2 => n7127, ZN => n6488);
   U7422 : OAI211_X1 port map( C1 => n7322, C2 => n7327, A => n6481, B => n6480
                           , ZN => n6487);
   U7423 : AOI22_X1 port map( A1 => n6962, A2 => n6483, B1 => n6482, B2 => 
                           intadd_25xBx0x, ZN => n6485);
   U7424 : INV_X1 port map( A => n6720, ZN => n6706);
   U7425 : OAI221_X1 port map( B1 => n7236, B2 => n6485, C1 => ashr_25xSHx3x, 
                           C2 => n6484, A => n6706, ZN => n6486);
   U7426 : NAND4_X1 port map( A1 => n6489, A2 => n6488, A3 => n6487, A4 => 
                           n6486, ZN => n6490);
   U7427 : AOI211_X1 port map( C1 => n7409, C2 => n7094, A => n6491, B => n6490
                           , ZN => n6492);
   U7428 : OAI211_X1 port map( C1 => n6495, C2 => n6494, A => n6493, B => n6492
                           , ZN => n6497);
   U7429 : INV_X1 port map( A => n6495, ZN => n6496);
   U7430 : AOI22_X1 port map( A1 => n7029, A2 => n6497, B1 => n6596, B2 => 
                           n6496, ZN => n6498);
   U7431 : OAI211_X1 port map( C1 => n7083, C2 => n6591, A => n6499, B => n6498
                           , ZN => IF_ISAxN10946);
   U7432 : INV_X1 port map( A => n6500, ZN => n7124);
   U7433 : INV_X1 port map( A => intadd_25xSUMx8x, ZN => n6543);
   U7434 : OAI21_X1 port map( B1 => n7466, B2 => ashr_25xAx10x, A => n6501, ZN 
                           => n6506);
   U7435 : INV_X1 port map( A => n6502, ZN => n6505);
   U7436 : AOI22_X1 port map( A1 => n7414, A2 => ashr_25xAx10x, B1 => 
                           ashr_25xAx9x, B2 => n7412, ZN => n6605);
   U7437 : AOI22_X1 port map( A1 => n7418, A2 => n6605, B1 => n6503, B2 => 
                           n7231, ZN => n6696);
   U7438 : AOI22_X1 port map( A1 => n6962, A2 => n6696, B1 => n6504, B2 => 
                           intadd_25xBx0x, ZN => n6853);
   U7439 : OAI22_X1 port map( A1 => n6505, A2 => n6562, B1 => n6853, B2 => 
                           ashr_25xSHx3x, ZN => n7139);
   U7440 : AOI22_X1 port map( A1 => n7073, A2 => n6506, B1 => n7420, B2 => 
                           n7139, ZN => n6542);
   U7441 : AOI22_X1 port map( A1 => add_x_26xBx10x, A2 => n7251, B1 => n6507, 
                           B2 => n7447, ZN => n6511);
   U7442 : OAI221_X1 port map( B1 => n7236, B2 => n6509, C1 => ashr_25xSHx3x, 
                           C2 => n6508, A => n6706, ZN => n6510);
   U7443 : OAI211_X1 port map( C1 => n7316, C2 => n6512, A => n6511, B => n6510
                           , ZN => n6539);
   U7444 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn79, A2 => n7159, ZN 
                           => n6537);
   U7445 : INV_X1 port map( A => n6513, ZN => n6516);
   U7446 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx10x, B1 => 
                           ashr_25xAx9x, B2 => n7086, ZN => n6599);
   U7447 : AOI22_X1 port map( A1 => n7404, A2 => n6599, B1 => n6514, B2 => 
                           n7402, ZN => n6700);
   U7448 : AOI22_X1 port map( A1 => n6941, A2 => n6700, B1 => n6515, B2 => 
                           n7309, ZN => n6849);
   U7449 : OAI22_X1 port map( A1 => n6516, A2 => n6568, B1 => n6849, B2 => 
                           n7207, ZN => n7138);
   U7450 : NAND2_X1 port map( A1 => n7236, A2 => n6517, ZN => n7143);
   U7451 : INV_X1 port map( A => n7143, ZN => n6518);
   U7452 : AOI22_X1 port map( A1 => n7409, A2 => n7138, B1 => n6598, B2 => 
                           n6518, ZN => n6536);
   U7453 : INV_X1 port map( A => n6519, ZN => n6522);
   U7454 : INV_X1 port map( A => n6520, ZN => n6521);
   U7455 : OAI21_X1 port map( B1 => n6522, B2 => n7207, A => n6521, ZN => n7121
                           );
   U7456 : AND2_X1 port map( A1 => n6523, A2 => n7376, ZN => n6524);
   U7457 : AOI21_X1 port map( B1 => n6525, B2 => n7207, A => n6524, ZN => n6527
                           );
   U7458 : INV_X1 port map( A => n6527, ZN => n6533);
   U7459 : INV_X1 port map( A => n6633, ZN => n6675);
   U7460 : NAND3_X1 port map( A1 => n6675, A2 => n6526, A3 => n7143, ZN => 
                           n7135);
   U7461 : AOI22_X1 port map( A1 => n6653, A2 => n6527, B1 => n6734, B2 => 
                           n7135, ZN => n6532);
   U7462 : OAI21_X1 port map( B1 => n6528, B2 => n7389, A => n7398, ZN => n6529
                           );
   U7463 : NAND2_X1 port map( A1 => n6530, A2 => n6529, ZN => n6531);
   U7464 : OAI211_X1 port map( C1 => n7427, C2 => n6533, A => n6532, B => n6531
                           , ZN => n6534);
   U7465 : AOI21_X1 port map( B1 => n6678, B2 => n7121, A => n6534, ZN => n6535
                           );
   U7466 : NAND3_X1 port map( A1 => n6537, A2 => n6536, A3 => n6535, ZN => 
                           n6538);
   U7467 : AOI211_X1 port map( C1 => n6540, C2 => n7320, A => n6539, B => n6538
                           , ZN => n6541);
   U7468 : OAI211_X1 port map( C1 => n6543, C2 => n7384, A => n6542, B => n6541
                           , ZN => n6544);
   U7469 : AOI22_X1 port map( A1 => n6597, A2 => fromMemoryPortxLOADEDDATAx(10)
                           , B1 => n7029, B2 => n6544, ZN => n6546);
   U7470 : NAND2_X1 port map( A1 => n6547, A2 => ashr_25xAx10x, ZN => n6545);
   U7471 : OAI211_X1 port map( C1 => n6591, C2 => n7124, A => n6546, B => n6545
                           , ZN => IF_ISAxN10947);
   U7472 : AOI22_X1 port map( A1 => n6941, A2 => n6574, B1 => n6723, B2 => 
                           n7309, ZN => n7194);
   U7473 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(11), A2 => n6597
                           , B1 => n6547, B2 => ashr_25xAx11x, ZN => n6590);
   U7474 : INV_X1 port map( A => n6548, ZN => n6549);
   U7475 : AOI21_X1 port map( B1 => intadd_29xBx2x, B2 => n6549, A => n6633, ZN
                           => n7165);
   U7476 : NOR2_X1 port map( A1 => intadd_27xAx0x, A2 => add_x_26xBx11x, ZN => 
                           n6550);
   U7477 : AOI22_X1 port map( A1 => intadd_25xSUMx9x, A2 => n7276, B1 => n6550,
                           B2 => n7410, ZN => n6586);
   U7478 : AOI221_X1 port map( B1 => intadd_27xAx0x, B2 => n7398, C1 => n7389, 
                           C2 => n7398, A => n7467, ZN => n6584);
   U7479 : NAND2_X1 port map( A1 => intadd_27xAx0x, A2 => add_x_26xBx11x, ZN =>
                           n6556);
   U7480 : OAI221_X1 port map( B1 => n7236, B2 => n6552, C1 => ashr_25xSHx3x, 
                           C2 => n6551, A => n6706, ZN => n6555);
   U7481 : OAI221_X1 port map( B1 => intadd_27xAx0x, B2 => n7467, C1 => 
                           ashr_25xAx11x, C2 => n6553, A => n7327, ZN => n6554)
                           ;
   U7482 : OAI211_X1 port map( C1 => n7316, C2 => n6556, A => n6555, B => n6554
                           , ZN => n6583);
   U7483 : OAI221_X1 port map( B1 => n7251, B2 => n7320, C1 => n7251, C2 => 
                           ashr_25xAx11x, A => add_x_26xBx11x, ZN => n6571);
   U7484 : AOI22_X1 port map( A1 => n7418, A2 => n6558, B1 => n6557, B2 => 
                           n7259, ZN => n6726);
   U7485 : AND2_X1 port map( A1 => n6726, A2 => intadd_29xBx1x, ZN => n6559);
   U7486 : AOI21_X1 port map( B1 => n6560, B2 => intadd_25xBx0x, A => n6559, ZN
                           => n6908);
   U7487 : INV_X1 port map( A => n6908, ZN => n6561);
   U7488 : OAI22_X1 port map( A1 => n6563, A2 => n6562, B1 => n6561, B2 => 
                           ashr_25xSHx3x, ZN => n7163);
   U7489 : INV_X1 port map( A => n6564, ZN => n6569);
   U7490 : AOI22_X1 port map( A1 => n7404, A2 => n6566, B1 => n6565, B2 => 
                           n7402, ZN => n6732);
   U7491 : AOI22_X1 port map( A1 => n6941, A2 => n6732, B1 => n6567, B2 => 
                           n6900, ZN => n6903);
   U7492 : OAI22_X1 port map( A1 => n6569, A2 => n6568, B1 => n6903, B2 => 
                           n7207, ZN => n7189);
   U7493 : AOI22_X1 port map( A1 => n7420, A2 => n7163, B1 => n7409, B2 => 
                           n7189, ZN => n6570);
   U7494 : OAI211_X1 port map( C1 => n7118, C2 => n6572, A => n6571, B => n6570
                           , ZN => n6582);
   U7495 : NAND2_X1 port map( A1 => n7413, A2 => n7269, ZN => n6677);
   U7496 : INV_X1 port map( A => n6677, ZN => n6573);
   U7497 : AOI21_X1 port map( B1 => n7400, B2 => n6574, A => n6573, ZN => n7191
                           );
   U7498 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn80, A2 => n7368, ZN 
                           => n6579);
   U7499 : MUX2_X1 port map( A => n6576, B => n6575, S => n7376, Z => n6587);
   U7500 : NOR2_X1 port map( A1 => n6577, A2 => ashr_25xSHx3x, ZN => n7167);
   U7501 : AOI22_X1 port map( A1 => n6653, A2 => n6587, B1 => n6598, B2 => 
                           n7167, ZN => n6578);
   U7502 : OAI211_X1 port map( C1 => n7191, C2 => n6580, A => n6579, B => n6578
                           , ZN => n6581);
   U7503 : NOR4_X1 port map( A1 => n6584, A2 => n6583, A3 => n6582, A4 => n6581
                           , ZN => n6585);
   U7504 : OAI211_X1 port map( C1 => n7165, C2 => n6938, A => n6586, B => n6585
                           , ZN => n6588);
   U7505 : AOI22_X1 port map( A1 => n7029, A2 => n6588, B1 => n6596, B2 => 
                           n6587, ZN => n6589);
   U7506 : OAI211_X1 port map( C1 => n7194, C2 => n6591, A => n6590, B => n6589
                           , ZN => IF_ISAxN10948);
   U7507 : NAND2_X1 port map( A1 => n7400, A2 => n6592, ZN => n7239);
   U7508 : INV_X1 port map( A => n6593, ZN => n6594);
   U7509 : AOI22_X1 port map( A1 => n7376, A2 => n6595, B1 => n6594, B2 => 
                           n7207, ZN => n6603);
   U7510 : AOI22_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(12), A2 => n6597
                           , B1 => n6596, B2 => n6603, ZN => n6631);
   U7511 : NAND2_X1 port map( A1 => n7341, A2 => n6598, ZN => n6741);
   U7512 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx12x, B1 => 
                           ashr_25xAx11x, B2 => n7399, ZN => n6699);
   U7513 : AOI22_X1 port map( A1 => n7404, A2 => n6699, B1 => n6599, B2 => 
                           n7402, ZN => n6761);
   U7514 : AOI22_X1 port map( A1 => n6941, A2 => n6761, B1 => n6600, B2 => 
                           n7309, ZN => n6931);
   U7515 : NOR2_X1 port map( A1 => n6601, A2 => n7376, ZN => n6602);
   U7516 : AOI21_X1 port map( B1 => n7376, B2 => n6931, A => n6602, ZN => n7216
                           );
   U7517 : AOI22_X1 port map( A1 => n7216, A2 => n7409, B1 => n6603, B2 => 
                           n6653, ZN => n6604);
   U7518 : INV_X1 port map( A => n6604, ZN => n6621);
   U7519 : AOI22_X1 port map( A1 => n7333, A2 => ashr_25xAx12x, B1 => 
                           ashr_25xAx11x, B2 => n7412, ZN => n6695);
   U7520 : AOI22_X1 port map( A1 => n7418, A2 => n6695, B1 => n6605, B2 => 
                           n7259, ZN => n6769);
   U7521 : MUX2_X1 port map( A => n6606, B => n6769, S => intadd_29xBx1x, Z => 
                           n6942);
   U7522 : INV_X1 port map( A => n6607, ZN => n6930);
   U7523 : NOR2_X1 port map( A1 => n6930, A2 => intadd_29xBx2x, ZN => n6608);
   U7524 : AOI21_X1 port map( B1 => intadd_29xBx2x, B2 => n6942, A => n6608, ZN
                           => n7214);
   U7525 : AOI21_X1 port map( B1 => n7236, B2 => n6609, A => n6633, ZN => n7221
                           );
   U7526 : OAI22_X1 port map( A1 => n7214, A2 => n7343, B1 => n7221, B2 => 
                           n6938, ZN => n6620);
   U7527 : OAI22_X1 port map( A1 => n6611, A2 => n7384, B1 => n6610, B2 => 
                           n7316, ZN => n6619);
   U7528 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn81, A2 => n7159, ZN 
                           => n6617);
   U7529 : NAND2_X1 port map( A1 => n6677, A2 => n7239, ZN => n7228);
   U7530 : AOI22_X1 port map( A1 => n6678, A2 => n7228, B1 => n6612, B2 => 
                           n7447, ZN => n6616);
   U7531 : OAI22_X1 port map( A1 => intadd_27xBx1x, A2 => n7227, B1 => n6613, 
                           B2 => n7397, ZN => n6614);
   U7532 : AOI21_X1 port map( B1 => n7322, B2 => n6626, A => n6614, ZN => n6615
                           );
   U7533 : NAND3_X1 port map( A1 => n6617, A2 => n6616, A3 => n6615, ZN => 
                           n6618);
   U7534 : NOR4_X1 port map( A1 => n6621, A2 => n6620, A3 => n6619, A4 => n6618
                           , ZN => n6625);
   U7535 : OAI221_X1 port map( B1 => intadd_29xBx2x, B2 => n6623, C1 => 
                           ashr_25xSHx3x, C2 => n6622, A => n6706, ZN => n6624)
                           ;
   U7536 : OAI211_X1 port map( C1 => n7245, C2 => n6741, A => n6625, B => n6624
                           , ZN => n6629);
   U7537 : AOI221_X1 port map( B1 => n7327, B2 => n7468, C1 => n7253, C2 => 
                           n6626, A => n7251, ZN => n6627);
   U7538 : OAI221_X1 port map( B1 => intadd_27xBx1x, B2 => n7386, C1 => 
                           add_x_26xBx12x, C2 => n7255, A => n6627, ZN => n6628
                           );
   U7539 : OAI221_X1 port map( B1 => n6629, B2 => ashr_25xAx12x, C1 => n6629, 
                           C2 => n6628, A => n7029, ZN => n6630);
   U7540 : OAI211_X1 port map( C1 => n6632, C2 => n7239, A => n6631, B => n6630
                           , ZN => IF_ISAxN10949);
   U7541 : AOI21_X1 port map( B1 => intadd_29xBx2x, B2 => n6634, A => n6633, ZN
                           => n7287);
   U7542 : INV_X1 port map( A => n7227, ZN => n7380);
   U7543 : AOI22_X1 port map( A1 => n6635, A2 => n7447, B1 => add_x_26xBx13x, 
                           B2 => n7380, ZN => n6639);
   U7544 : OAI221_X1 port map( B1 => intadd_29xBx2x, B2 => n6637, C1 => 
                           ashr_25xSHx3x, C2 => n6636, A => n6706, ZN => n6638)
                           ;
   U7545 : OAI211_X1 port map( C1 => n7287, C2 => n6938, A => n6639, B => n6638
                           , ZN => n6668);
   U7546 : AND2_X1 port map( A1 => n6640, A2 => n7376, ZN => n6641);
   U7547 : AOI21_X1 port map( B1 => n6642, B2 => n7207, A => n6641, ZN => n6666
                           );
   U7548 : AOI22_X1 port map( A1 => n7376, A2 => n6644, B1 => n6643, B2 => 
                           n7207, ZN => n7282);
   U7549 : NAND2_X1 port map( A1 => n7400, A2 => n6645, ZN => n7284);
   U7550 : AOI22_X1 port map( A1 => n7236, A2 => n6647, B1 => n6646, B2 => 
                           ashr_25xSHx3x, ZN => n7283);
   U7551 : OAI22_X1 port map( A1 => n6729, A2 => n7284, B1 => n7343, B2 => 
                           n7283, ZN => n6648);
   U7552 : AOI21_X1 port map( B1 => n7409, B2 => n7282, A => n6648, ZN => n6665
                           );
   U7553 : INV_X1 port map( A => intadd_25xSUMx11x, ZN => n6650);
   U7554 : OAI22_X1 port map( A1 => n6650, A2 => n7384, B1 => n6649, B2 => 
                           n7316, ZN => n6663);
   U7555 : INV_X1 port map( A => n6666, ZN => n6654);
   U7556 : INV_X1 port map( A => n6651, ZN => n6652);
   U7557 : OAI21_X1 port map( B1 => n6652, B2 => n7269, A => n6677, ZN => n7277
                           );
   U7558 : AOI222_X1 port map( A1 => n6654, A2 => n6653, B1 => n6678, B2 => 
                           n7277, C1 => n7368, C2 => DP_OP_719J14_125_1055xn82,
                           ZN => n6655);
   U7559 : INV_X1 port map( A => n6655, ZN => n6662);
   U7560 : AOI21_X1 port map( B1 => n6657, B2 => n6656, A => n7397, ZN => n6661
                           );
   U7561 : OAI221_X1 port map( B1 => intadd_27xBx2x, B2 => n7386, C1 => 
                           add_x_26xBx13x, C2 => n7255, A => n7387, ZN => n6658
                           );
   U7562 : AOI21_X1 port map( B1 => n7253, B2 => n6669, A => n6658, ZN => n6659
                           );
   U7563 : OAI22_X1 port map( A1 => n7286, A2 => n6741, B1 => intadd_27xAx2x, 
                           B2 => n6659, ZN => n6660);
   U7564 : NOR4_X1 port map( A1 => n6663, A2 => n6662, A3 => n6661, A4 => n6660
                           , ZN => n6664);
   U7565 : OAI211_X1 port map( C1 => n7427, C2 => n6666, A => n6665, B => n6664
                           , ZN => n6667);
   U7566 : AOI211_X1 port map( C1 => n7322, C2 => n6669, A => n6668, B => n6667
                           , ZN => n6671);
   U7567 : OAI22_X1 port map( A1 => n6671, A2 => n6717, B1 => n6670, B2 => 
                           n7439, ZN => IF_ISAxN10950);
   U7568 : NAND2_X1 port map( A1 => n7400, A2 => n6672, ZN => n7342);
   U7569 : INV_X1 port map( A => n7342, ZN => n6714);
   U7570 : OR2_X1 port map( A1 => n6673, A2 => ashr_25xSHx3x, ZN => n6674);
   U7571 : AND2_X1 port map( A1 => n6675, A2 => n6674, ZN => n7330);
   U7572 : INV_X1 port map( A => n7330, ZN => n6679);
   U7573 : NAND3_X1 port map( A1 => n7342, A2 => n6677, A3 => n6676, ZN => 
                           n7350);
   U7574 : AOI222_X1 port map( A1 => n6679, A2 => n6734, B1 => n7350, B2 => 
                           n6678, C1 => n7368, C2 => DP_OP_719J14_125_1055xn83,
                           ZN => n6680);
   U7575 : INV_X1 port map( A => n6680, ZN => n6713);
   U7576 : AOI22_X1 port map( A1 => n6941, A2 => n6682, B1 => n6681, B2 => 
                           n6900, ZN => n6685);
   U7577 : INV_X1 port map( A => n6683, ZN => n6684);
   U7578 : AOI221_X1 port map( B1 => n6686, B2 => n7376, C1 => n6685, C2 => 
                           n7207, A => n6684, ZN => n6705);
   U7579 : OAI22_X1 port map( A1 => intadd_27xBx3x, A2 => n7227, B1 => n7118, 
                           B2 => n6687, ZN => n6692);
   U7580 : OAI221_X1 port map( B1 => n7470, B2 => n7389, C1 => n6693, C2 => 
                           n7115, A => n7387, ZN => n6688);
   U7581 : AOI221_X1 port map( B1 => n7410, B2 => intadd_27xBx3x, C1 => n7320, 
                           C2 => add_x_26xBx14x, A => n6688, ZN => n6690);
   U7582 : OAI22_X1 port map( A1 => intadd_27xAx3x, A2 => n6690, B1 => n7316, 
                           B2 => n6689, ZN => n6691);
   U7583 : AOI211_X1 port map( C1 => n7322, C2 => n6693, A => n6692, B => n6691
                           , ZN => n6703);
   U7584 : NOR2_X1 port map( A1 => n7470, A2 => ashr_25xAx14x, ZN => n6694);
   U7585 : AOI22_X1 port map( A1 => n6694, A2 => n7073, B1 => intadd_25xSUMx12x
                           , B2 => n7276, ZN => n6702);
   U7586 : AOI22_X1 port map( A1 => n7333, A2 => ashr_25xAx14x, B1 => 
                           ashr_25xAx13x, B2 => n7412, ZN => n6767);
   U7587 : AOI22_X1 port map( A1 => n7418, A2 => n6767, B1 => n6695, B2 => 
                           n7259, ZN => n6847);
   U7588 : AOI22_X1 port map( A1 => n6962, A2 => n6847, B1 => n6696, B2 => 
                           intadd_25xBx0x, ZN => n6966);
   U7589 : AND2_X1 port map( A1 => n6697, A2 => ashr_25xSHx3x, ZN => n6698);
   U7590 : AOI21_X1 port map( B1 => intadd_29xBx2x, B2 => n6966, A => n6698, ZN
                           => n7351);
   U7591 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx14x, B1 => 
                           ashr_25xAx13x, B2 => n7399, ZN => n6762);
   U7592 : AOI22_X1 port map( A1 => n7404, A2 => n6762, B1 => n6699, B2 => 
                           n7402, ZN => n6852);
   U7593 : AOI22_X1 port map( A1 => n6941, A2 => n6852, B1 => n6700, B2 => 
                           n6900, ZN => n6977);
   U7594 : AOI22_X1 port map( A1 => n7376, A2 => n6977, B1 => n6978, B2 => 
                           n7207, ZN => n7347);
   U7595 : AOI22_X1 port map( A1 => n7420, A2 => n7351, B1 => n7409, B2 => 
                           n7347, ZN => n6701);
   U7596 : NAND3_X1 port map( A1 => n6703, A2 => n6702, A3 => n6701, ZN => 
                           n6704);
   U7597 : NOR2_X1 port map( A1 => n6705, A2 => n6704, ZN => n6710);
   U7598 : OAI221_X1 port map( B1 => intadd_29xBx2x, B2 => n6708, C1 => 
                           ashr_25xSHx3x, C2 => n6707, A => n6706, ZN => n6709)
                           ;
   U7599 : OAI211_X1 port map( C1 => n6741, C2 => n6711, A => n6710, B => n6709
                           , ZN => n6712);
   U7600 : AOI211_X1 port map( C1 => n6715, C2 => n6714, A => n6713, B => n6712
                           , ZN => n6718);
   U7601 : OAI22_X1 port map( A1 => n6718, A2 => n6717, B1 => n6716, B2 => 
                           n7439, ZN => IF_ISAxN10951);
   U7602 : INV_X1 port map( A => n6719, ZN => n6721);
   U7603 : AOI221_X1 port map( B1 => n6722, B2 => ashr_25xSHx3x, C1 => n6721, 
                           C2 => intadd_29xBx2x, A => n6720, ZN => n6758);
   U7604 : NAND2_X1 port map( A1 => n7400, A2 => n6723, ZN => n7426);
   U7605 : AOI22_X1 port map( A1 => n7418, A2 => n6725, B1 => n6724, B2 => 
                           n7259, ZN => n6896);
   U7606 : AOI22_X1 port map( A1 => n6962, A2 => n6896, B1 => n6726, B2 => 
                           intadd_25xBx0x, ZN => n7017);
   U7607 : INV_X1 port map( A => n7001, ZN => n6727);
   U7608 : NOR2_X1 port map( A1 => n6727, A2 => intadd_29xBx2x, ZN => n6728);
   U7609 : AOI21_X1 port map( B1 => intadd_29xBx2x, B2 => n7017, A => n6728, ZN
                           => n7371);
   U7610 : OAI22_X1 port map( A1 => n6729, A2 => n7426, B1 => n7343, B2 => 
                           n7371, ZN => n6757);
   U7611 : AOI22_X1 port map( A1 => n7404, A2 => n6731, B1 => n6730, B2 => 
                           n7402, ZN => n6901);
   U7612 : AOI22_X1 port map( A1 => n6941, A2 => n6901, B1 => n6732, B2 => 
                           n6900, ZN => n7375);
   U7613 : NOR2_X1 port map( A1 => n7471, A2 => ashr_25xAx15x, ZN => n6733);
   U7614 : AOI22_X1 port map( A1 => n6733, A2 => n7073, B1 => intadd_25xSUMx13x
                           , B2 => n7276, ZN => n6736);
   U7615 : AOI22_X1 port map( A1 => n7394, A2 => n7372, B1 => n6734, B2 => 
                           n7413, ZN => n6735);
   U7616 : OAI211_X1 port map( C1 => n7375, C2 => n6967, A => n6736, B => n6735
                           , ZN => n6737);
   U7617 : AOI21_X1 port map( B1 => DP_OP_719J14_125_1055xn84, B2 => n7159, A 
                           => n6737, ZN => n6738);
   U7618 : INV_X1 port map( A => n6738, ZN => n6756);
   U7619 : OAI221_X1 port map( B1 => n7471, B2 => n7389, C1 => n6739, C2 => 
                           n7115, A => n7387, ZN => n6740);
   U7620 : AOI21_X1 port map( B1 => n7320, B2 => add_x_26xBx15x, A => n6740, ZN
                           => n6754);
   U7621 : INV_X1 port map( A => n6741, ZN => n6747);
   U7622 : OAI22_X1 port map( A1 => n6743, A2 => n7227, B1 => n7118, B2 => 
                           n6742, ZN => n6746);
   U7623 : OAI22_X1 port map( A1 => n6744, A2 => n7316, B1 => n7471, B2 => 
                           n7398, ZN => n6745);
   U7624 : AOI211_X1 port map( C1 => n7396, C2 => n6747, A => n6746, B => n6745
                           , ZN => n6753);
   U7625 : INV_X1 port map( A => n6748, ZN => n6749);
   U7626 : OAI221_X1 port map( B1 => n7376, B2 => n6750, C1 => n7207, C2 => 
                           n6749, A => n7192, ZN => n6751);
   U7627 : OAI21_X1 port map( B1 => n7046, B2 => n7353, A => n6751, ZN => n6752
                           );
   U7628 : OAI211_X1 port map( C1 => n6766, C2 => n6754, A => n6753, B => n6752
                           , ZN => n6755);
   U7629 : NOR4_X1 port map( A1 => n6758, A2 => n6757, A3 => n6756, A4 => n6755
                           , ZN => n6760);
   U7630 : OAI22_X1 port map( A1 => n6760, A2 => n7533, B1 => n6759, B2 => 
                           n7439, ZN => IF_ISAxN10952);
   U7631 : NAND2_X1 port map( A1 => n6761, A2 => n7309, ZN => n6764);
   U7632 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx16x, B1 => 
                           ashr_25xAx15x, B2 => n7267, ZN => n6851);
   U7633 : AOI22_X1 port map( A1 => n7404, A2 => n6851, B1 => n6762, B2 => 
                           n7402, ZN => n6940);
   U7634 : NAND2_X1 port map( A1 => n6940, A2 => n7311, ZN => n6763);
   U7635 : AND2_X1 port map( A1 => n6764, A2 => n6763, ZN => n7052);
   U7636 : INV_X1 port map( A => n7431, ZN => n6965);
   U7637 : OAI22_X1 port map( A1 => n7052, A2 => n6967, B1 => n6765, B2 => 
                           n6965, ZN => n6799);
   U7638 : AOI22_X1 port map( A1 => n7333, A2 => n6774, B1 => n6766, B2 => 
                           n7412, ZN => n6846);
   U7639 : INV_X1 port map( A => n6767, ZN => n6768);
   U7640 : AOI22_X1 port map( A1 => n7418, A2 => n6846, B1 => n6768, B2 => 
                           n7259, ZN => n6936);
   U7641 : INV_X1 port map( A => n6936, ZN => n6770);
   U7642 : AOI22_X1 port map( A1 => n6962, A2 => n6770, B1 => n6769, B2 => 
                           intadd_25xBx0x, ZN => n7038);
   U7643 : INV_X1 port map( A => n7018, ZN => n6850);
   U7644 : OAI22_X1 port map( A1 => n7038, A2 => n6850, B1 => n6771, B2 => 
                           n7314, ZN => n6798);
   U7645 : AOI22_X1 port map( A1 => n7320, A2 => add_x_26xBx16x, B1 => n7253, 
                           B2 => n6777, ZN => n6773);
   U7646 : OAI21_X1 port map( B1 => n6786, B2 => n7349, A => n7353, ZN => n6772
                           );
   U7647 : OAI221_X1 port map( B1 => n6774, B2 => n6773, C1 => n6774, C2 => 
                           n7387, A => n6772, ZN => n6797);
   U7648 : AOI22_X1 port map( A1 => n7276, A2 => intadd_25xSUMx14x, B1 => n7410
                           , B2 => n6775, ZN => n6793);
   U7649 : AOI21_X1 port map( B1 => n7331, B2 => n6789, A => n7329, ZN => n6785
                           );
   U7650 : AOI22_X1 port map( A1 => n7322, A2 => n6777, B1 => n6776, B2 => 
                           n7447, ZN => n6782);
   U7651 : INV_X1 port map( A => n6778, ZN => n6780);
   U7652 : OAI21_X1 port map( B1 => n6780, B2 => n6779, A => n7327, ZN => n6781
                           );
   U7653 : OAI211_X1 port map( C1 => n6783, C2 => n7227, A => n6782, B => n6781
                           , ZN => n6784);
   U7654 : AOI211_X1 port map( C1 => n7046, C2 => n6786, A => n6785, B => n6784
                           , ZN => n6792);
   U7655 : AOI22_X1 port map( A1 => n6788, A2 => n7352, B1 => n6787, B2 => 
                           n7348, ZN => n6791);
   U7656 : OR2_X1 port map( A1 => n6789, A2 => n7220, ZN => n6790);
   U7657 : NAND4_X1 port map( A1 => n6793, A2 => n6792, A3 => n6791, A4 => 
                           n6790, ZN => n6794);
   U7658 : AOI21_X1 port map( B1 => n7368, B2 => DP_OP_719J14_125_1055xn85, A 
                           => n6794, ZN => n6795);
   U7659 : INV_X1 port map( A => n6795, ZN => n6796);
   U7660 : NOR4_X1 port map( A1 => n6799, A2 => n6798, A3 => n6797, A4 => n6796
                           , ZN => n6801);
   U7661 : OAI22_X1 port map( A1 => n6801, A2 => n7533, B1 => n6800, B2 => 
                           n7439, ZN => IF_ISAxN10953);
   U7662 : AOI22_X1 port map( A1 => n6802, A2 => n7073, B1 => intadd_25xSUMx15x
                           , B2 => n7276, ZN => n6804);
   U7663 : AOI22_X1 port map( A1 => n7322, A2 => n6806, B1 => add_x_26xBx17x, 
                           B2 => n7380, ZN => n6803);
   U7664 : OAI211_X1 port map( C1 => n7118, C2 => n6805, A => n6804, B => n6803
                           , ZN => n6838);
   U7665 : OAI221_X1 port map( B1 => n7473, B2 => n7389, C1 => n6806, C2 => 
                           n7115, A => n7387, ZN => n6807);
   U7666 : AOI221_X1 port map( B1 => n7410, B2 => intadd_26xBx0x, C1 => n7320, 
                           C2 => add_x_26xBx17x, A => n6807, ZN => n6810);
   U7667 : INV_X1 port map( A => n6808, ZN => n6809);
   U7668 : OAI22_X1 port map( A1 => intadd_26xAx0x, A2 => n6810, B1 => n7316, 
                           B2 => n6809, ZN => n6837);
   U7669 : AOI22_X1 port map( A1 => n6962, A2 => n6813, B1 => n6812, B2 => 
                           n6811, ZN => n7112);
   U7670 : AOI22_X1 port map( A1 => n7431, A2 => n6814, B1 => n7018, B2 => 
                           n7112, ZN => n6817);
   U7671 : OAI21_X1 port map( B1 => n6815, B2 => n7349, A => n7353, ZN => n6816
                           );
   U7672 : OAI211_X1 port map( C1 => n7314, C2 => n6818, A => n6817, B => n6816
                           , ZN => n6836);
   U7673 : AND2_X1 port map( A1 => DP_OP_719J14_125_1055xn86, A2 => n7368, ZN 
                           => n6834);
   U7674 : INV_X1 port map( A => n7348, ZN => n7373);
   U7675 : OAI22_X1 port map( A1 => n7373, A2 => n6820, B1 => n7220, B2 => 
                           n6819, ZN => n6833);
   U7676 : OR2_X1 port map( A1 => n6821, A2 => n7309, ZN => n6824);
   U7677 : NAND2_X1 port map( A1 => n6822, A2 => n7309, ZN => n6823);
   U7678 : AND2_X1 port map( A1 => n6824, A2 => n6823, ZN => n7084);
   U7679 : INV_X1 port map( A => n7084, ZN => n6825);
   U7680 : NAND2_X1 port map( A1 => n7307, A2 => n6825, ZN => n6826);
   U7681 : NOR2_X1 port map( A1 => n7329, A2 => n7331, ZN => n7289);
   U7682 : INV_X1 port map( A => n7289, ZN => n7101);
   U7683 : OAI211_X1 port map( C1 => n7329, C2 => n6827, A => n6826, B => n7101
                           , ZN => n6832);
   U7684 : AOI22_X1 port map( A1 => n7046, A2 => n6829, B1 => n7352, B2 => 
                           n6828, ZN => n6830);
   U7685 : INV_X1 port map( A => n6830, ZN => n6831);
   U7686 : OR4_X1 port map( A1 => n6834, A2 => n6833, A3 => n6832, A4 => n6831,
                           ZN => n6835);
   U7687 : NOR4_X1 port map( A1 => n6838, A2 => n6837, A3 => n6836, A4 => n6835
                           , ZN => n6840);
   U7688 : OAI22_X1 port map( A1 => n6840, A2 => n7533, B1 => n6839, B2 => 
                           n7439, ZN => IF_ISAxN10954);
   U7689 : NAND2_X1 port map( A1 => n7192, A2 => n6841, ZN => n6842);
   U7690 : AOI22_X1 port map( A1 => n7166, A2 => n6843, B1 => n7353, B2 => 
                           n6842, ZN => n6844);
   U7691 : OAI21_X1 port map( B1 => n7373, B2 => n6845, A => n6844, ZN => n6876
                           );
   U7692 : AOI22_X1 port map( A1 => n7333, A2 => intadd_26xAx1x, B1 => 
                           intadd_26xAx0x, B2 => n7412, ZN => n6935);
   U7693 : AOI22_X1 port map( A1 => n7418, A2 => n6935, B1 => n6846, B2 => 
                           n7231, ZN => n6961);
   U7694 : INV_X1 port map( A => n6961, ZN => n6848);
   U7695 : AOI22_X1 port map( A1 => n6962, A2 => n6848, B1 => n6847, B2 => 
                           intadd_25xBx0x, ZN => n7136);
   U7696 : OAI22_X1 port map( A1 => n7136, A2 => n6850, B1 => n6849, B2 => 
                           n7314, ZN => n6875);
   U7697 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx18x, B1 => 
                           ashr_25xAx17x, B2 => n7267, ZN => n6939);
   U7698 : AOI22_X1 port map( A1 => n7404, A2 => n6939, B1 => n6851, B2 => 
                           n7402, ZN => n6964);
   U7699 : AOI22_X1 port map( A1 => n6941, A2 => n6964, B1 => n6852, B2 => 
                           n6900, ZN => n7125);
   U7700 : OAI22_X1 port map( A1 => n7125, A2 => n6967, B1 => n6853, B2 => 
                           n6965, ZN => n6874);
   U7701 : INV_X1 port map( A => intadd_25xSUMx16x, ZN => n6854);
   U7702 : OAI22_X1 port map( A1 => n6855, A2 => n7115, B1 => n6854, B2 => 
                           n7384, ZN => n6871);
   U7703 : AOI221_X1 port map( B1 => n7327, B2 => n7474, C1 => n7253, C2 => 
                           n6861, A => n7251, ZN => n6856);
   U7704 : OAI221_X1 port map( B1 => intadd_26xBx1x, B2 => n7386, C1 => 
                           add_x_26xBx18x, C2 => n7255, A => n6856, ZN => n6868
                           );
   U7705 : INV_X1 port map( A => n7352, ZN => n7370);
   U7706 : OAI22_X1 port map( A1 => n6858, A2 => n7427, B1 => n7370, B2 => 
                           n6857, ZN => n6867);
   U7707 : OAI22_X1 port map( A1 => intadd_26xBx1x, A2 => n7227, B1 => n7118, 
                           B2 => n6859, ZN => n6860);
   U7708 : AOI211_X1 port map( C1 => n7322, C2 => n6861, A => n6860, B => n7289
                           , ZN => n6865);
   U7709 : INV_X1 port map( A => n7329, ZN => n7174);
   U7710 : NOR2_X1 port map( A1 => intadd_26xBx1x, A2 => ashr_25xAx18x, ZN => 
                           n6862);
   U7711 : AOI22_X1 port map( A1 => n7174, A2 => n6863, B1 => n6862, B2 => 
                           n7410, ZN => n6864);
   U7712 : NAND2_X1 port map( A1 => n6865, A2 => n6864, ZN => n6866);
   U7713 : AOI211_X1 port map( C1 => n6868, C2 => ashr_25xAx18x, A => n6867, B 
                           => n6866, ZN => n6869);
   U7714 : INV_X1 port map( A => n6869, ZN => n6870);
   U7715 : AOI211_X1 port map( C1 => DP_OP_719J14_125_1055xn87, C2 => n7159, A 
                           => n6871, B => n6870, ZN => n6872);
   U7716 : INV_X1 port map( A => n6872, ZN => n6873);
   U7717 : NOR4_X1 port map( A1 => n6876, A2 => n6875, A3 => n6874, A4 => n6873
                           , ZN => n6878);
   U7718 : OAI22_X1 port map( A1 => n6878, A2 => n7533, B1 => n6877, B2 => 
                           n7439, ZN => IF_ISAxN10955);
   U7719 : AOI22_X1 port map( A1 => n7046, A2 => n6880, B1 => n7166, B2 => 
                           n6879, ZN => n6883);
   U7720 : OAI21_X1 port map( B1 => n6881, B2 => ashr_25xSHx4x, A => n7174, ZN 
                           => n6882);
   U7721 : OAI211_X1 port map( C1 => n6884, C2 => n7373, A => n6883, B => n6882
                           , ZN => n6915);
   U7722 : INV_X1 port map( A => n6885, ZN => n6886);
   U7723 : OAI22_X1 port map( A1 => n6887, A2 => n7397, B1 => n6886, B2 => 
                           n7316, ZN => n6914);
   U7724 : AOI22_X1 port map( A1 => n7322, A2 => n6888, B1 => add_x_26xBx19x, 
                           B2 => n7380, ZN => n6892);
   U7725 : AOI221_X1 port map( B1 => n7327, B2 => n7475, C1 => n7253, C2 => 
                           n6888, A => n7251, ZN => n6889);
   U7726 : OAI221_X1 port map( B1 => intadd_26xBx2x, B2 => n7386, C1 => 
                           add_x_26xBx19x, C2 => n7255, A => n6889, ZN => n6890
                           );
   U7727 : AOI22_X1 port map( A1 => n7276, A2 => intadd_25xSUMx17x, B1 => 
                           ashr_25xAx19x, B2 => n6890, ZN => n6891);
   U7728 : OAI211_X1 port map( C1 => n7118, C2 => n6893, A => n6892, B => n6891
                           , ZN => n6913);
   U7729 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn88, A2 => n7368, ZN 
                           => n6911);
   U7730 : AOI22_X1 port map( A1 => n7418, A2 => n6895, B1 => n6894, B2 => 
                           n7231, ZN => n7016);
   U7731 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n7016, B1 => n6896, 
                           B2 => intadd_25xBx0x, ZN => n7198);
   U7732 : AOI21_X1 port map( B1 => n7192, B2 => n6897, A => n7190, ZN => n6905
                           );
   U7733 : AOI22_X1 port map( A1 => n7404, A2 => n6899, B1 => n6898, B2 => 
                           n7402, ZN => n6999);
   U7734 : INV_X1 port map( A => n6999, ZN => n6902);
   U7735 : AOI22_X1 port map( A1 => n6941, A2 => n6902, B1 => n6901, B2 => 
                           n6900, ZN => n7195);
   U7736 : OAI22_X1 port map( A1 => n7195, A2 => n6967, B1 => n6903, B2 => 
                           n7314, ZN => n6904);
   U7737 : AOI211_X1 port map( C1 => n7018, C2 => n7198, A => n6905, B => n6904
                           , ZN => n6910);
   U7738 : INV_X1 port map( A => n6906, ZN => n6907);
   U7739 : AOI22_X1 port map( A1 => n7431, A2 => n6908, B1 => n7352, B2 => 
                           n6907, ZN => n6909);
   U7740 : NAND3_X1 port map( A1 => n6911, A2 => n6910, A3 => n6909, ZN => 
                           n6912);
   U7741 : NOR4_X1 port map( A1 => n6915, A2 => n6914, A3 => n6913, A4 => n6912
                           , ZN => n6917);
   U7742 : OAI22_X1 port map( A1 => n6917, A2 => n7533, B1 => n6916, B2 => 
                           n7439, ZN => IF_ISAxN10956);
   U7743 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn89, A2 => n7368, ZN 
                           => n6925);
   U7744 : AOI22_X1 port map( A1 => intadd_25xSUMx18x, A2 => n7276, B1 => n6918
                           , B2 => n7410, ZN => n6924);
   U7745 : INV_X1 port map( A => n6919, ZN => n6922);
   U7746 : INV_X1 port map( A => n6920, ZN => n6921);
   U7747 : AOI22_X1 port map( A1 => n7046, A2 => n6922, B1 => n7166, B2 => 
                           n6921, ZN => n6923);
   U7748 : NAND3_X1 port map( A1 => n6925, A2 => n6924, A3 => n6923, ZN => 
                           n6953);
   U7749 : OAI211_X1 port map( C1 => n7322, C2 => n7327, A => intadd_26xAx3x, B
                           => n6933, ZN => n6928);
   U7750 : AOI22_X1 port map( A1 => n6926, A2 => n7447, B1 => add_x_26xBx20x, 
                           B2 => n7380, ZN => n6927);
   U7751 : OAI211_X1 port map( C1 => n6930, C2 => n6929, A => n6928, B => n6927
                           , ZN => n6952);
   U7752 : OAI22_X1 port map( A1 => n6932, A2 => n7004, B1 => n6931, B2 => 
                           n7314, ZN => n6951);
   U7753 : OAI221_X1 port map( B1 => n7476, B2 => n7389, C1 => n6933, C2 => 
                           n7115, A => n7387, ZN => n6934);
   U7754 : AOI221_X1 port map( B1 => n7410, B2 => intadd_26xBx3x, C1 => n7320, 
                           C2 => add_x_26xBx20x, A => n6934, ZN => n6949);
   U7755 : AOI22_X1 port map( A1 => n7333, A2 => intadd_26xAx3x, B1 => 
                           intadd_26xAx2x, B2 => n7412, ZN => n6960);
   U7756 : AOI22_X1 port map( A1 => n7418, A2 => n6960, B1 => n6935, B2 => 
                           n7416, ZN => n7039);
   U7757 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n7039, B1 => n6936, 
                           B2 => intadd_25xBx0x, ZN => n7235);
   U7758 : AOI22_X1 port map( A1 => n7435, A2 => ashr_25xSHx4x, B1 => n6938, B2
                           => n6937, ZN => n6945);
   U7759 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx20x, B1 => 
                           ashr_25xAx19x, B2 => n7267, ZN => n6963);
   U7760 : AOI22_X1 port map( A1 => n7404, A2 => n6963, B1 => n6939, B2 => 
                           n7402, ZN => n7036);
   U7761 : AOI22_X1 port map( A1 => n6941, A2 => n7036, B1 => n6940, B2 => 
                           n7309, ZN => n7208);
   U7762 : INV_X1 port map( A => n6942, ZN => n6943);
   U7763 : OAI22_X1 port map( A1 => n7208, A2 => n6967, B1 => n6943, B2 => 
                           n6965, ZN => n6944);
   U7764 : AOI211_X1 port map( C1 => n7018, C2 => n7235, A => n6945, B => n6944
                           , ZN => n6948);
   U7765 : OAI21_X1 port map( B1 => n7349, B2 => n6946, A => n7353, ZN => n6947
                           );
   U7766 : OAI211_X1 port map( C1 => intadd_26xAx3x, C2 => n6949, A => n6948, B
                           => n6947, ZN => n6950);
   U7767 : NOR4_X1 port map( A1 => n6953, A2 => n6952, A3 => n6951, A4 => n6950
                           , ZN => n6955);
   U7768 : OAI22_X1 port map( A1 => n6955, A2 => n7533, B1 => n6954, B2 => 
                           n7439, ZN => IF_ISAxN10957);
   U7769 : AOI221_X1 port map( B1 => n7327, B2 => n7478, C1 => n7253, C2 => 
                           n6958, A => n7251, ZN => n6956);
   U7770 : OAI221_X1 port map( B1 => intadd_26xBx5x, B2 => n7386, C1 => 
                           add_x_26xBx22x, C2 => n7255, A => n6956, ZN => n6957
                           );
   U7771 : AOI22_X1 port map( A1 => n7276, A2 => intadd_25xSUMx20x, B1 => 
                           ashr_25xAx22x, B2 => n6957, ZN => n6973);
   U7772 : AOI22_X1 port map( A1 => n7166, A2 => n6959, B1 => n7322, B2 => 
                           n6958, ZN => n6972);
   U7773 : AOI22_X1 port map( A1 => n7333, A2 => intadd_26xAx5x, B1 => 
                           intadd_26xAx4x, B2 => n7412, ZN => n7037);
   U7774 : AOI22_X1 port map( A1 => n7418, A2 => n7037, B1 => n6960, B2 => 
                           n7416, ZN => n7133);
   U7775 : AOI22_X1 port map( A1 => n6962, A2 => n7133, B1 => n6961, B2 => 
                           intadd_25xBx0x, ZN => n7299);
   U7776 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx22x, B1 => 
                           ashr_25xAx21x, B2 => n7267, ZN => n7035);
   U7777 : AOI22_X1 port map( A1 => n7404, A2 => n7035, B1 => n6963, B2 => 
                           n7402, ZN => n7142);
   U7778 : AOI22_X1 port map( A1 => n7311, A2 => n7142, B1 => n6964, B2 => 
                           n7309, ZN => n7315);
   U7779 : OAI22_X1 port map( A1 => n7315, A2 => n6967, B1 => n6966, B2 => 
                           n6965, ZN => n6968);
   U7780 : AOI21_X1 port map( B1 => n7018, B2 => n7299, A => n6968, ZN => n6971
                           );
   U7781 : OAI21_X1 port map( B1 => n7349, B2 => n6969, A => n7353, ZN => n6970
                           );
   U7782 : NAND4_X1 port map( A1 => n6973, A2 => n6972, A3 => n6971, A4 => 
                           n6970, ZN => n6993);
   U7783 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn91, A2 => n7368, ZN 
                           => n6991);
   U7784 : INV_X1 port map( A => n6974, ZN => n6976);
   U7785 : OAI22_X1 port map( A1 => n6976, A2 => n7397, B1 => n6975, B2 => 
                           n7316, ZN => n6980);
   U7786 : OAI22_X1 port map( A1 => n6978, A2 => n7004, B1 => n6977, B2 => 
                           n7314, ZN => n6979);
   U7787 : AOI211_X1 port map( C1 => n7000, C2 => n6981, A => n6980, B => n6979
                           , ZN => n6990);
   U7788 : NAND2_X1 port map( A1 => n7046, A2 => n6982, ZN => n6986);
   U7789 : NOR2_X1 port map( A1 => n7118, A2 => n6983, ZN => n6984);
   U7790 : AOI21_X1 port map( B1 => add_x_26xBx22x, B2 => n7380, A => n6984, ZN
                           => n6985);
   U7791 : NAND2_X1 port map( A1 => n6986, A2 => n6985, ZN => n6987);
   U7792 : AOI211_X1 port map( C1 => n6988, C2 => n7174, A => n7289, B => n6987
                           , ZN => n6989);
   U7793 : NAND3_X1 port map( A1 => n6991, A2 => n6990, A3 => n6989, ZN => 
                           n6992);
   U7794 : OAI21_X1 port map( B1 => n6993, B2 => n6992, A => n7029, ZN => n6994
                           );
   U7795 : OAI21_X1 port map( B1 => n7439, B2 => n6995, A => n6994, ZN => 
                           IF_ISAxN10959);
   U7796 : AOI22_X1 port map( A1 => n7073, A2 => n6997, B1 => n6996, B2 => 
                           n7447, ZN => n7003);
   U7797 : AOI22_X1 port map( A1 => n7268, A2 => intadd_26xAx6x, B1 => 
                           intadd_26xAx5x, B2 => n7267, ZN => n7087);
   U7798 : AOI22_X1 port map( A1 => n7404, A2 => n7087, B1 => n6998, B2 => 
                           n7402, ZN => n7162);
   U7799 : AOI22_X1 port map( A1 => n7311, A2 => n7162, B1 => n6999, B2 => 
                           n7309, ZN => n7393);
   U7800 : AOI22_X1 port map( A1 => n7001, A2 => n7000, B1 => n7307, B2 => 
                           n7393, ZN => n7002);
   U7801 : OAI211_X1 port map( C1 => n7005, C2 => n7004, A => n7003, B => n7002
                           , ZN => n7031);
   U7802 : AOI22_X1 port map( A1 => intadd_25xSUMx21x, A2 => n7276, B1 => n7006
                           , B2 => n7410, ZN => n7007);
   U7803 : OAI21_X1 port map( B1 => n7008, B2 => n7220, A => n7007, ZN => n7027
                           );
   U7804 : AOI221_X1 port map( B1 => n7327, B2 => n7479, C1 => n7253, C2 => 
                           n7009, A => n7251, ZN => n7010);
   U7805 : OAI221_X1 port map( B1 => intadd_26xBx6x, B2 => n7386, C1 => 
                           add_x_26xBx23x, C2 => n7255, A => n7010, ZN => n7024
                           );
   U7806 : OAI22_X1 port map( A1 => n7427, A2 => n7011, B1 => n7227, B2 => 
                           intadd_26xBx6x, ZN => n7014);
   U7807 : OAI22_X1 port map( A1 => n7398, A2 => n7479, B1 => n7329, B2 => 
                           n7012, ZN => n7013);
   U7808 : OR3_X1 port map( A1 => n7014, A2 => n7289, A3 => n7013, ZN => n7023)
                           ;
   U7809 : AOI22_X1 port map( A1 => n7333, A2 => intadd_26xAx6x, B1 => 
                           intadd_26xAx5x, B2 => n7412, ZN => n7091);
   U7810 : AOI22_X1 port map( A1 => n7418, A2 => n7091, B1 => n7015, B2 => 
                           n7259, ZN => n7179);
   U7811 : AOI22_X1 port map( A1 => intadd_29xBx1x, A2 => n7179, B1 => n7016, 
                           B2 => intadd_25xBx0x, ZN => n7430);
   U7812 : AOI22_X1 port map( A1 => n7018, A2 => n7430, B1 => n7431, B2 => 
                           n7017, ZN => n7021);
   U7813 : OAI21_X1 port map( B1 => n7349, B2 => n7019, A => n7353, ZN => n7020
                           );
   U7814 : OAI211_X1 port map( C1 => n7375, C2 => n7314, A => n7021, B => n7020
                           , ZN => n7022);
   U7815 : AOI211_X1 port map( C1 => n7024, C2 => ashr_25xAx23x, A => n7023, B 
                           => n7022, ZN => n7025);
   U7816 : INV_X1 port map( A => n7025, ZN => n7026);
   U7817 : AOI211_X1 port map( C1 => DP_OP_719J14_125_1055xn92, C2 => n7159, A 
                           => n7027, B => n7026, ZN => n7028);
   U7818 : INV_X1 port map( A => n7028, ZN => n7030);
   U7819 : OAI21_X1 port map( B1 => n7031, B2 => n7030, A => n7029, ZN => n7032
                           );
   U7820 : OAI21_X1 port map( B1 => n7439, B2 => n7033, A => n7032, ZN => 
                           IF_ISAxN10960);
   U7821 : AOI21_X1 port map( B1 => n7192, B2 => n7034, A => n7190, ZN => n7070
                           );
   U7822 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx24x, B1 => 
                           ashr_25xAx23x, B2 => n7086, ZN => n7141);
   U7823 : AOI22_X1 port map( A1 => n7404, A2 => n7141, B1 => n7035, B2 => 
                           n7402, ZN => n7213);
   U7824 : AOI22_X1 port map( A1 => n7275, A2 => n7036, B1 => n7400, B2 => 
                           n7213, ZN => n7045);
   U7825 : OAI22_X1 port map( A1 => n7130, A2 => intadd_26xAx7x, B1 => 
                           intadd_26xAx6x, B2 => n7414, ZN => n7131);
   U7826 : AOI22_X1 port map( A1 => n7418, A2 => n7131, B1 => n7037, B2 => 
                           n7416, ZN => n7229);
   U7827 : OAI222_X1 port map( A1 => n7132, A2 => n7039, B1 => n7415, B2 => 
                           n7229, C1 => n7038, C2 => n7236, ZN => n7041);
   U7828 : AOI22_X1 port map( A1 => n7420, A2 => n7041, B1 => n7352, B2 => 
                           n7040, ZN => n7044);
   U7829 : NAND3_X1 port map( A1 => intadd_29xBx2x, A2 => n7166, A3 => n7042, 
                           ZN => n7043);
   U7830 : OAI211_X1 port map( C1 => n7045, C2 => n7206, A => n7044, B => n7043
                           , ZN => n7069);
   U7831 : NAND2_X1 port map( A1 => n7376, A2 => n7046, ZN => n7193);
   U7832 : OAI221_X1 port map( B1 => n7480, B2 => n7389, C1 => n7053, C2 => 
                           n7115, A => n7387, ZN => n7047);
   U7833 : AOI221_X1 port map( B1 => n7410, B2 => intadd_26xBx7x, C1 => n7320, 
                           C2 => add_x_26xBx24x, A => n7047, ZN => n7048);
   U7834 : OAI22_X1 port map( A1 => n7049, A2 => n7193, B1 => intadd_26xAx7x, 
                           B2 => n7048, ZN => n7068);
   U7835 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn93, A2 => n7368, ZN 
                           => n7066);
   U7836 : NOR2_X1 port map( A1 => n7480, A2 => ashr_25xAx24x, ZN => n7050);
   U7837 : AOI22_X1 port map( A1 => n7050, A2 => n7073, B1 => intadd_25xSUMx22x
                           , B2 => n7276, ZN => n7065);
   U7838 : AOI22_X1 port map( A1 => n7410, A2 => n7051, B1 => add_x_26xBx24x, 
                           B2 => n7380, ZN => n7063);
   U7839 : INV_X1 port map( A => n7052, ZN => n7059);
   U7840 : NAND2_X1 port map( A1 => n7322, A2 => n7053, ZN => n7057);
   U7841 : AOI22_X1 port map( A1 => n7348, A2 => n7055, B1 => n7054, B2 => 
                           n7447, ZN => n7056);
   U7842 : NAND2_X1 port map( A1 => n7057, A2 => n7056, ZN => n7058);
   U7843 : AOI21_X1 port map( B1 => n7394, B2 => n7059, A => n7058, ZN => n7062
                           );
   U7844 : NAND2_X1 port map( A1 => n7174, A2 => n7060, ZN => n7061);
   U7845 : AND4_X1 port map( A1 => n7063, A2 => n7062, A3 => n7101, A4 => n7061
                           , ZN => n7064);
   U7846 : NAND3_X1 port map( A1 => n7066, A2 => n7065, A3 => n7064, ZN => 
                           n7067);
   U7847 : NOR4_X1 port map( A1 => n7070, A2 => n7069, A3 => n7068, A4 => n7067
                           , ZN => n7072);
   U7848 : OAI22_X1 port map( A1 => n7072, A2 => n7533, B1 => n7071, B2 => 
                           n7439, ZN => IF_ISAxN10961);
   U7849 : AOI22_X1 port map( A1 => n7074, A2 => n7073, B1 => intadd_25xSUMx23x
                           , B2 => n7276, ZN => n7078);
   U7850 : OAI22_X1 port map( A1 => n7080, A2 => n7227, B1 => n7481, B2 => 
                           n7398, ZN => n7075);
   U7851 : AOI21_X1 port map( B1 => n7076, B2 => n7410, A => n7075, ZN => n7077
                           );
   U7852 : OAI211_X1 port map( C1 => n7118, C2 => n7079, A => n7078, B => n7077
                           , ZN => n7111);
   U7853 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn94, A2 => n7159, ZN 
                           => n7109);
   U7854 : OAI221_X1 port map( B1 => n7080, B2 => n7320, C1 => add_x_26xBx25x, 
                           C2 => n7127, A => ashr_25xAx25x, ZN => n7081);
   U7855 : OAI21_X1 port map( B1 => n7220, B2 => n7082, A => n7081, ZN => n7107
                           );
   U7856 : OAI22_X1 port map( A1 => n7084, A2 => n7314, B1 => n7083, B2 => 
                           n7193, ZN => n7106);
   U7857 : AOI21_X1 port map( B1 => n7192, B2 => n7085, A => n7190, ZN => n7105
                           );
   U7858 : AOI22_X1 port map( A1 => n7268, A2 => n7129, B1 => intadd_26xAx7x, 
                           B2 => n7086, ZN => n7161);
   U7859 : AOI22_X1 port map( A1 => n7404, A2 => n7161, B1 => n7087, B2 => 
                           n7402, ZN => n7274);
   U7860 : OAI22_X1 port map( A1 => n7088, A2 => n7406, B1 => n7274, B2 => 
                           n7269, ZN => n7090);
   U7861 : AOI22_X1 port map( A1 => n7409, A2 => n7090, B1 => n7352, B2 => 
                           n7089, ZN => n7103);
   U7862 : AOI22_X1 port map( A1 => n7333, A2 => ashr_25xAx25x, B1 => 
                           ashr_25xAx24x, B2 => n7412, ZN => n7178);
   U7863 : INV_X1 port map( A => n7178, ZN => n7092);
   U7864 : AOI22_X1 port map( A1 => n7418, A2 => n7092, B1 => n7091, B2 => 
                           n7259, ZN => n7258);
   U7865 : OAI22_X1 port map( A1 => n7093, A2 => n7132, B1 => n7258, B2 => 
                           n7415, ZN => n7095);
   U7866 : AOI22_X1 port map( A1 => n7420, A2 => n7095, B1 => n7348, B2 => 
                           n7094, ZN => n7102);
   U7867 : INV_X1 port map( A => n7096, ZN => n7099);
   U7868 : OAI221_X1 port map( B1 => n7481, B2 => n7389, C1 => n7097, C2 => 
                           n7115, A => n7387, ZN => n7098);
   U7869 : AOI22_X1 port map( A1 => n7174, A2 => n7099, B1 => n7098, B2 => 
                           ashr_25xAx25x, ZN => n7100);
   U7870 : NAND4_X1 port map( A1 => n7103, A2 => n7102, A3 => n7101, A4 => 
                           n7100, ZN => n7104);
   U7871 : NOR4_X1 port map( A1 => n7107, A2 => n7106, A3 => n7105, A4 => n7104
                           , ZN => n7108);
   U7872 : NAND2_X1 port map( A1 => n7109, A2 => n7108, ZN => n7110);
   U7873 : AOI211_X1 port map( C1 => n7431, C2 => n7112, A => n7111, B => n7110
                           , ZN => n7114);
   U7874 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(25), ZN => n7113);
   U7875 : OAI22_X1 port map( A1 => n7114, A2 => n7533, B1 => n7113, B2 => 
                           n7439, ZN => IF_ISAxN10962);
   U7876 : OAI221_X1 port map( B1 => n7482, B2 => n7389, C1 => n7120, C2 => 
                           n7115, A => n7387, ZN => n7116);
   U7877 : AOI221_X1 port map( B1 => n7410, B2 => n7126, C1 => n7320, C2 => 
                           add_x_26xBx26x, A => n7116, ZN => n7119);
   U7878 : OAI22_X1 port map( A1 => n7160, A2 => n7119, B1 => n7118, B2 => 
                           n7117, ZN => n7156);
   U7879 : OAI211_X1 port map( C1 => n7322, C2 => n7327, A => n7160, B => n7120
                           , ZN => n7123);
   U7880 : OAI21_X1 port map( B1 => n7349, B2 => n7121, A => n7353, ZN => n7122
                           );
   U7881 : OAI211_X1 port map( C1 => n7126, C2 => n7227, A => n7123, B => n7122
                           , ZN => n7155);
   U7882 : OAI22_X1 port map( A1 => n7125, A2 => n7314, B1 => n7124, B2 => 
                           n7193, ZN => n7154);
   U7883 : NOR2_X1 port map( A1 => n7126, A2 => ashr_25xAx26x, ZN => n7128);
   U7884 : AOI22_X1 port map( A1 => intadd_25xSUMx24x, A2 => n7276, B1 => n7128
                           , B2 => n7127, ZN => n7150);
   U7885 : OAI22_X1 port map( A1 => n7130, A2 => n7160, B1 => n7129, B2 => 
                           n7414, ZN => n7230);
   U7886 : OAI22_X1 port map( A1 => n7231, A2 => n7230, B1 => n7131, B2 => 
                           n7418, ZN => n7338);
   U7887 : OAI22_X1 port map( A1 => n7338, A2 => n7415, B1 => n7133, B2 => 
                           n7132, ZN => n7134);
   U7888 : AOI22_X1 port map( A1 => n7174, A2 => n7135, B1 => n7420, B2 => 
                           n7134, ZN => n7149);
   U7889 : INV_X1 port map( A => n7136, ZN => n7137);
   U7890 : AOI21_X1 port map( B1 => n7431, B2 => n7137, A => n7289, ZN => n7148
                           );
   U7891 : AOI22_X1 port map( A1 => n7352, A2 => n7139, B1 => n7348, B2 => 
                           n7138, ZN => n7140);
   U7892 : INV_X1 port map( A => n7140, ZN => n7146);
   U7893 : AOI22_X1 port map( A1 => n7268, A2 => ashr_25xAx26x, B1 => 
                           ashr_25xAx25x, B2 => n7399, ZN => n7210);
   U7894 : AOI22_X1 port map( A1 => n7404, A2 => n7210, B1 => n7141, B2 => 
                           n7402, ZN => n7310);
   U7895 : AOI22_X1 port map( A1 => n7275, A2 => n7142, B1 => n7400, B2 => 
                           n7310, ZN => n7144);
   U7896 : OAI22_X1 port map( A1 => n7144, A2 => n7206, B1 => n7220, B2 => 
                           n7143, ZN => n7145);
   U7897 : NOR2_X1 port map( A1 => n7146, A2 => n7145, ZN => n7147);
   U7898 : NAND4_X1 port map( A1 => n7150, A2 => n7149, A3 => n7148, A4 => 
                           n7147, ZN => n7151);
   U7899 : AOI21_X1 port map( B1 => DP_OP_719J14_125_1055xn95, B2 => n7159, A 
                           => n7151, ZN => n7152);
   U7900 : INV_X1 port map( A => n7152, ZN => n7153);
   U7901 : NOR4_X1 port map( A1 => n7156, A2 => n7155, A3 => n7154, A4 => n7153
                           , ZN => n7158);
   U7902 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(26), ZN => n7157);
   U7903 : OAI22_X1 port map( A1 => n7158, A2 => n7533, B1 => n7157, B2 => 
                           n7439, ZN => IF_ISAxN10963);
   U7904 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn96, A2 => n7159, ZN 
                           => n7177);
   U7905 : AOI22_X1 port map( A1 => n7209, A2 => n7184, B1 => n7160, B2 => 
                           n7399, ZN => n7270);
   U7906 : AOI22_X1 port map( A1 => n7404, A2 => n7270, B1 => n7161, B2 => 
                           n7402, ZN => n7407);
   U7907 : OAI22_X1 port map( A1 => n7162, A2 => n7406, B1 => n7407, B2 => 
                           n7269, ZN => n7164);
   U7908 : AOI22_X1 port map( A1 => n7409, A2 => n7164, B1 => n7352, B2 => 
                           n7163, ZN => n7176);
   U7909 : INV_X1 port map( A => n7165, ZN => n7173);
   U7910 : AOI22_X1 port map( A1 => n7167, A2 => n7166, B1 => add_x_26xBx27x, 
                           B2 => n7380, ZN => n7171);
   U7911 : OAI22_X1 port map( A1 => n7483, A2 => n7389, B1 => n7168, B2 => 
                           n7386, ZN => n7169);
   U7912 : OAI21_X1 port map( B1 => n7251, B2 => n7169, A => ashr_25xAx27x, ZN 
                           => n7170);
   U7913 : OAI211_X1 port map( C1 => n7398, C2 => n7483, A => n7171, B => n7170
                           , ZN => n7172);
   U7914 : AOI211_X1 port map( C1 => n7174, C2 => n7173, A => n7289, B => n7172
                           , ZN => n7175);
   U7915 : NAND3_X1 port map( A1 => n7177, A2 => n7176, A3 => n7175, ZN => 
                           n7203);
   U7916 : AOI22_X1 port map( A1 => n7333, A2 => ashr_25xAx27x, B1 => 
                           ashr_25xAx26x, B2 => n7412, ZN => n7260);
   U7917 : AOI22_X1 port map( A1 => n7418, A2 => n7260, B1 => n7178, B2 => 
                           n7231, ZN => n7421);
   U7918 : INV_X1 port map( A => n7179, ZN => n7180);
   U7919 : AOI22_X1 port map( A1 => n7341, A2 => n7421, B1 => n7422, B2 => 
                           n7180, ZN => n7201);
   U7920 : OAI22_X1 port map( A1 => n7182, A2 => n7316, B1 => n7181, B2 => 
                           n7397, ZN => n7188);
   U7921 : NAND2_X1 port map( A1 => n7184, A2 => n7183, ZN => n7186);
   U7922 : OAI22_X1 port map( A1 => n7186, A2 => n7397, B1 => n7185, B2 => 
                           n7384, ZN => n7187);
   U7923 : AOI211_X1 port map( C1 => n7348, C2 => n7189, A => n7188, B => n7187
                           , ZN => n7200);
   U7924 : AOI21_X1 port map( B1 => n7192, B2 => n7191, A => n7190, ZN => n7197
                           );
   U7925 : OAI22_X1 port map( A1 => n7195, A2 => n7314, B1 => n7194, B2 => 
                           n7193, ZN => n7196);
   U7926 : AOI211_X1 port map( C1 => n7431, C2 => n7198, A => n7197, B => n7196
                           , ZN => n7199);
   U7927 : OAI211_X1 port map( C1 => n7201, C2 => n7343, A => n7200, B => n7199
                           , ZN => n7202);
   U7928 : AOI211_X1 port map( C1 => n7204, C2 => n7447, A => n7203, B => n7202
                           , ZN => n7205);
   U7929 : OAI22_X1 port map( A1 => n7205, A2 => n7533, B1 => n3646, B2 => 
                           n7439, ZN => IF_ISAxN10964);
   U7930 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn97, A2 => n7368, ZN 
                           => n7219);
   U7931 : AOI21_X1 port map( B1 => n7208, B2 => n7207, A => n7206, ZN => n7212
                           );
   U7932 : AOI22_X1 port map( A1 => n7209, A2 => ashr_25xAx28x, B1 => 
                           ashr_25xAx27x, B2 => n7267, ZN => n7301);
   U7933 : OAI221_X1 port map( B1 => n7304, B2 => n7210, C1 => n7402, C2 => 
                           n7301, A => n7400, ZN => n7211);
   U7934 : OAI211_X1 port map( C1 => n7406, C2 => n7213, A => n7212, B => n7211
                           , ZN => n7218);
   U7935 : INV_X1 port map( A => n7214, ZN => n7215);
   U7936 : AOI22_X1 port map( A1 => n7348, A2 => n7216, B1 => n7352, B2 => 
                           n7215, ZN => n7217);
   U7937 : NAND3_X1 port map( A1 => n7219, A2 => n7218, A3 => n7217, ZN => 
                           n7247);
   U7938 : NOR2_X1 port map( A1 => n7415, A2 => n7220, ZN => n7395);
   U7939 : INV_X1 port map( A => n7395, ZN => n7285);
   U7940 : AOI21_X1 port map( B1 => n7331, B2 => n7221, A => n7329, ZN => n7226
                           );
   U7941 : OAI221_X1 port map( B1 => n7484, B2 => n7389, C1 => n7242, C2 => 
                           n7397, A => n7387, ZN => n7222);
   U7942 : AOI221_X1 port map( B1 => n7410, B2 => intadd_28xBx0x, C1 => n7320, 
                           C2 => add_x_26xBx28x, A => n7222, ZN => n7224);
   U7943 : NAND2_X1 port map( A1 => intadd_28xAx0x, A2 => n7242, ZN => n7223);
   U7944 : OAI22_X1 port map( A1 => intadd_28xAx0x, A2 => n7224, B1 => n7397, 
                           B2 => n7223, ZN => n7225);
   U7945 : AOI211_X1 port map( C1 => n7276, C2 => intadd_25xSUMx26x, A => n7226
                           , B => n7225, ZN => n7244);
   U7946 : AOI221_X1 port map( B1 => ashr_25xAx28x, B2 => n7227, C1 => n7316, 
                           C2 => n7227, A => intadd_28xBx0x, ZN => n7241);
   U7947 : OAI21_X1 port map( B1 => n7349, B2 => n7228, A => n7353, ZN => n7238
                           );
   U7948 : AOI21_X1 port map( B1 => n7422, B2 => n7229, A => n7343, ZN => n7234
                           );
   U7949 : INV_X1 port map( A => n7230, ZN => n7232);
   U7950 : AOI22_X1 port map( A1 => n7333, A2 => ashr_25xAx28x, B1 => 
                           ashr_25xAx27x, B2 => n7412, ZN => n7332);
   U7951 : OAI221_X1 port map( B1 => n7418, B2 => n7232, C1 => n7231, C2 => 
                           n7332, A => n7341, ZN => n7233);
   U7952 : OAI211_X1 port map( C1 => n7236, C2 => n7235, A => n7234, B => n7233
                           , ZN => n7237);
   U7953 : OAI211_X1 port map( C1 => n7239, C2 => n7427, A => n7238, B => n7237
                           , ZN => n7240);
   U7954 : AOI211_X1 port map( C1 => n7322, C2 => n7242, A => n7241, B => n7240
                           , ZN => n7243);
   U7955 : OAI211_X1 port map( C1 => n7245, C2 => n7285, A => n7244, B => n7243
                           , ZN => n7246);
   U7956 : AOI211_X1 port map( C1 => n7248, C2 => n7447, A => n7247, B => n7246
                           , ZN => n7250);
   U7957 : OAI22_X1 port map( A1 => n7250, A2 => n7533, B1 => n7249, B2 => 
                           n7439, ZN => IF_ISAxN10965);
   U7958 : NAND2_X1 port map( A1 => intadd_28xAx1x, A2 => n7252, ZN => n7266);
   U7959 : AOI221_X1 port map( B1 => n7327, B2 => n7485, C1 => n7253, C2 => 
                           n7252, A => n7251, ZN => n7254);
   U7960 : OAI221_X1 port map( B1 => intadd_28xBx1x, B2 => n7386, C1 => 
                           add_x_26xBx29x, C2 => n7255, A => n7254, ZN => n7256
                           );
   U7961 : AOI22_X1 port map( A1 => n7410, A2 => n7257, B1 => ashr_25xAx29x, B2
                           => n7256, ZN => n7265);
   U7962 : AOI21_X1 port map( B1 => n7422, B2 => n7258, A => n7343, ZN => n7262
                           );
   U7963 : AOI22_X1 port map( A1 => n7333, A2 => ashr_25xAx29x, B1 => 
                           ashr_25xAx28x, B2 => n7130, ZN => n7417);
   U7964 : OAI221_X1 port map( B1 => n7418, B2 => n7260, C1 => n7259, C2 => 
                           n7417, A => n7341, ZN => n7261);
   U7965 : OAI211_X1 port map( C1 => intadd_29xBx2x, C2 => n7263, A => n7262, B
                           => n7261, ZN => n7264);
   U7966 : OAI211_X1 port map( C1 => n7397, C2 => n7266, A => n7265, B => n7264
                           , ZN => n7295);
   U7967 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn98, A2 => n7368, ZN 
                           => n7293);
   U7968 : AOI22_X1 port map( A1 => n7268, A2 => intadd_28xAx1x, B1 => 
                           intadd_28xAx0x, B2 => n7267, ZN => n7403);
   U7969 : AOI221_X1 port map( B1 => n7403, B2 => n7304, C1 => n7270, C2 => 
                           n5711, A => n7269, ZN => n7273);
   U7970 : OAI21_X1 port map( B1 => n7376, B2 => n7271, A => n7409, ZN => n7272
                           );
   U7971 : AOI211_X1 port map( C1 => n7275, C2 => n7274, A => n7273, B => n7272
                           , ZN => n7281);
   U7972 : AOI22_X1 port map( A1 => intadd_25xSUMx27x, A2 => n7276, B1 => 
                           add_x_26xBx29x, B2 => n7380, ZN => n7279);
   U7973 : OAI21_X1 port map( B1 => n7349, B2 => n7277, A => n7353, ZN => n7278
                           );
   U7974 : OAI211_X1 port map( C1 => n7485, C2 => n7398, A => n7279, B => n7278
                           , ZN => n7280);
   U7975 : AOI211_X1 port map( C1 => n7348, C2 => n7282, A => n7281, B => n7280
                           , ZN => n7292);
   U7976 : OAI22_X1 port map( A1 => n7427, A2 => n7284, B1 => n7370, B2 => 
                           n7283, ZN => n7290);
   U7977 : OAI22_X1 port map( A1 => n7329, A2 => n7287, B1 => n7286, B2 => 
                           n7285, ZN => n7288);
   U7978 : NOR3_X1 port map( A1 => n7290, A2 => n7289, A3 => n7288, ZN => n7291
                           );
   U7979 : NAND3_X1 port map( A1 => n7293, A2 => n7292, A3 => n7291, ZN => 
                           n7294);
   U7980 : AOI211_X1 port map( C1 => n7296, C2 => n7447, A => n7295, B => n7294
                           , ZN => n7298);
   U7981 : INV_X1 port map( A => fromMemoryPortxLOADEDDATAx(29), ZN => n7297);
   U7982 : OAI22_X1 port map( A1 => n7298, A2 => n7533, B1 => n7297, B2 => 
                           n7439, ZN => IF_ISAxN10966);
   U7983 : AOI22_X1 port map( A1 => n7395, A2 => n7300, B1 => n7431, B2 => 
                           n7299, ZN => n7313);
   U7984 : INV_X1 port map( A => n7301, ZN => n7306);
   U7985 : NOR2_X1 port map( A1 => n7399, A2 => ashr_25xAx30x, ZN => n7303);
   U7986 : NOR2_X1 port map( A1 => n7209, A2 => ashr_25xAx29x, ZN => n7302);
   U7987 : NOR2_X1 port map( A1 => n7303, A2 => n7302, ZN => n7305);
   U7988 : MUX2_X1 port map( A => n7306, B => n7305, S => n7304, Z => n7308);
   U7989 : OAI221_X1 port map( B1 => n7311, B2 => n7310, C1 => n7309, C2 => 
                           n7308, A => n7307, ZN => n7312);
   U7990 : OAI211_X1 port map( C1 => n7315, C2 => n7314, A => n7313, B => n7312
                           , ZN => n7360);
   U7991 : NAND2_X1 port map( A1 => DP_OP_719J14_125_1055xn99, A2 => n7368, ZN 
                           => n7358);
   U7992 : INV_X1 port map( A => intadd_25xSUMx28x, ZN => n7318);
   U7993 : OAI22_X1 port map( A1 => n7318, A2 => n7384, B1 => n7317, B2 => 
                           n7316, ZN => n7326);
   U7994 : OAI221_X1 port map( B1 => n7487, B2 => n7389, C1 => n7321, C2 => 
                           n7397, A => n7387, ZN => n7319);
   U7995 : AOI221_X1 port map( B1 => n7410, B2 => intadd_28xBx2x, C1 => n7320, 
                           C2 => add_x_26xBx30x, A => n7319, ZN => n7324);
   U7996 : AOI22_X1 port map( A1 => n7322, A2 => n7321, B1 => add_x_26xBx30x, 
                           B2 => n7380, ZN => n7323);
   U7997 : OAI21_X1 port map( B1 => intadd_28xAx2x, B2 => n7324, A => n7323, ZN
                           => n7325);
   U7998 : AOI211_X1 port map( C1 => n7328, C2 => n7327, A => n7326, B => n7325
                           , ZN => n7357);
   U7999 : AOI21_X1 port map( B1 => n7331, B2 => n7330, A => n7329, ZN => n7346
                           );
   U8000 : INV_X1 port map( A => n7332, ZN => n7337);
   U8001 : NOR2_X1 port map( A1 => ashr_25xAx30x, A2 => n7130, ZN => n7335);
   U8002 : NOR2_X1 port map( A1 => n7333, A2 => ashr_25xAx29x, ZN => n7334);
   U8003 : NOR2_X1 port map( A1 => n7335, A2 => n7334, ZN => n7336);
   U8004 : MUX2_X1 port map( A => n7337, B => n7336, S => n7418, Z => n7340);
   U8005 : INV_X1 port map( A => n7338, ZN => n7339);
   U8006 : AOI22_X1 port map( A1 => n7341, A2 => n7340, B1 => n7422, B2 => 
                           n7339, ZN => n7344);
   U8007 : OAI22_X1 port map( A1 => n7344, A2 => n7343, B1 => n7427, B2 => 
                           n7342, ZN => n7345);
   U8008 : AOI211_X1 port map( C1 => n7348, C2 => n7347, A => n7346, B => n7345
                           , ZN => n7356);
   U8009 : OR2_X1 port map( A1 => n7350, A2 => n7349, ZN => n7354);
   U8010 : AOI22_X1 port map( A1 => n7354, A2 => n7353, B1 => n7352, B2 => 
                           n7351, ZN => n7355);
   U8011 : NAND4_X1 port map( A1 => n7358, A2 => n7357, A3 => n7356, A4 => 
                           n7355, ZN => n7359);
   U8012 : AOI211_X1 port map( C1 => n7361, C2 => n7447, A => n7360, B => n7359
                           , ZN => n7363);
   U8013 : OAI22_X1 port map( A1 => n7363, A2 => n7533, B1 => n7362, B2 => 
                           n7439, ZN => IF_ISAxN10967);
   U8014 : OAI21_X1 port map( B1 => n7364, B2 => n7489, A => n7392, ZN => n7365
                           );
   U8015 : XOR2_X1 port map( A => n7550, B => n7365, Z => n7366);
   U8016 : XOR2_X1 port map( A => n7366, B => n7413, Z => n7367);
   U8017 : XOR2_X1 port map( A => DP_OP_719J14_125_1055xn2, B => n7367, Z => 
                           n7369);
   U8018 : NAND2_X1 port map( A1 => n7369, A2 => n7368, ZN => n7382);
   U8019 : NOR2_X1 port map( A1 => n7371, A2 => n7370, ZN => n7378);
   U8020 : NOR2_X1 port map( A1 => n7372, A2 => n7376, ZN => n7374);
   U8021 : AOI211_X1 port map( C1 => n7376, C2 => n7375, A => n7374, B => n7373
                           , ZN => n7377);
   U8022 : AOI211_X1 port map( C1 => n7380, C2 => n7379, A => n7378, B => n7377
                           , ZN => n7381);
   U8023 : OAI211_X1 port map( C1 => n7384, C2 => n7383, A => n7382, B => n7381
                           , ZN => n7437);
   U8024 : OAI21_X1 port map( B1 => n7392, B2 => n7386, A => n7385, ZN => n7391
                           );
   U8025 : OAI221_X1 port map( B1 => n7489, B2 => n7389, C1 => n7388, C2 => 
                           n7397, A => n7387, ZN => n7390);
   U8026 : AOI211_X1 port map( C1 => n7410, C2 => n7392, A => n7391, B => n7390
                           , ZN => n7434);
   U8027 : AOI22_X1 port map( A1 => n7396, A2 => n7395, B1 => n7394, B2 => 
                           n7393, ZN => n7433);
   U8028 : AOI211_X1 port map( C1 => n7398, C2 => n7397, A => n7413, B => n7489
                           , ZN => n7429);
   U8029 : AOI22_X1 port map( A1 => n7209, A2 => n7435, B1 => intadd_28xAx2x, 
                           B2 => n7399, ZN => n7401);
   U8030 : OAI221_X1 port map( B1 => n7404, B2 => n7403, C1 => n7402, C2 => 
                           n7401, A => n7400, ZN => n7405);
   U8031 : OAI21_X1 port map( B1 => n7407, B2 => n7406, A => n7405, ZN => n7408
                           );
   U8032 : AOI22_X1 port map( A1 => n7411, A2 => n7410, B1 => n7409, B2 => 
                           n7408, ZN => n7425);
   U8033 : AOI22_X1 port map( A1 => n7414, A2 => n7413, B1 => ashr_25xAx30x, B2
                           => n7412, ZN => n7419);
   U8034 : AOI221_X1 port map( B1 => n7419, B2 => n7418, C1 => n7417, C2 => 
                           n7416, A => n7415, ZN => n7423);
   U8035 : OAI221_X1 port map( B1 => n7423, B2 => n7422, C1 => n7423, C2 => 
                           n7421, A => n7420, ZN => n7424);
   U8036 : OAI211_X1 port map( C1 => n7427, C2 => n7426, A => n7425, B => n7424
                           , ZN => n7428);
   U8037 : AOI211_X1 port map( C1 => n7431, C2 => n7430, A => n7429, B => n7428
                           , ZN => n7432);
   U8038 : OAI211_X1 port map( C1 => n7435, C2 => n7434, A => n7433, B => n7432
                           , ZN => n7436);
   U8039 : AOI211_X1 port map( C1 => n7438, C2 => n7447, A => n7437, B => n7436
                           , ZN => n7441);
   U8040 : OAI22_X1 port map( A1 => n7441, A2 => n7533, B1 => n7440, B2 => 
                           n7439, ZN => IF_ISAxN10968);
   U8041 : NOR2_X1 port map( A1 => rst, A2 => n7442, ZN => IF_ISAxN10970);
   U8042 : NOR2_X1 port map( A1 => rst, A2 => n7443, ZN => IF_ISAxN10971);
   U8043 : AND2_X1 port map( A1 => n7509, A2 => fromMemoryPortxLOADEDDATAx(9), 
                           ZN => IF_ISAxN10972);
   U8044 : AND2_X1 port map( A1 => n7509, A2 => fromMemoryPortxLOADEDDATAx(10),
                           ZN => IF_ISAxN10973);
   U8045 : AND2_X1 port map( A1 => n7523, A2 => fromMemoryPortxLOADEDDATAx(11),
                           ZN => IF_ISAxN10974);
   U8046 : NAND3_X1 port map( A1 => n7538, A2 => n7535, A3 => n7455, ZN => 
                           n7492);
   U8047 : NOR2_X1 port map( A1 => fromMemoryPortxLOADEDDATAx(2), A2 => 
                           fromMemoryPortxLOADEDDATAx(4), ZN => n7451);
   U8048 : INV_X1 port map( A => n7492, ZN => n7450);
   U8049 : NOR3_X1 port map( A1 => n7446, A2 => n7445, A3 => n7444, ZN => n7448
                           );
   U8050 : NAND2_X1 port map( A1 => n7448, A2 => n7447, ZN => n7449);
   U8051 : NAND2_X1 port map( A1 => n7450, A2 => n7449, ZN => n7491);
   U8052 : NOR2_X1 port map( A1 => n7451, A2 => n7491, ZN => n7456);
   U8053 : NOR2_X1 port map( A1 => rst, A2 => n7456, ZN => n7527);
   U8054 : OAI21_X1 port map( B1 => n7452, B2 => n7492, A => n7527, ZN => 
                           IF_ISAxN10969);
   U8055 : INV_X1 port map( A => n7453, ZN => n7454);
   U8056 : AOI21_X1 port map( B1 => n7455, B2 => n7454, A => rst, ZN => n7493);
   U8057 : INV_X1 port map( A => n7456, ZN => n7532);
   U8058 : OAI211_X1 port map( C1 => n7457, C2 => n7492, A => n7493, B => n7532
                           , ZN => IF_ISAxN10902);
   U8059 : NAND2_X1 port map( A1 => n7458, A2 => IF_ISAxsection_0_port, ZN => 
                           n7459);
   U8060 : NAND3_X1 port map( A1 => n7460, A2 => n7493, A3 => n7459, ZN => 
                           n7488);
   U8061 : CLKBUF_X1 port map( A => n7488, Z => n7486);
   U8062 : NOR2_X1 port map( A1 => n7461, A2 => n7486, ZN => IF_ISAxN10842);
   U8063 : NOR2_X1 port map( A1 => n7462, A2 => n7486, ZN => IF_ISAxN10843);
   U8064 : NOR2_X1 port map( A1 => n7463, A2 => n7486, ZN => IF_ISAxN10844);
   U8065 : NOR2_X1 port map( A1 => n7464, A2 => n7486, ZN => IF_ISAxN10845);
   U8066 : NOR2_X1 port map( A1 => n7465, A2 => n7486, ZN => IF_ISAxN10846);
   U8067 : NOR2_X1 port map( A1 => n7466, A2 => n7486, ZN => IF_ISAxN10847);
   U8068 : NOR2_X1 port map( A1 => n7467, A2 => n7486, ZN => IF_ISAxN10848);
   U8069 : NOR2_X1 port map( A1 => n7468, A2 => n7486, ZN => IF_ISAxN10849);
   U8070 : NOR2_X1 port map( A1 => n7469, A2 => n7486, ZN => IF_ISAxN10850);
   U8071 : NOR2_X1 port map( A1 => n7470, A2 => n7486, ZN => IF_ISAxN10851);
   U8072 : NOR2_X1 port map( A1 => n7471, A2 => n7486, ZN => IF_ISAxN10852);
   U8073 : NOR2_X1 port map( A1 => n7472, A2 => n7486, ZN => IF_ISAxN10853);
   U8074 : NOR2_X1 port map( A1 => n7473, A2 => n7488, ZN => IF_ISAxN10854);
   U8075 : NOR2_X1 port map( A1 => n7474, A2 => n7488, ZN => IF_ISAxN10855);
   U8076 : NOR2_X1 port map( A1 => n7475, A2 => n7488, ZN => IF_ISAxN10856);
   U8077 : NOR2_X1 port map( A1 => n7476, A2 => n7488, ZN => IF_ISAxN10857);
   U8078 : NOR2_X1 port map( A1 => n7477, A2 => n7488, ZN => IF_ISAxN10858);
   U8079 : NOR2_X1 port map( A1 => n7478, A2 => n7488, ZN => IF_ISAxN10859);
   U8080 : NOR2_X1 port map( A1 => n7479, A2 => n7488, ZN => IF_ISAxN10860);
   U8081 : NOR2_X1 port map( A1 => n7480, A2 => n7488, ZN => IF_ISAxN10861);
   U8082 : NOR2_X1 port map( A1 => n7481, A2 => n7488, ZN => IF_ISAxN10862);
   U8083 : NOR2_X1 port map( A1 => n7482, A2 => n7488, ZN => IF_ISAxN10863);
   U8084 : NOR2_X1 port map( A1 => n7483, A2 => n7488, ZN => IF_ISAxN10864);
   U8085 : NOR2_X1 port map( A1 => n7484, A2 => n7486, ZN => IF_ISAxN10865);
   U8086 : NOR2_X1 port map( A1 => n7485, A2 => n7488, ZN => IF_ISAxN10866);
   U8087 : NOR2_X1 port map( A1 => n7487, A2 => n7486, ZN => IF_ISAxN10867);
   U8088 : NOR2_X1 port map( A1 => n7489, A2 => n7488, ZN => IF_ISAxN10868);
   U8089 : OAI21_X1 port map( B1 => n7490, B2 => n7492, A => n7493, ZN => 
                           IF_ISAxN10832);
   U8090 : NAND2_X1 port map( A1 => n7493, A2 => n7491, ZN => IF_ISAxN10869);
   U8091 : OAI21_X1 port map( B1 => n7538, B2 => n7535, A => 
                           toMemoryPort_sync_port, ZN => n7494);
   U8092 : OAI211_X1 port map( C1 => IF_ISAxsection_0_port, C2 => n7494, A => 
                           n7493, B => n7492, ZN => IF_ISAxN10829);
   U8093 : NAND2_X1 port map( A1 => toRegsPortxDSTxx3x, A2 => 
                           toRegsPortxDSTxx2x, ZN => n7496);
   U8094 : NOR2_X1 port map( A1 => n7534, A2 => n7496, ZN => n7508);
   U8095 : INV_X1 port map( A => n7508, ZN => n7495);
   U8096 : NAND2_X1 port map( A1 => toRegsPortxDSTxx0x, A2 => 
                           toRegsPortxDSTxx4x, ZN => n7506);
   U8097 : OR2_X1 port map( A1 => n7540, A2 => n7506, ZN => n7497);
   U8098 : OAI21_X1 port map( B1 => n7495, B2 => n7497, A => n7509, ZN => 
                           IF_RegsxN659);
   U8099 : NAND2_X1 port map( A1 => toRegsPortxDSTxx4x, A2 => n7536, ZN => 
                           n7507);
   U8100 : OR2_X1 port map( A1 => n7540, A2 => n7507, ZN => n7505);
   U8101 : OAI21_X1 port map( B1 => n7495, B2 => n7505, A => n7520, ZN => 
                           IF_RegsxN692);
   U8102 : NOR2_X1 port map( A1 => toRegsPortxDSTxx1x, A2 => n7496, ZN => n7511
                           );
   U8103 : INV_X1 port map( A => n7511, ZN => n7498);
   U8104 : OAI21_X1 port map( B1 => n7498, B2 => n7497, A => n7523, ZN => 
                           IF_RegsxN693);
   U8105 : OAI21_X1 port map( B1 => n7498, B2 => n7505, A => n7520, ZN => 
                           IF_RegsxN694);
   U8106 : NAND4_X1 port map( A1 => toRegsPortxDSTxx1x, A2 => toRegsPort_notify
                           , A3 => toRegsPortxDSTxx3x, A4 => n7537, ZN => n7513
                           );
   U8107 : OAI21_X1 port map( B1 => n7506, B2 => n7513, A => n7509, ZN => 
                           IF_RegsxN695);
   U8108 : OAI21_X1 port map( B1 => n7507, B2 => n7513, A => n7523, ZN => 
                           IF_RegsxN696);
   U8109 : NAND2_X1 port map( A1 => toRegsPort_notify, A2 => toRegsPortxDSTxx0x
                           , ZN => n7503);
   U8110 : OAI21_X1 port map( B1 => n7503, B2 => n7499, A => n7523, ZN => 
                           IF_RegsxN697);
   U8111 : NAND2_X1 port map( A1 => toRegsPortxDSTxx2x, A2 => n7541, ZN => 
                           n7501);
   U8112 : NOR2_X1 port map( A1 => n7534, A2 => n7501, ZN => n7515);
   U8113 : NAND2_X1 port map( A1 => toRegsPort_notify, A2 => n7515, ZN => n7500
                           );
   U8114 : OAI21_X1 port map( B1 => n7506, B2 => n7500, A => n7509, ZN => 
                           IF_RegsxN699);
   U8115 : OAI21_X1 port map( B1 => n7500, B2 => n7507, A => n7509, ZN => 
                           IF_RegsxN700);
   U8116 : NOR2_X1 port map( A1 => toRegsPortxDSTxx1x, A2 => n7501, ZN => n7504
                           );
   U8117 : NAND2_X1 port map( A1 => toRegsPortxDSTxx4x, A2 => n7504, ZN => 
                           n7502);
   U8118 : OAI21_X1 port map( B1 => n7503, B2 => n7502, A => n7509, ZN => 
                           IF_RegsxN701);
   U8119 : INV_X1 port map( A => n7504, ZN => n7519);
   U8120 : OAI21_X1 port map( B1 => n7505, B2 => n7519, A => n7520, ZN => 
                           IF_RegsxN702);
   U8121 : NAND4_X1 port map( A1 => toRegsPortxDSTxx1x, A2 => toRegsPort_notify
                           , A3 => n7541, A4 => n7537, ZN => n7522);
   U8122 : OAI21_X1 port map( B1 => n7506, B2 => n7522, A => n7520, ZN => 
                           IF_RegsxN703);
   U8123 : OAI21_X1 port map( B1 => n7507, B2 => n7522, A => n7509, ZN => 
                           IF_RegsxN704);
   U8124 : NAND4_X1 port map( A1 => toRegsPort_notify, A2 => n7541, A3 => n7534
                           , A4 => n7537, ZN => n7525);
   U8125 : OAI21_X1 port map( B1 => n7506, B2 => n7525, A => n7520, ZN => 
                           IF_RegsxN705);
   U8126 : OAI21_X1 port map( B1 => n7507, B2 => n7525, A => n7523, ZN => 
                           IF_RegsxN706);
   U8127 : NAND3_X1 port map( A1 => toRegsPort_notify, A2 => n7508, A3 => n7539
                           , ZN => n7510);
   U8128 : OAI21_X1 port map( B1 => n7536, B2 => n7510, A => n7509, ZN => 
                           IF_RegsxN707);
   U8129 : OAI21_X1 port map( B1 => toRegsPortxDSTxx0x, B2 => n7510, A => n7520
                           , ZN => IF_RegsxN708);
   U8130 : NAND3_X1 port map( A1 => toRegsPort_notify, A2 => n7511, A3 => n7539
                           , ZN => n7512);
   U8131 : OAI21_X1 port map( B1 => n7536, B2 => n7512, A => n7520, ZN => 
                           IF_RegsxN709);
   U8132 : OAI21_X1 port map( B1 => toRegsPortxDSTxx0x, B2 => n7512, A => n7520
                           , ZN => IF_RegsxN710);
   U8133 : NAND2_X1 port map( A1 => toRegsPortxDSTxx0x, A2 => n7539, ZN => 
                           n7524);
   U8134 : OAI21_X1 port map( B1 => n7513, B2 => n7524, A => n7523, ZN => 
                           IF_RegsxN711);
   U8135 : NAND2_X1 port map( A1 => n7536, A2 => n7539, ZN => n7521);
   U8136 : OAI21_X1 port map( B1 => n7513, B2 => n7521, A => n7520, ZN => 
                           IF_RegsxN712);
   U8137 : OR2_X1 port map( A1 => n7540, A2 => n7524, ZN => n7517);
   U8138 : OAI21_X1 port map( B1 => n7514, B2 => n7517, A => n7520, ZN => 
                           IF_RegsxN713);
   U8139 : OR2_X1 port map( A1 => n7540, A2 => n7521, ZN => n7518);
   U8140 : OAI21_X1 port map( B1 => n7514, B2 => n7518, A => n7520, ZN => 
                           IF_RegsxN714);
   U8141 : INV_X1 port map( A => n7515, ZN => n7516);
   U8142 : OAI21_X1 port map( B1 => n7516, B2 => n7517, A => n7520, ZN => 
                           IF_RegsxN715);
   U8143 : OAI21_X1 port map( B1 => n7516, B2 => n7518, A => n7520, ZN => 
                           IF_RegsxN716);
   U8144 : OAI21_X1 port map( B1 => n7519, B2 => n7517, A => n7520, ZN => 
                           IF_RegsxN717);
   U8145 : OAI21_X1 port map( B1 => n7519, B2 => n7518, A => n7520, ZN => 
                           IF_RegsxN718);
   U8146 : OAI21_X1 port map( B1 => n7522, B2 => n7524, A => n7520, ZN => 
                           IF_RegsxN719);
   U8147 : OAI21_X1 port map( B1 => n7522, B2 => n7521, A => n7520, ZN => 
                           IF_RegsxN720);
   U8148 : OAI21_X1 port map( B1 => n7525, B2 => n7524, A => n7523, ZN => 
                           IF_RegsxN721);
   U8149 : NAND2_X1 port map( A1 => n7527, A2 => n7526, ZN => IF_ISAxN10935);
   U8150 : NAND2_X1 port map( A1 => n7538, A2 => n7535, ZN => n7529);
   U8151 : INV_X1 port map( A => IF_ISAxN10935, ZN => n7528);
   U8152 : OAI211_X1 port map( C1 => IF_ISAxsection_0_port, C2 => n7529, A => 
                           n7528, B => toRegsPort_notify, ZN => n7530);
   U8153 : OAI211_X1 port map( C1 => n7533, C2 => n7532, A => n7531, B => n7530
                           , ZN => n3458);
   clk_gate_IF_ISAxtoMemoryPort_notify_reg : SNPS_CLOCK_GATE_HIGH_CPU_0 port 
                           map( CLK => clk, EN => IF_ISAxN10829, ENCLK => 
                           net325226);
   clk_gate_IF_ISAxtoRegsPort_regxDSTDATAx : SNPS_CLOCK_GATE_HIGH_CPU_36 port 
                           map( CLK => clk, EN => IF_ISAxN10935, ENCLK => 
                           net325231);
   clk_gate_IF_ISAxtoRegsPort_regxDSTx : SNPS_CLOCK_GATE_HIGH_CPU_35 port map( 
                           CLK => clk, EN => IF_ISAxN10969, ENCLK => net325236)
                           ;
   clk_gate_IF_ISAxpcReg_signal_reg : SNPS_CLOCK_GATE_HIGH_CPU_34 port map( CLK
                           => clk, EN => IF_ISAxN10902, ENCLK => net325241);
   clk_gate_IF_ISAxtoMemoryPort_regxREQx : SNPS_CLOCK_GATE_HIGH_CPU_33 port 
                           map( CLK => clk, EN => IF_ISAxN10832, ENCLK => 
                           net325246);
   clk_gate_IF_ISAxtoMemoryPort_regxADDRINx : SNPS_CLOCK_GATE_HIGH_CPU_32 port 
                           map( CLK => clk, EN => IF_ISAxN10869, ENCLK => 
                           net325251);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_31x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_31 port map( CLK => clk, EN
                           => IF_RegsxN659, ENCLK => net325256);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_30x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_30 port map( CLK => clk, EN
                           => IF_RegsxN692, ENCLK => net325261);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_29x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_29 port map( CLK => clk, EN
                           => IF_RegsxN693, ENCLK => net325266);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_28x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_28 port map( CLK => clk, EN
                           => IF_RegsxN694, ENCLK => net325271);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_27x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_27 port map( CLK => clk, EN
                           => IF_RegsxN695, ENCLK => net325276);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_26x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_26 port map( CLK => clk, EN
                           => IF_RegsxN696, ENCLK => net325281);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_25x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_25 port map( CLK => clk, EN
                           => IF_RegsxN697, ENCLK => net325286);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_24x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_24 port map( CLK => clk, EN
                           => IF_RegsxN698, ENCLK => net325291);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_23x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_23 port map( CLK => clk, EN
                           => IF_RegsxN699, ENCLK => net325296);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_22x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_22 port map( CLK => clk, EN
                           => IF_RegsxN700, ENCLK => net325301);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_21x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_21 port map( CLK => clk, EN
                           => IF_RegsxN701, ENCLK => net325306);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_20x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_20 port map( CLK => clk, EN
                           => IF_RegsxN702, ENCLK => net325311);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_19x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_19 port map( CLK => clk, EN
                           => IF_RegsxN703, ENCLK => net325316);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_18x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_18 port map( CLK => clk, EN
                           => IF_RegsxN704, ENCLK => net325321);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_17x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_17 port map( CLK => clk, EN
                           => IF_RegsxN705, ENCLK => net325326);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_16x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_16 port map( CLK => clk, EN
                           => IF_RegsxN706, ENCLK => net325331);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_15x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_15 port map( CLK => clk, EN
                           => IF_RegsxN707, ENCLK => net325336);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_14x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_14 port map( CLK => clk, EN
                           => IF_RegsxN708, ENCLK => net325341);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_13x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_13 port map( CLK => clk, EN
                           => IF_RegsxN709, ENCLK => net325346);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_12x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_12 port map( CLK => clk, EN
                           => IF_RegsxN710, ENCLK => net325351);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_11x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_11 port map( CLK => clk, EN
                           => IF_RegsxN711, ENCLK => net325356);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_10x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_10 port map( CLK => clk, EN
                           => IF_RegsxN712, ENCLK => net325361);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_09x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_9 port map( CLK => clk, EN 
                           => IF_RegsxN713, ENCLK => net325366);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_08x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_8 port map( CLK => clk, EN 
                           => IF_RegsxN714, ENCLK => net325371);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_07x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_7 port map( CLK => clk, EN 
                           => IF_RegsxN715, ENCLK => net325376);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_06x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_6 port map( CLK => clk, EN 
                           => IF_RegsxN716, ENCLK => net325381);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_05x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_5 port map( CLK => clk, EN 
                           => IF_RegsxN717, ENCLK => net325386);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_04x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_4 port map( CLK => clk, EN 
                           => IF_RegsxN718, ENCLK => net325391);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_03x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_3 port map( CLK => clk, EN 
                           => IF_RegsxN719, ENCLK => net325396);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_02x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_2 port map( CLK => clk, EN 
                           => IF_RegsxN720, ENCLK => net325401);
   clk_gate_IF_RegsxRegsToCtl_port_regxREG_FILE_01x : 
                           SNPS_CLOCK_GATE_HIGH_CPU_1 port map( CLK => clk, EN 
                           => IF_RegsxN721, ENCLK => net325406);
   U3773 : INV_X1 port map( A => n7628, ZN => toMemoryPortxREQxx1x(0));
   n7628 <= '1';

end SYN_CPU_arch;
