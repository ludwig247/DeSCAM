package testbasic15_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic15_SECTIONS;

endpackage
