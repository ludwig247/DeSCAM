package testmasterslave1_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave1_SECTIONS;

endpackage
