library ieee;
use IEEE.numeric_std.all;

package TestFunction0_types is
type TestFunction0_SECTIONS is (run);
end package TestFunction0_types;
