package testbasic13_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic13_SECTIONS;

endpackage
