library ieee;
use IEEE.numeric_std.all;
use work.SCAM_Model_types.all;

package TestBasic13_types is
type Sections is (SECTION_A, SECTION_B);
end package TestBasic13_types;