package testbasic6_types;

endpackage