package testmasterslave9_types;

	typedef enum logic {
		section_a,
		section_b
	} TestMasterSlave9_SECTIONS;

endpackage
