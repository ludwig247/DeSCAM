library ieee;
use IEEE.numeric_std.all;

package TestBasic23_types is
type TestBasic23_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic23_types;
