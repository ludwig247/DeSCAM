package testbasic11_types;

	typedef enum logic {
		section_a,
		section_b
	} TestBasic11_SECTIONS;

endpackage
