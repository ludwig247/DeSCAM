package SCAM_Model_types is
subtype bool is Boolean;
subtype int is Integer;
type Mip_SECTIONS is (run);
end package SCAM_Model_types;
