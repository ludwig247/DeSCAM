package testbasic3_types;

	import scam_model_types::*;
endpackage