package testbasic5_types;

endpackage