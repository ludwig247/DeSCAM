package testfunction1_types;

	typedef enum logic {
		run
	} TestFunction1_SECTIONS;

endpackage
