library ieee;
use IEEE.numeric_std.all;

package TestMasterSlave7_types is
type TestMasterSlave7_SECTIONS is (SECTION_A, SECTION_B);
end package TestMasterSlave7_types;

