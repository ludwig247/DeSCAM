library ieee;
use IEEE.numeric_std.all;

package TestBasic15_types is
type TestBasic15_SECTIONS is (SECTION_A, SECTION_B);
end package TestBasic15_types;
