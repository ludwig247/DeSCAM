library ieee;
use IEEE.numeric_std.all;
use work.top_level_types.all;

package TestMasterSlave00_types is
type Phases is (SECTION_A, SECTION_B);
end package TestMasterSlave00_types;