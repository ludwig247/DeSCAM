library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.SCAM_Model_types.all;

entity Regs is
port(	
	RFtoISA_port_sig: out RegfileType;
	ISAtoRF_port_sig: in RegfileWriteType;
	ISAtoRF_port_sync: in boolean;
	clk: in std_logic;
	rst: in std_logic
);
end Regs;

architecture Regs_arch of Regs is
	-- Define internal data types
	type Regs_assign_t is (assign_0, assign_1, assign_2, assign_3, assign_4, assign_5, assign_6, assign_7, assign_8, assign_9, assign_10, assign_11, assign_12, assign_13, assign_14, assign_15, assign_16, assign_17, assign_18, assign_19, assign_20, assign_21, assign_22, assign_23, assign_24);
	type Regs_state_t is (st_run_0);

	-- Declare signals
	signal active_state: Regs_state_t;
	signal active_assignment: Regs_assign_t;
	--signal --reg_file_01: unsigned(31 downto 0);
	--signal --reg_file_02: unsigned(31 downto 0);
	--signal --reg_file_06: unsigned(31 downto 0);
	--signal --reg_file_07: unsigned(31 downto 0);
	--signal --reg_file_08: unsigned(31 downto 0);
	--signal --reg_file_09: unsigned(31 downto 0);
	--signal --reg_file_10: unsigned(31 downto 0);
	--signal --reg_file_11: unsigned(31 downto 0);
	--signal --reg_file_12: unsigned(31 downto 0);
	--signal --reg_file_13: unsigned(31 downto 0);
	--signal --reg_file_14: unsigned(31 downto 0);
	--signal --reg_file_15: unsigned(31 downto 0);
	--signal --reg_file_16: unsigned(31 downto 0);
	--signal --reg_file_17: unsigned(31 downto 0);
	--signal --reg_file_18: unsigned(31 downto 0);
	--signal --reg_file_19: unsigned(31 downto 0);
	--signal --reg_file_20: unsigned(31 downto 0);
	--signal --reg_file_21: unsigned(31 downto 0);
	--signal --reg_file_22: unsigned(31 downto 0);
	--signal --reg_file_23: unsigned(31 downto 0);
	--signal --reg_file_24: unsigned(31 downto 0);
	--signal --reg_file_25: unsigned(31 downto 0);
	--signal --reg_file_26: unsigned(31 downto 0);
	--signal --reg_file_27: unsigned(31 downto 0);

	-- Declare state signals that are used by ITL properties for OneSpin
	signal run_0: boolean;


begin
	-- Combinational logic that selects current operation
	process (active_state, ISAtoRF_port_sync, ISAtoRF_port_sig.dst)
	begin
		case active_state is
		when st_run_0 =>
			if (not(ISAtoRF_port_sync)) then 
				-- Operation: op_run_0_write_0;
				active_assignment <= assign_0;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000000") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_1;
				active_assignment <= assign_0;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000001") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_2;
				active_assignment <= assign_1;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000002") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_3;
				active_assignment <= assign_2;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000006") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_4;
				active_assignment <= assign_3;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000007") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_5;
				active_assignment <= assign_4;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000008") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_6;
				active_assignment <= assign_5;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000009") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_7;
				active_assignment <= assign_6;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000000a") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_8;
				active_assignment <= assign_7;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000000b") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_9;
				active_assignment <= assign_8;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000000c") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_10;
				active_assignment <= assign_9;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000000d") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_11;
				active_assignment <= assign_10;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000000e") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_12;
				active_assignment <= assign_11;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000000f") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_13;
				active_assignment <= assign_12;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000010") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_14;
				active_assignment <= assign_13;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000011") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_15;
				active_assignment <= assign_14;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000012") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_16;
				active_assignment <= assign_15;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000013") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_17;
				active_assignment <= assign_16;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000014") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_18;
				active_assignment <= assign_17;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000015") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_19;
				active_assignment <= assign_18;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000016") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_20;
				active_assignment <= assign_19;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000017") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_21;
				active_assignment <= assign_20;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000018") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_22;
				active_assignment <= assign_21;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"00000019") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_23;
				active_assignment <= assign_22;
			elsif (ISAtoRF_port_sync and (ISAtoRF_port_sig.dst = x"0000001a") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_24;
				active_assignment <= assign_23;
			else--if(ISAtoRF_port_sync and not(ISAtoRF_port_sig.dst = x"00000000") and not(ISAtoRF_port_sig.dst = x"00000001") and not(ISAtoRF_port_sig.dst = x"00000002") and not(ISAtoRF_port_sig.dst = x"00000006") and not(ISAtoRF_port_sig.dst = x"00000007") and not(ISAtoRF_port_sig.dst = x"00000008") and not(ISAtoRF_port_sig.dst = x"00000009") and not(ISAtoRF_port_sig.dst = x"0000000a") and not(ISAtoRF_port_sig.dst = x"0000000b") and not(ISAtoRF_port_sig.dst = x"0000000c") and not(ISAtoRF_port_sig.dst = x"0000000d") and not(ISAtoRF_port_sig.dst = x"0000000e") and not(ISAtoRF_port_sig.dst = x"0000000f") and not(ISAtoRF_port_sig.dst = x"00000010") and not(ISAtoRF_port_sig.dst = x"00000011") and not(ISAtoRF_port_sig.dst = x"00000012") and not(ISAtoRF_port_sig.dst = x"00000013") and not(ISAtoRF_port_sig.dst = x"00000014") and not(ISAtoRF_port_sig.dst = x"00000015") and not(ISAtoRF_port_sig.dst = x"00000016") and not(ISAtoRF_port_sig.dst = x"00000017") and not(ISAtoRF_port_sig.dst = x"00000018") and not(ISAtoRF_port_sig.dst = x"00000019") and not(ISAtoRF_port_sig.dst = x"0000001a") and ISAtoRF_port_sync) then 
				-- Operation: op_run_0_write_25;
				active_assignment <= assign_24;
			end if;
		end case;
	end process;

	-- Main process
	process (clk, rst)
	begin
		if (rst = '1') then
			RFtoISA_port_sig.reg_file_25 <= x"00000000";
			RFtoISA_port_sig.reg_file_18 <= x"00000000";
			RFtoISA_port_sig.reg_file_17 <= x"00000000";
			RFtoISA_port_sig.reg_file_02 <= x"00000000";
			RFtoISA_port_sig.reg_file_13 <= x"00000000";
			--reg_file_15 <= x"00000000";
			--reg_file_02 <= x"00000000";
			RFtoISA_port_sig.reg_file_19 <= x"00000000";
			--reg_file_27 <= x"00000000";
			--reg_file_23 <= x"00000000";
			RFtoISA_port_sig.reg_file_20 <= x"00000000";
			RFtoISA_port_sig.reg_file_08 <= x"00000000";
			RFtoISA_port_sig.reg_file_27 <= x"00000000";
			RFtoISA_port_sig.reg_file_21 <= x"00000000";
			RFtoISA_port_sig.reg_file_22 <= x"00000000";
			RFtoISA_port_sig.reg_file_15 <= x"00000000";
			RFtoISA_port_sig.reg_file_23 <= x"00000000";
			RFtoISA_port_sig.reg_file_14 <= x"00000000";
			--reg_file_08 <= x"00000000";
			--reg_file_13 <= x"00000000";
			RFtoISA_port_sig.reg_file_11 <= x"00000000";
			--reg_file_01 <= x"00000000";
			--reg_file_25 <= x"00000000";
			RFtoISA_port_sig.reg_file_26 <= x"00000000";
			--reg_file_21 <= x"00000000";
			active_state <= st_run_0;
			RFtoISA_port_sig.reg_file_12 <= x"00000000";
			--reg_file_22 <= x"00000000";
			RFtoISA_port_sig.reg_file_16 <= x"00000000";
			RFtoISA_port_sig.reg_file_01 <= x"00000000";
			--reg_file_12 <= x"00000000";
			--reg_file_10 <= x"00000000";
			--reg_file_18 <= x"00000000";
			--reg_file_16 <= x"00000000";
			--reg_file_26 <= x"00000000";
			--reg_file_20 <= x"00000000";
			--reg_file_07 <= x"00000000";
			--reg_file_11 <= x"00000000";
			--reg_file_14 <= x"00000000";
			--reg_file_09 <= x"00000000";
			RFtoISA_port_sig.reg_file_07 <= x"00000000";
			--reg_file_06 <= x"00000000";
			RFtoISA_port_sig.reg_file_09 <= x"00000000";
			RFtoISA_port_sig.reg_file_06 <= x"00000000";
			--reg_file_17 <= x"00000000";
			RFtoISA_port_sig.reg_file_24 <= x"00000000";
			--reg_file_24 <= x"00000000";
			RFtoISA_port_sig.reg_file_10 <= x"00000000";
			--reg_file_19 <= x"00000000";
		elsif (clk = '1' and clk'event) then
			case active_assignment is
			when assign_0 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_1 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				RFtoISA_port_sig.reg_file_01 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--reg_file_01 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_2 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				RFtoISA_port_sig.reg_file_02 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--reg_file_02 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_3 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--reg_file_06 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				RFtoISA_port_sig.reg_file_06 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_4 =>
				RFtoISA_port_sig.reg_file_07 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--reg_file_07 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_5 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--reg_file_08 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				RFtoISA_port_sig.reg_file_08 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_6 =>
				RFtoISA_port_sig.reg_file_09 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--reg_file_09 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
			when assign_7 =>
				--reg_file_10 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				RFtoISA_port_sig.reg_file_10 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_8 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				RFtoISA_port_sig.reg_file_11 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--reg_file_11 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_9 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--reg_file_12 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
				RFtoISA_port_sig.reg_file_12 <= ISAtoRF_port_sig.dstData;
			when assign_10 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				RFtoISA_port_sig.reg_file_13 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--reg_file_13 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_11 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--reg_file_14 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				RFtoISA_port_sig.reg_file_14 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_12 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--reg_file_15 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				RFtoISA_port_sig.reg_file_15 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_13 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				RFtoISA_port_sig.reg_file_16 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--reg_file_16 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_14 =>
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				RFtoISA_port_sig.reg_file_17 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--reg_file_17 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_15 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--reg_file_18 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				RFtoISA_port_sig.reg_file_18 <= ISAtoRF_port_sig.dstData;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_16 =>
				RFtoISA_port_sig.reg_file_19 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--reg_file_19 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_17 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--reg_file_20 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				RFtoISA_port_sig.reg_file_20 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_18 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				RFtoISA_port_sig.reg_file_21 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--reg_file_21 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_19 =>
				--reg_file_22 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				RFtoISA_port_sig.reg_file_22 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_20 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				RFtoISA_port_sig.reg_file_23 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--reg_file_23 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_21 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--reg_file_24 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				RFtoISA_port_sig.reg_file_24 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_22 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				RFtoISA_port_sig.reg_file_25 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--reg_file_25 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_23 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_27 <= --reg_file_27;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--reg_file_26 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				RFtoISA_port_sig.reg_file_26 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			when assign_24 =>
				--RFtoISA_port_sig.reg_file_17 <= --reg_file_17;
				--RFtoISA_port_sig.reg_file_13 <= --reg_file_13;
				--RFtoISA_port_sig.reg_file_16 <= --reg_file_16;
				--RFtoISA_port_sig.reg_file_06 <= --reg_file_06;
				--RFtoISA_port_sig.reg_file_07 <= --reg_file_07;
				--RFtoISA_port_sig.reg_file_08 <= --reg_file_08;
				--RFtoISA_port_sig.reg_file_11 <= --reg_file_11;
				RFtoISA_port_sig.reg_file_27 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_25 <= --reg_file_25;
				--RFtoISA_port_sig.reg_file_14 <= --reg_file_14;
				--RFtoISA_port_sig.reg_file_18 <= --reg_file_18;
				--RFtoISA_port_sig.reg_file_21 <= --reg_file_21;
				--RFtoISA_port_sig.reg_file_20 <= --reg_file_20;
				active_state <= st_run_0;
				--RFtoISA_port_sig.reg_file_15 <= --reg_file_15;
				--RFtoISA_port_sig.reg_file_26 <= --reg_file_26;
				--RFtoISA_port_sig.reg_file_23 <= --reg_file_23;
				--reg_file_27 <= ISAtoRF_port_sig.dstData;
				--RFtoISA_port_sig.reg_file_10 <= --reg_file_10;
				--RFtoISA_port_sig.reg_file_01 <= --reg_file_01;
				--RFtoISA_port_sig.reg_file_02 <= --reg_file_02;
				--RFtoISA_port_sig.reg_file_12 <= --reg_file_12;
				--RFtoISA_port_sig.reg_file_22 <= --reg_file_22;
				--RFtoISA_port_sig.reg_file_24 <= --reg_file_24;
				--RFtoISA_port_sig.reg_file_19 <= --reg_file_19;
				--RFtoISA_port_sig.reg_file_09 <= --reg_file_09;
			end case;
		end if;
	end process;

	-- Assigning state signals that are used by ITL properties for OneSpin
	run_0 <= active_state = st_run_0;

end Regs_arch;

